module osc_core (
    input glob_en,
    input [3:0] delay_con_lsb,
    input [6:0] delay_con_msb,
    input [3:0] con_perb,

    output osc_000,
    output osc_036,
    output osc_072,
    output osc_144,
    output osc_180

// 
// waiting to integrate the ref_injector
//  

// 
// buffered output phase, goes to phase blender
// 

)



