###########################
# Greatest Common Divisor #
###########################
