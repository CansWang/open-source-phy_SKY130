magic
tech sky130A
<<<<<<< HEAD
timestamp 1619949044
<< dnwell >>
rect 759 5481 877 5599
rect 534 4966 652 5084
rect 776 5003 894 5121
rect 1012 4985 1130 5103
rect 1255 4965 1373 5083
rect 1441 4969 1559 5087
rect 1631 4976 1749 5094
<< metal3 >>
rect 2939 -652 4545 66
<< via4 >>
rect 88 5407 206 5525
rect 526 5420 644 5538
rect 759 5481 877 5599
rect 534 4966 652 5084
rect 776 5003 894 5121
rect 1012 4985 1130 5103
rect 1255 4965 1373 5083
rect 1441 4969 1559 5087
rect 1631 4976 1749 5094
<< metal5 >>
rect 2908 19715 4514 20433
rect -1030 19099 -467 19126
rect -1030 17920 1759 19099
rect -1030 6258 -467 17920
rect 2882 15120 4488 15838
rect 7922 7728 8606 7782
rect 6951 7213 8606 7728
rect 0 6744 427 7130
rect -1408 5525 468 6258
rect -1408 5407 88 5525
rect 206 5407 468 5525
rect -1408 3981 468 5407
rect -1408 3890 541 3981
rect -1408 2597 468 3890
rect 7922 2383 8606 7213
rect 385 319 1347 2349
rect 7206 2042 8606 2383
rect 7206 2035 8539 2042
use test  test_0
timestamp 1619945680
transform 1 0 0 0 1 0
box 0 0 7500 20000
<< labels >>
flabel metal5 385 319 1347 2349 1 FreeSans 3200 0 0 0 VDD
port 3 n
flabel metal3 2939 -652 4545 66 1 FreeSans 3200 0 0 0 in
port 1 n
flabel metal5 2882 15120 4488 15838 1 FreeSans 3200 0 0 0 out
port 2 n
flabel metal5 2908 19715 4514 20433 1 FreeSans 3200 0 0 0 GND
port 4 n
=======
magscale 1 2
timestamp 1619375533
<< error_p >>
rect 16381 38796 16826 39032
rect 16590 37120 16826 38796
rect 16490 37090 16826 37120
rect 16562 37062 16628 37090
<< error_s >>
rect 3868 39959 9658 40320
rect 3832 39796 9658 39959
rect 9713 39796 9742 39959
rect 14603 38987 16381 39032
rect 235 38804 471 38987
rect 562 38804 798 38987
rect 889 38804 1125 38987
rect 1216 38804 1452 38987
rect 1543 38804 1779 38987
rect 1870 38804 2106 38987
rect 2197 38804 2433 38987
rect 2524 38804 2760 38987
rect 2851 38804 3087 38987
rect 3178 38804 3414 38987
rect 3505 38804 3741 38987
rect 3832 38804 4068 38987
rect 4159 38804 4395 38987
rect 4486 38804 4722 38987
rect 4813 38804 5049 38987
rect 5140 38804 5376 38987
rect 5467 38804 5703 38987
rect 5794 38804 6030 38987
rect 6121 38804 6357 38987
rect 6448 38804 6684 38987
rect 6775 38804 7011 38987
rect 7102 38804 7338 38987
rect 7429 38804 7665 38987
rect 7756 38804 7992 38987
rect 8083 38804 8319 38987
rect 8409 38804 8645 38987
rect 8735 38804 8971 38987
rect 9061 38804 9297 38987
rect 9387 38804 9623 38987
rect 9713 38804 9949 38987
rect 10039 38804 10275 38987
rect 10365 38804 10601 38987
rect 10691 38804 10927 38987
rect 11017 38804 11253 38987
rect 11343 38804 11579 38987
rect 11669 38804 11905 38987
rect 11995 38804 12231 38987
rect 12321 38804 12557 38987
rect 12647 38804 12883 38987
rect 12973 38804 13209 38987
rect 13299 38804 13535 38987
rect 13625 38804 13861 38987
rect 13951 38804 14187 38987
rect 14277 38804 14513 38987
rect 14588 38804 16381 38987
rect -174 38796 16381 38804
rect -174 38784 14839 38796
rect 0 38751 14839 38784
rect 0 38663 14824 38751
rect 0 38427 14839 38663
rect 14890 38427 14923 38608
rect 0 38339 14824 38427
rect 14890 38423 14908 38427
rect 0 38103 14839 38339
rect 14890 38103 14923 38423
rect 0 38015 14824 38103
rect 14890 38099 14908 38103
rect 0 37779 14839 38015
rect 14890 37779 14923 38099
rect 0 37691 14824 37779
rect 14890 37775 14908 37779
rect 0 37455 14839 37691
rect 14890 37455 14923 37775
rect 0 37367 14824 37455
rect 14890 37451 14908 37455
rect 0 37131 14839 37367
rect 14890 37238 14923 37451
rect 0 37110 14824 37131
rect -174 37086 14824 37110
rect 53 18966 118 19030
rect 14812 18966 15258 19030
rect 137 18730 202 18966
rect 14599 18730 15258 18966
rect 53 18630 118 18714
rect 14812 18630 15258 18730
rect 137 18394 202 18630
rect 14599 18394 15258 18630
rect 53 18294 118 18378
rect 14812 18294 15258 18394
rect 137 18058 202 18294
rect 14599 18058 15258 18294
rect 53 17958 118 18042
rect 14812 17958 15258 18058
rect 137 17722 202 17958
rect 14599 17722 15258 17958
rect 53 17622 118 17706
rect 14812 17622 15258 17722
rect 137 17386 202 17622
rect 14599 17386 15258 17622
rect 53 17286 118 17370
rect 14812 17286 15258 17386
rect 137 17050 202 17286
rect 14599 17050 15258 17286
rect 53 16950 118 17034
rect 14812 16950 15258 17050
rect 137 16714 202 16950
rect 14599 16714 15258 16950
rect 53 16614 118 16698
rect 14812 16614 15258 16714
rect 137 16378 202 16614
rect 14599 16378 15258 16614
rect 53 16278 118 16362
rect 14812 16278 15258 16378
rect 137 16042 202 16278
rect 14599 16042 15258 16278
rect 53 15942 118 16026
rect 14812 15942 15258 16042
rect 137 15706 202 15942
rect 14599 15706 15258 15942
rect 53 15606 118 15690
rect 14812 15606 15258 15706
rect 137 15370 202 15606
rect 14599 15370 15258 15606
rect 53 15270 118 15354
rect 14812 15270 15258 15370
rect 137 15034 202 15270
rect 14599 15034 15258 15270
rect 53 14934 118 15018
rect 14812 14934 15258 15034
rect 137 14698 202 14934
rect 14599 14698 15258 14934
rect 53 14598 118 14682
rect 14812 14598 15258 14698
rect 137 14362 202 14598
rect 14599 14362 15258 14598
rect 53 14262 118 14346
rect 14812 14262 15258 14362
rect 137 14026 202 14262
rect 14599 14026 15258 14262
rect 53 13657 118 13741
rect 14812 13657 15258 14026
rect 137 13421 202 13657
rect 14597 13421 15258 13657
rect 53 13091 118 13175
rect 14812 13091 15258 13421
rect 137 12918 202 13091
rect -358 12855 459 12890
rect 14597 12855 15258 13091
rect -358 12831 568 12855
rect 14812 12832 15258 12855
rect 14420 12831 15282 12832
rect -358 12828 254 12831
rect 14812 12830 15282 12831
rect 15258 12806 15282 12830
rect -568 12533 248 12570
rect -569 12532 248 12533
rect -568 12511 248 12532
rect 14740 12511 14812 12512
rect -568 12508 574 12511
rect 15258 12510 15554 12512
rect -568 5202 -544 12508
rect 0 12487 176 12508
rect 0 12251 373 12487
rect 14740 12290 14746 12296
rect 14833 12290 14976 12487
rect 15554 12296 15580 12314
rect 15550 12291 15580 12296
rect 14994 12290 15580 12291
rect 14597 12251 15580 12290
rect 0 11921 176 12251
rect 14740 11921 15580 12251
rect 0 11685 373 11921
rect 14597 11685 15580 11921
rect 0 11641 176 11685
rect 0 11341 177 11641
rect 0 11275 176 11341
rect 0 11215 177 11275
rect 0 10619 176 11215
rect 0 10559 177 10619
rect 14740 10559 15580 11685
rect 0 10323 278 10559
rect 14705 10323 15580 10559
rect 0 10263 177 10323
rect 0 9667 176 10263
rect 0 9607 177 9667
rect 0 9541 176 9607
rect 0 9241 177 9541
rect 0 9197 176 9241
rect 14740 9197 15580 10323
rect 0 8961 373 9197
rect 14599 8961 15580 9197
rect 0 8591 176 8961
rect 14740 8591 15580 8961
rect 0 8355 373 8591
rect 14599 8355 15580 8591
rect 0 8311 176 8355
rect 0 8031 177 8311
rect 0 7987 176 8031
rect 14740 7987 15580 8355
rect 0 7751 373 7987
rect 14599 7751 15580 7987
rect 0 7621 176 7751
rect 14740 7621 15580 7751
rect 0 7385 373 7621
rect 14599 7385 15580 7621
rect 0 7341 176 7385
rect 0 7061 177 7341
rect 0 7017 176 7061
rect 14740 7017 15580 7385
rect 0 6781 373 7017
rect 14599 6781 15580 7017
rect 0 6651 176 6781
rect 14740 6651 15580 6781
rect 0 6415 373 6651
rect 14599 6415 15580 6651
rect 0 6371 176 6415
rect 0 6091 177 6371
rect 0 6047 176 6091
rect 14740 6047 15580 6415
rect 0 5811 373 6047
rect 14599 5811 15580 6047
rect 0 5441 176 5811
rect 14740 5441 15580 5811
rect 0 5205 373 5441
rect 14599 5240 15580 5441
rect 14514 5205 15580 5240
rect 0 5202 176 5205
rect -568 5181 568 5202
rect 14386 5181 15580 5205
rect -568 5166 248 5181
rect -574 5160 248 5166
rect -568 5154 -562 5160
rect 170 5159 177 5160
rect 170 5154 176 5159
rect 14740 5148 15580 5181
rect 14734 5142 15580 5148
rect 14740 5136 14746 5142
rect 15550 5136 15580 5142
rect 15556 5118 15580 5136
rect 14706 4900 14740 4920
rect 176 4861 248 4882
rect 14706 4861 15484 4900
rect 176 4840 568 4861
rect 14732 4837 15484 4861
rect 0 4601 373 4837
rect 14599 4601 15484 4837
rect 0 4231 222 4601
rect 14732 4231 15484 4601
rect 0 3995 373 4231
rect 14599 3995 15484 4231
rect 0 3627 222 3995
rect 14732 3627 15484 3995
rect 0 3391 373 3627
rect 14599 3391 15484 3627
rect 0 3261 222 3391
rect 14732 3261 15484 3391
rect 0 3025 373 3261
rect 14599 3025 15484 3261
rect 0 2657 222 3025
rect 14732 2657 15484 3025
rect 0 2421 373 2657
rect 14599 2421 15484 2657
rect 0 2051 222 2421
rect 14732 2051 15484 2421
rect 0 1815 373 2051
rect 14599 1815 15484 2051
rect 0 1446 222 1815
rect 14732 1446 15484 1815
rect 0 1210 373 1446
rect 14599 1210 15484 1446
rect 0 1064 222 1210
rect 14732 1186 15484 1210
rect 14732 1181 15490 1186
rect 14732 1180 15491 1181
rect 14732 1064 15514 1180
rect 0 828 373 1064
rect 14599 828 15514 1064
rect 0 682 222 828
rect 14732 682 15514 828
rect 0 446 373 682
rect 14599 462 15514 682
rect 14599 446 15491 462
rect 0 310 222 446
rect 14732 386 15491 446
rect 14738 0 15491 386
rect 14738 -868 14739 0
rect 15489 -520 15491 0
rect 15466 -542 15491 -520
rect 15182 -544 15828 -542
rect 15182 -838 15514 -544
rect 15182 -862 15532 -838
rect 14732 -873 14739 -868
rect 15442 -873 15566 -862
rect 14732 -874 15566 -873
rect 14738 -880 14744 -874
rect 15484 -875 15491 -874
rect 15484 -880 15490 -875
rect 15502 -880 15532 -874
rect 15508 -898 15532 -880
<< psubdiff >>
rect 3382 39796 3868 40496
rect 9658 39796 10356 40496
rect 3382 39522 10356 39796
<< psubdiffcont >>
rect 3868 39796 9658 40496
<< locali >>
rect 3382 40496 10356 40856
rect 3382 39796 3868 40496
rect 9658 39796 10356 40496
rect 3382 39522 10356 39796
<< viali >>
rect 3868 39796 9658 40496
<< metal1 >>
rect 3382 40496 10356 40856
rect 3382 39796 3868 40496
rect 9658 39796 10356 40496
rect 3382 39522 10356 39796
<< via1 >>
rect 3868 39796 9658 40496
<< metal2 >>
rect 3382 40496 10356 40856
rect 3382 39796 3868 40496
rect 9658 39796 10356 40496
rect 3382 39522 10356 39796
<< via2 >>
rect 3868 39796 9658 40496
<< metal3 >>
rect 3382 40496 10356 40856
rect 3382 39796 3868 40496
rect 9658 39796 10356 40496
rect 3382 39522 10356 39796
rect -3174 38808 -162 38818
rect -3174 38608 18208 38808
rect -3174 38590 14890 38608
rect -3174 37214 -1478 38590
rect -108 37238 14890 38590
rect 16440 37238 18208 38608
rect -108 37214 18208 37238
rect -3174 37090 18208 37214
rect -3174 15370 -1632 37090
rect -3174 13964 -1628 15370
rect -400 13964 118 15370
rect -3174 12532 -1632 13964
rect -3174 11002 -568 12532
rect -570 10578 -568 11002
rect 17060 11450 18208 37090
rect 15556 11446 18486 11450
rect 15556 9990 18488 11446
rect 15556 9940 16936 9990
rect 4144 -424 10462 192
rect 5606 -986 8772 -424
<< via3 >>
rect 3868 39796 9658 40496
rect -1478 37214 -108 38590
rect 14890 37238 16440 38608
rect -568 5160 176 12532
rect 14740 5142 15556 12290
rect 14738 -874 15490 1180
rect 15502 -874 15508 -862
<< mimcap >>
rect 14744 38796 16594 38798
rect 16590 37120 16594 38796
rect 16590 37090 16600 37120
<< metal4 >>
rect 3382 40496 10356 40856
rect 3382 39796 3868 40496
rect 9658 39796 10356 40496
rect 3382 39522 10356 39796
rect -1626 38804 258 38812
rect 14714 38804 16598 38808
rect -1626 38590 -174 38804
rect 14824 38798 16598 38804
rect 14824 38608 16590 38796
rect -1626 37214 -1478 38590
rect 14824 37238 14890 38608
rect 16440 37238 16590 38608
rect -1626 37086 -174 37214
rect 14824 37090 16590 37238
rect 16594 37120 16598 38798
rect 14824 37086 16598 37090
rect 14714 37082 16598 37086
rect 4354 29812 10364 30094
rect 4354 27544 5108 29812
rect 9590 27544 10364 29812
rect 4354 27012 10364 27544
rect 222 2940 2300 3716
rect 12772 2944 14732 3720
<< via4 >>
rect 3868 39796 9658 40496
rect -174 38798 14824 38804
rect -174 38796 16594 38798
rect -174 38590 14824 38796
rect -1478 37214 -108 38590
rect -108 37214 14824 38590
rect 14890 37238 16440 38608
rect -174 37086 14824 37214
rect 16590 37120 16594 38796
rect 16590 37090 16600 37120
rect 5108 27544 9590 29812
rect -226 12918 118 19030
rect 14812 12830 15258 19030
rect -568 5160 176 12532
rect 14740 5142 15556 12290
rect -490 310 222 4818
rect 14732 1180 15484 4900
rect 14732 386 14738 1180
rect 14738 -874 15490 1180
rect 15502 -874 15508 -862
<< metal5 >>
rect 3382 40496 10356 40856
rect 3382 39796 3868 40496
rect 9658 39796 10356 40496
rect 3382 39522 10356 39796
rect -1634 38804 208 38808
rect 3856 38804 8982 39522
rect -1634 38590 -174 38804
rect 14824 38798 16596 38802
rect 14824 38608 16590 38796
rect -1634 37214 -1478 38590
rect 14824 37238 14890 38608
rect 16440 37238 16590 38608
rect -1634 37086 -174 37214
rect 14824 37090 16590 37238
rect 16594 37120 16596 38798
rect 4354 29812 10364 30094
rect -1008 28520 -180 29640
rect -1008 24690 1558 28520
rect 4354 27544 5108 29812
rect 9590 27544 10364 29812
rect 4354 27012 10364 27544
rect -1008 23980 -180 24690
rect -358 19030 254 19096
rect -358 18770 -226 19030
rect -1554 16280 -226 18770
rect -1628 15858 -226 16280
rect -2480 13774 -226 15858
rect -2480 12430 -1216 13774
rect -358 12918 -226 13774
rect 118 12918 254 19030
rect -358 12828 254 12918
rect 14740 19030 15352 19092
rect 14740 12832 14812 19030
rect 15258 16030 15352 19030
rect 16420 16030 17094 16174
rect 15258 14882 17094 16030
rect 15258 12832 15352 14882
rect -568 12532 248 12570
rect -2480 1968 -1230 12430
rect 176 5160 248 12532
rect 14740 12290 15554 12512
rect 14706 4900 15492 4920
rect -538 4818 248 4882
rect -538 1968 -490 4818
rect -2480 432 -490 1968
rect -538 310 -490 432
rect 222 310 248 4818
rect -538 -1560 248 310
rect 14706 386 14732 4900
rect 15484 1212 15492 4900
rect 15484 1180 15490 1212
rect 16420 462 17094 14882
rect 14706 -874 14738 386
rect 15490 -544 17754 462
rect 14706 -1560 15492 -874
rect -538 -5424 15512 -1560
rect -538 -5490 248 -5424
rect 14706 -5452 15492 -5424
use test  test_0
timestamp 1619375533
transform 1 0 -6 0 1 -6
box 0 0 15000 40000
<< labels >>
flabel metal5 3382 40496 10356 40856 1 FreeSans 6400 0 0 0 GND
port 4 n
flabel metal5 -1008 23980 -180 29640 1 FreeSans 6400 0 0 0 out
port 2 n
flabel metal5 -538 -5424 15512 -1560 1 FreeSans 6400 0 0 0 VDD
port 3 n
flabel metal3 5606 -986 8772 -380 1 FreeSans 6400 0 0 0 in
port 1 n
>>>>>>> 4fc8ec152ed10a0bfcaa5005507078aaca6a9b6b
<< end >>
