magic
tech sky130A
magscale 1 2
timestamp 1619862920
<< checkpaint >>
rect -1267 -1488 2778 3936
<< nwell >>
rect 0 2537 670 2676
rect -5 1465 670 2537
rect -7 -52 643 1189
<< pwell >>
rect 800 1556 1436 2208
rect 835 1142 1249 1149
rect 835 97 1365 1142
rect 1279 93 1365 97
<< nmos >>
rect 879 1582 929 2182
rect 985 1582 1035 2182
rect 1201 1582 1251 2182
rect 1307 1582 1357 2182
<< mvnmos >>
rect 914 123 1014 1123
rect 1070 123 1170 1123
<< mvpmos >>
rect 112 123 212 1123
rect 268 123 368 1123
rect 424 123 524 1123
<< pmoshvt >>
rect 84 1501 134 2501
rect 190 1501 240 2501
rect 407 1501 457 2501
rect 513 1501 563 2501
<< ndiff >>
rect 826 2170 879 2182
rect 826 2136 834 2170
rect 868 2136 879 2170
rect 826 2102 879 2136
rect 826 2068 834 2102
rect 868 2068 879 2102
rect 826 2034 879 2068
rect 826 2000 834 2034
rect 868 2000 879 2034
rect 826 1966 879 2000
rect 826 1932 834 1966
rect 868 1932 879 1966
rect 826 1898 879 1932
rect 826 1864 834 1898
rect 868 1864 879 1898
rect 826 1830 879 1864
rect 826 1796 834 1830
rect 868 1796 879 1830
rect 826 1762 879 1796
rect 826 1728 834 1762
rect 868 1728 879 1762
rect 826 1694 879 1728
rect 826 1660 834 1694
rect 868 1660 879 1694
rect 826 1582 879 1660
rect 929 2170 985 2182
rect 929 2136 940 2170
rect 974 2136 985 2170
rect 929 2102 985 2136
rect 929 2068 940 2102
rect 974 2068 985 2102
rect 929 2034 985 2068
rect 929 2000 940 2034
rect 974 2000 985 2034
rect 929 1966 985 2000
rect 929 1932 940 1966
rect 974 1932 985 1966
rect 929 1898 985 1932
rect 929 1864 940 1898
rect 974 1864 985 1898
rect 929 1830 985 1864
rect 929 1796 940 1830
rect 974 1796 985 1830
rect 929 1762 985 1796
rect 929 1728 940 1762
rect 974 1728 985 1762
rect 929 1694 985 1728
rect 929 1660 940 1694
rect 974 1660 985 1694
rect 929 1582 985 1660
rect 1035 2170 1088 2182
rect 1035 2136 1046 2170
rect 1080 2136 1088 2170
rect 1035 2102 1088 2136
rect 1035 2068 1046 2102
rect 1080 2068 1088 2102
rect 1035 2034 1088 2068
rect 1035 2000 1046 2034
rect 1080 2000 1088 2034
rect 1035 1966 1088 2000
rect 1035 1932 1046 1966
rect 1080 1932 1088 1966
rect 1035 1898 1088 1932
rect 1035 1864 1046 1898
rect 1080 1864 1088 1898
rect 1035 1830 1088 1864
rect 1035 1796 1046 1830
rect 1080 1796 1088 1830
rect 1035 1762 1088 1796
rect 1035 1728 1046 1762
rect 1080 1728 1088 1762
rect 1035 1694 1088 1728
rect 1035 1660 1046 1694
rect 1080 1660 1088 1694
rect 1035 1582 1088 1660
rect 1148 2170 1201 2182
rect 1148 2136 1156 2170
rect 1190 2136 1201 2170
rect 1148 2102 1201 2136
rect 1148 2068 1156 2102
rect 1190 2068 1201 2102
rect 1148 2034 1201 2068
rect 1148 2000 1156 2034
rect 1190 2000 1201 2034
rect 1148 1966 1201 2000
rect 1148 1932 1156 1966
rect 1190 1932 1201 1966
rect 1148 1898 1201 1932
rect 1148 1864 1156 1898
rect 1190 1864 1201 1898
rect 1148 1830 1201 1864
rect 1148 1796 1156 1830
rect 1190 1796 1201 1830
rect 1148 1762 1201 1796
rect 1148 1728 1156 1762
rect 1190 1728 1201 1762
rect 1148 1694 1201 1728
rect 1148 1660 1156 1694
rect 1190 1660 1201 1694
rect 1148 1582 1201 1660
rect 1251 2170 1307 2182
rect 1251 2136 1262 2170
rect 1296 2136 1307 2170
rect 1251 2102 1307 2136
rect 1251 2068 1262 2102
rect 1296 2068 1307 2102
rect 1251 2034 1307 2068
rect 1251 2000 1262 2034
rect 1296 2000 1307 2034
rect 1251 1966 1307 2000
rect 1251 1932 1262 1966
rect 1296 1932 1307 1966
rect 1251 1898 1307 1932
rect 1251 1864 1262 1898
rect 1296 1864 1307 1898
rect 1251 1830 1307 1864
rect 1251 1796 1262 1830
rect 1296 1796 1307 1830
rect 1251 1762 1307 1796
rect 1251 1728 1262 1762
rect 1296 1728 1307 1762
rect 1251 1694 1307 1728
rect 1251 1660 1262 1694
rect 1296 1660 1307 1694
rect 1251 1582 1307 1660
rect 1357 2170 1410 2182
rect 1357 2136 1368 2170
rect 1402 2136 1410 2170
rect 1357 2102 1410 2136
rect 1357 2068 1368 2102
rect 1402 2068 1410 2102
rect 1357 2034 1410 2068
rect 1357 2000 1368 2034
rect 1402 2000 1410 2034
rect 1357 1966 1410 2000
rect 1357 1932 1368 1966
rect 1402 1932 1410 1966
rect 1357 1898 1410 1932
rect 1357 1864 1368 1898
rect 1402 1864 1410 1898
rect 1357 1830 1410 1864
rect 1357 1796 1368 1830
rect 1402 1796 1410 1830
rect 1357 1762 1410 1796
rect 1357 1728 1368 1762
rect 1402 1728 1410 1762
rect 1357 1694 1410 1728
rect 1357 1660 1368 1694
rect 1402 1660 1410 1694
rect 1357 1582 1410 1660
<< pdiff >>
rect 31 2431 84 2501
rect 31 2397 39 2431
rect 73 2397 84 2431
rect 31 2363 84 2397
rect 31 2329 39 2363
rect 73 2329 84 2363
rect 31 2295 84 2329
rect 31 2261 39 2295
rect 73 2261 84 2295
rect 31 2227 84 2261
rect 31 2193 39 2227
rect 73 2193 84 2227
rect 31 2159 84 2193
rect 31 2125 39 2159
rect 73 2125 84 2159
rect 31 2091 84 2125
rect 31 2057 39 2091
rect 73 2057 84 2091
rect 31 2023 84 2057
rect 31 1989 39 2023
rect 73 1989 84 2023
rect 31 1955 84 1989
rect 31 1921 39 1955
rect 73 1921 84 1955
rect 31 1887 84 1921
rect 31 1853 39 1887
rect 73 1853 84 1887
rect 31 1819 84 1853
rect 31 1785 39 1819
rect 73 1785 84 1819
rect 31 1751 84 1785
rect 31 1717 39 1751
rect 73 1717 84 1751
rect 31 1683 84 1717
rect 31 1649 39 1683
rect 73 1649 84 1683
rect 31 1615 84 1649
rect 31 1581 39 1615
rect 73 1581 84 1615
rect 31 1547 84 1581
rect 31 1513 39 1547
rect 73 1513 84 1547
rect 31 1501 84 1513
rect 134 2431 190 2501
rect 134 2397 145 2431
rect 179 2397 190 2431
rect 134 2363 190 2397
rect 134 2329 145 2363
rect 179 2329 190 2363
rect 134 2295 190 2329
rect 134 2261 145 2295
rect 179 2261 190 2295
rect 134 2227 190 2261
rect 134 2193 145 2227
rect 179 2193 190 2227
rect 134 2159 190 2193
rect 134 2125 145 2159
rect 179 2125 190 2159
rect 134 2091 190 2125
rect 134 2057 145 2091
rect 179 2057 190 2091
rect 134 2023 190 2057
rect 134 1989 145 2023
rect 179 1989 190 2023
rect 134 1955 190 1989
rect 134 1921 145 1955
rect 179 1921 190 1955
rect 134 1887 190 1921
rect 134 1853 145 1887
rect 179 1853 190 1887
rect 134 1819 190 1853
rect 134 1785 145 1819
rect 179 1785 190 1819
rect 134 1751 190 1785
rect 134 1717 145 1751
rect 179 1717 190 1751
rect 134 1683 190 1717
rect 134 1649 145 1683
rect 179 1649 190 1683
rect 134 1615 190 1649
rect 134 1581 145 1615
rect 179 1581 190 1615
rect 134 1547 190 1581
rect 134 1513 145 1547
rect 179 1513 190 1547
rect 134 1501 190 1513
rect 240 2431 293 2501
rect 240 2397 251 2431
rect 285 2397 293 2431
rect 240 2363 293 2397
rect 240 2329 251 2363
rect 285 2329 293 2363
rect 240 2295 293 2329
rect 240 2261 251 2295
rect 285 2261 293 2295
rect 240 2227 293 2261
rect 240 2193 251 2227
rect 285 2193 293 2227
rect 240 2159 293 2193
rect 240 2125 251 2159
rect 285 2125 293 2159
rect 240 2091 293 2125
rect 240 2057 251 2091
rect 285 2057 293 2091
rect 240 2023 293 2057
rect 240 1989 251 2023
rect 285 1989 293 2023
rect 240 1955 293 1989
rect 240 1921 251 1955
rect 285 1921 293 1955
rect 240 1887 293 1921
rect 240 1853 251 1887
rect 285 1853 293 1887
rect 240 1819 293 1853
rect 240 1785 251 1819
rect 285 1785 293 1819
rect 240 1751 293 1785
rect 240 1717 251 1751
rect 285 1717 293 1751
rect 240 1683 293 1717
rect 240 1649 251 1683
rect 285 1649 293 1683
rect 240 1615 293 1649
rect 240 1581 251 1615
rect 285 1581 293 1615
rect 240 1547 293 1581
rect 240 1513 251 1547
rect 285 1513 293 1547
rect 240 1501 293 1513
rect 354 2431 407 2501
rect 354 2397 362 2431
rect 396 2397 407 2431
rect 354 2363 407 2397
rect 354 2329 362 2363
rect 396 2329 407 2363
rect 354 2295 407 2329
rect 354 2261 362 2295
rect 396 2261 407 2295
rect 354 2227 407 2261
rect 354 2193 362 2227
rect 396 2193 407 2227
rect 354 2159 407 2193
rect 354 2125 362 2159
rect 396 2125 407 2159
rect 354 2091 407 2125
rect 354 2057 362 2091
rect 396 2057 407 2091
rect 354 2023 407 2057
rect 354 1989 362 2023
rect 396 1989 407 2023
rect 354 1955 407 1989
rect 354 1921 362 1955
rect 396 1921 407 1955
rect 354 1887 407 1921
rect 354 1853 362 1887
rect 396 1853 407 1887
rect 354 1819 407 1853
rect 354 1785 362 1819
rect 396 1785 407 1819
rect 354 1751 407 1785
rect 354 1717 362 1751
rect 396 1717 407 1751
rect 354 1683 407 1717
rect 354 1649 362 1683
rect 396 1649 407 1683
rect 354 1615 407 1649
rect 354 1581 362 1615
rect 396 1581 407 1615
rect 354 1547 407 1581
rect 354 1513 362 1547
rect 396 1513 407 1547
rect 354 1501 407 1513
rect 457 2431 513 2501
rect 457 2397 468 2431
rect 502 2397 513 2431
rect 457 2363 513 2397
rect 457 2329 468 2363
rect 502 2329 513 2363
rect 457 2295 513 2329
rect 457 2261 468 2295
rect 502 2261 513 2295
rect 457 2227 513 2261
rect 457 2193 468 2227
rect 502 2193 513 2227
rect 457 2159 513 2193
rect 457 2125 468 2159
rect 502 2125 513 2159
rect 457 2091 513 2125
rect 457 2057 468 2091
rect 502 2057 513 2091
rect 457 2023 513 2057
rect 457 1989 468 2023
rect 502 1989 513 2023
rect 457 1955 513 1989
rect 457 1921 468 1955
rect 502 1921 513 1955
rect 457 1887 513 1921
rect 457 1853 468 1887
rect 502 1853 513 1887
rect 457 1819 513 1853
rect 457 1785 468 1819
rect 502 1785 513 1819
rect 457 1751 513 1785
rect 457 1717 468 1751
rect 502 1717 513 1751
rect 457 1683 513 1717
rect 457 1649 468 1683
rect 502 1649 513 1683
rect 457 1615 513 1649
rect 457 1581 468 1615
rect 502 1581 513 1615
rect 457 1547 513 1581
rect 457 1513 468 1547
rect 502 1513 513 1547
rect 457 1501 513 1513
rect 563 2431 616 2501
rect 563 2397 574 2431
rect 608 2397 616 2431
rect 563 2363 616 2397
rect 563 2329 574 2363
rect 608 2329 616 2363
rect 563 2295 616 2329
rect 563 2261 574 2295
rect 608 2261 616 2295
rect 563 2227 616 2261
rect 563 2193 574 2227
rect 608 2193 616 2227
rect 563 2159 616 2193
rect 563 2125 574 2159
rect 608 2125 616 2159
rect 563 2091 616 2125
rect 563 2057 574 2091
rect 608 2057 616 2091
rect 563 2023 616 2057
rect 563 1989 574 2023
rect 608 1989 616 2023
rect 563 1955 616 1989
rect 563 1921 574 1955
rect 608 1921 616 1955
rect 563 1887 616 1921
rect 563 1853 574 1887
rect 608 1853 616 1887
rect 563 1819 616 1853
rect 563 1785 574 1819
rect 608 1785 616 1819
rect 563 1751 616 1785
rect 563 1717 574 1751
rect 608 1717 616 1751
rect 563 1683 616 1717
rect 563 1649 574 1683
rect 608 1649 616 1683
rect 563 1615 616 1649
rect 563 1581 574 1615
rect 608 1581 616 1615
rect 563 1547 616 1581
rect 563 1513 574 1547
rect 608 1513 616 1547
rect 563 1501 616 1513
<< mvndiff >>
rect 861 1053 914 1123
rect 861 1019 869 1053
rect 903 1019 914 1053
rect 861 985 914 1019
rect 861 951 869 985
rect 903 951 914 985
rect 861 917 914 951
rect 861 883 869 917
rect 903 883 914 917
rect 861 849 914 883
rect 861 815 869 849
rect 903 815 914 849
rect 861 781 914 815
rect 861 747 869 781
rect 903 747 914 781
rect 861 713 914 747
rect 861 679 869 713
rect 903 679 914 713
rect 861 645 914 679
rect 861 611 869 645
rect 903 611 914 645
rect 861 577 914 611
rect 861 543 869 577
rect 903 543 914 577
rect 861 509 914 543
rect 861 475 869 509
rect 903 475 914 509
rect 861 441 914 475
rect 861 407 869 441
rect 903 407 914 441
rect 861 373 914 407
rect 861 339 869 373
rect 903 339 914 373
rect 861 305 914 339
rect 861 271 869 305
rect 903 271 914 305
rect 861 237 914 271
rect 861 203 869 237
rect 903 203 914 237
rect 861 169 914 203
rect 861 135 869 169
rect 903 135 914 169
rect 861 123 914 135
rect 1014 1053 1070 1123
rect 1014 1019 1025 1053
rect 1059 1019 1070 1053
rect 1014 985 1070 1019
rect 1014 951 1025 985
rect 1059 951 1070 985
rect 1014 917 1070 951
rect 1014 883 1025 917
rect 1059 883 1070 917
rect 1014 849 1070 883
rect 1014 815 1025 849
rect 1059 815 1070 849
rect 1014 781 1070 815
rect 1014 747 1025 781
rect 1059 747 1070 781
rect 1014 713 1070 747
rect 1014 679 1025 713
rect 1059 679 1070 713
rect 1014 645 1070 679
rect 1014 611 1025 645
rect 1059 611 1070 645
rect 1014 577 1070 611
rect 1014 543 1025 577
rect 1059 543 1070 577
rect 1014 509 1070 543
rect 1014 475 1025 509
rect 1059 475 1070 509
rect 1014 441 1070 475
rect 1014 407 1025 441
rect 1059 407 1070 441
rect 1014 373 1070 407
rect 1014 339 1025 373
rect 1059 339 1070 373
rect 1014 305 1070 339
rect 1014 271 1025 305
rect 1059 271 1070 305
rect 1014 237 1070 271
rect 1014 203 1025 237
rect 1059 203 1070 237
rect 1014 169 1070 203
rect 1014 135 1025 169
rect 1059 135 1070 169
rect 1014 123 1070 135
rect 1170 1053 1223 1123
rect 1170 1019 1181 1053
rect 1215 1019 1223 1053
rect 1170 985 1223 1019
rect 1170 951 1181 985
rect 1215 951 1223 985
rect 1170 917 1223 951
rect 1170 883 1181 917
rect 1215 883 1223 917
rect 1170 849 1223 883
rect 1170 815 1181 849
rect 1215 815 1223 849
rect 1170 781 1223 815
rect 1170 747 1181 781
rect 1215 747 1223 781
rect 1170 713 1223 747
rect 1170 679 1181 713
rect 1215 679 1223 713
rect 1170 645 1223 679
rect 1170 611 1181 645
rect 1215 611 1223 645
rect 1170 577 1223 611
rect 1170 543 1181 577
rect 1215 543 1223 577
rect 1170 509 1223 543
rect 1170 475 1181 509
rect 1215 475 1223 509
rect 1170 441 1223 475
rect 1170 407 1181 441
rect 1215 407 1223 441
rect 1170 373 1223 407
rect 1170 339 1181 373
rect 1215 339 1223 373
rect 1170 305 1223 339
rect 1170 271 1181 305
rect 1215 271 1223 305
rect 1170 237 1223 271
rect 1170 203 1181 237
rect 1215 203 1223 237
rect 1170 169 1223 203
rect 1170 135 1181 169
rect 1215 135 1223 169
rect 1170 123 1223 135
<< mvpdiff >>
rect 59 1053 112 1123
rect 59 1019 67 1053
rect 101 1019 112 1053
rect 59 985 112 1019
rect 59 951 67 985
rect 101 951 112 985
rect 59 917 112 951
rect 59 883 67 917
rect 101 883 112 917
rect 59 849 112 883
rect 59 815 67 849
rect 101 815 112 849
rect 59 781 112 815
rect 59 747 67 781
rect 101 747 112 781
rect 59 713 112 747
rect 59 679 67 713
rect 101 679 112 713
rect 59 645 112 679
rect 59 611 67 645
rect 101 611 112 645
rect 59 577 112 611
rect 59 543 67 577
rect 101 543 112 577
rect 59 509 112 543
rect 59 475 67 509
rect 101 475 112 509
rect 59 441 112 475
rect 59 407 67 441
rect 101 407 112 441
rect 59 373 112 407
rect 59 339 67 373
rect 101 339 112 373
rect 59 305 112 339
rect 59 271 67 305
rect 101 271 112 305
rect 59 237 112 271
rect 59 203 67 237
rect 101 203 112 237
rect 59 169 112 203
rect 59 135 67 169
rect 101 135 112 169
rect 59 123 112 135
rect 212 1053 268 1123
rect 212 1019 223 1053
rect 257 1019 268 1053
rect 212 985 268 1019
rect 212 951 223 985
rect 257 951 268 985
rect 212 917 268 951
rect 212 883 223 917
rect 257 883 268 917
rect 212 849 268 883
rect 212 815 223 849
rect 257 815 268 849
rect 212 781 268 815
rect 212 747 223 781
rect 257 747 268 781
rect 212 713 268 747
rect 212 679 223 713
rect 257 679 268 713
rect 212 645 268 679
rect 212 611 223 645
rect 257 611 268 645
rect 212 577 268 611
rect 212 543 223 577
rect 257 543 268 577
rect 212 509 268 543
rect 212 475 223 509
rect 257 475 268 509
rect 212 441 268 475
rect 212 407 223 441
rect 257 407 268 441
rect 212 373 268 407
rect 212 339 223 373
rect 257 339 268 373
rect 212 305 268 339
rect 212 271 223 305
rect 257 271 268 305
rect 212 237 268 271
rect 212 203 223 237
rect 257 203 268 237
rect 212 169 268 203
rect 212 135 223 169
rect 257 135 268 169
rect 212 123 268 135
rect 368 1053 424 1123
rect 368 1019 379 1053
rect 413 1019 424 1053
rect 368 985 424 1019
rect 368 951 379 985
rect 413 951 424 985
rect 368 917 424 951
rect 368 883 379 917
rect 413 883 424 917
rect 368 849 424 883
rect 368 815 379 849
rect 413 815 424 849
rect 368 781 424 815
rect 368 747 379 781
rect 413 747 424 781
rect 368 713 424 747
rect 368 679 379 713
rect 413 679 424 713
rect 368 645 424 679
rect 368 611 379 645
rect 413 611 424 645
rect 368 577 424 611
rect 368 543 379 577
rect 413 543 424 577
rect 368 509 424 543
rect 368 475 379 509
rect 413 475 424 509
rect 368 441 424 475
rect 368 407 379 441
rect 413 407 424 441
rect 368 373 424 407
rect 368 339 379 373
rect 413 339 424 373
rect 368 305 424 339
rect 368 271 379 305
rect 413 271 424 305
rect 368 237 424 271
rect 368 203 379 237
rect 413 203 424 237
rect 368 169 424 203
rect 368 135 379 169
rect 413 135 424 169
rect 368 123 424 135
rect 524 1053 577 1123
rect 524 1019 535 1053
rect 569 1019 577 1053
rect 524 985 577 1019
rect 524 951 535 985
rect 569 951 577 985
rect 524 917 577 951
rect 524 883 535 917
rect 569 883 577 917
rect 524 849 577 883
rect 524 815 535 849
rect 569 815 577 849
rect 524 781 577 815
rect 524 747 535 781
rect 569 747 577 781
rect 524 713 577 747
rect 524 679 535 713
rect 569 679 577 713
rect 524 645 577 679
rect 524 611 535 645
rect 569 611 577 645
rect 524 577 577 611
rect 524 543 535 577
rect 569 543 577 577
rect 524 509 577 543
rect 524 475 535 509
rect 569 475 577 509
rect 524 441 577 475
rect 524 407 535 441
rect 569 407 577 441
rect 524 373 577 407
rect 524 339 535 373
rect 569 339 577 373
rect 524 305 577 339
rect 524 271 535 305
rect 569 271 577 305
rect 524 237 577 271
rect 524 203 535 237
rect 569 203 577 237
rect 524 169 577 203
rect 524 135 535 169
rect 569 135 577 169
rect 524 123 577 135
<< ndiffc >>
rect 834 2136 868 2170
rect 834 2068 868 2102
rect 834 2000 868 2034
rect 834 1932 868 1966
rect 834 1864 868 1898
rect 834 1796 868 1830
rect 834 1728 868 1762
rect 834 1660 868 1694
rect 940 2136 974 2170
rect 940 2068 974 2102
rect 940 2000 974 2034
rect 940 1932 974 1966
rect 940 1864 974 1898
rect 940 1796 974 1830
rect 940 1728 974 1762
rect 940 1660 974 1694
rect 1046 2136 1080 2170
rect 1046 2068 1080 2102
rect 1046 2000 1080 2034
rect 1046 1932 1080 1966
rect 1046 1864 1080 1898
rect 1046 1796 1080 1830
rect 1046 1728 1080 1762
rect 1046 1660 1080 1694
rect 1156 2136 1190 2170
rect 1156 2068 1190 2102
rect 1156 2000 1190 2034
rect 1156 1932 1190 1966
rect 1156 1864 1190 1898
rect 1156 1796 1190 1830
rect 1156 1728 1190 1762
rect 1156 1660 1190 1694
rect 1262 2136 1296 2170
rect 1262 2068 1296 2102
rect 1262 2000 1296 2034
rect 1262 1932 1296 1966
rect 1262 1864 1296 1898
rect 1262 1796 1296 1830
rect 1262 1728 1296 1762
rect 1262 1660 1296 1694
rect 1368 2136 1402 2170
rect 1368 2068 1402 2102
rect 1368 2000 1402 2034
rect 1368 1932 1402 1966
rect 1368 1864 1402 1898
rect 1368 1796 1402 1830
rect 1368 1728 1402 1762
rect 1368 1660 1402 1694
<< pdiffc >>
rect 39 2397 73 2431
rect 39 2329 73 2363
rect 39 2261 73 2295
rect 39 2193 73 2227
rect 39 2125 73 2159
rect 39 2057 73 2091
rect 39 1989 73 2023
rect 39 1921 73 1955
rect 39 1853 73 1887
rect 39 1785 73 1819
rect 39 1717 73 1751
rect 39 1649 73 1683
rect 39 1581 73 1615
rect 39 1513 73 1547
rect 145 2397 179 2431
rect 145 2329 179 2363
rect 145 2261 179 2295
rect 145 2193 179 2227
rect 145 2125 179 2159
rect 145 2057 179 2091
rect 145 1989 179 2023
rect 145 1921 179 1955
rect 145 1853 179 1887
rect 145 1785 179 1819
rect 145 1717 179 1751
rect 145 1649 179 1683
rect 145 1581 179 1615
rect 145 1513 179 1547
rect 251 2397 285 2431
rect 251 2329 285 2363
rect 251 2261 285 2295
rect 251 2193 285 2227
rect 251 2125 285 2159
rect 251 2057 285 2091
rect 251 1989 285 2023
rect 251 1921 285 1955
rect 251 1853 285 1887
rect 251 1785 285 1819
rect 251 1717 285 1751
rect 251 1649 285 1683
rect 251 1581 285 1615
rect 251 1513 285 1547
rect 362 2397 396 2431
rect 362 2329 396 2363
rect 362 2261 396 2295
rect 362 2193 396 2227
rect 362 2125 396 2159
rect 362 2057 396 2091
rect 362 1989 396 2023
rect 362 1921 396 1955
rect 362 1853 396 1887
rect 362 1785 396 1819
rect 362 1717 396 1751
rect 362 1649 396 1683
rect 362 1581 396 1615
rect 362 1513 396 1547
rect 468 2397 502 2431
rect 468 2329 502 2363
rect 468 2261 502 2295
rect 468 2193 502 2227
rect 468 2125 502 2159
rect 468 2057 502 2091
rect 468 1989 502 2023
rect 468 1921 502 1955
rect 468 1853 502 1887
rect 468 1785 502 1819
rect 468 1717 502 1751
rect 468 1649 502 1683
rect 468 1581 502 1615
rect 468 1513 502 1547
rect 574 2397 608 2431
rect 574 2329 608 2363
rect 574 2261 608 2295
rect 574 2193 608 2227
rect 574 2125 608 2159
rect 574 2057 608 2091
rect 574 1989 608 2023
rect 574 1921 608 1955
rect 574 1853 608 1887
rect 574 1785 608 1819
rect 574 1717 608 1751
rect 574 1649 608 1683
rect 574 1581 608 1615
rect 574 1513 608 1547
<< mvndiffc >>
rect 869 1019 903 1053
rect 869 951 903 985
rect 869 883 903 917
rect 869 815 903 849
rect 869 747 903 781
rect 869 679 903 713
rect 869 611 903 645
rect 869 543 903 577
rect 869 475 903 509
rect 869 407 903 441
rect 869 339 903 373
rect 869 271 903 305
rect 869 203 903 237
rect 869 135 903 169
rect 1025 1019 1059 1053
rect 1025 951 1059 985
rect 1025 883 1059 917
rect 1025 815 1059 849
rect 1025 747 1059 781
rect 1025 679 1059 713
rect 1025 611 1059 645
rect 1025 543 1059 577
rect 1025 475 1059 509
rect 1025 407 1059 441
rect 1025 339 1059 373
rect 1025 271 1059 305
rect 1025 203 1059 237
rect 1025 135 1059 169
rect 1181 1019 1215 1053
rect 1181 951 1215 985
rect 1181 883 1215 917
rect 1181 815 1215 849
rect 1181 747 1215 781
rect 1181 679 1215 713
rect 1181 611 1215 645
rect 1181 543 1215 577
rect 1181 475 1215 509
rect 1181 407 1215 441
rect 1181 339 1215 373
rect 1181 271 1215 305
rect 1181 203 1215 237
rect 1181 135 1215 169
<< mvpdiffc >>
rect 67 1019 101 1053
rect 67 951 101 985
rect 67 883 101 917
rect 67 815 101 849
rect 67 747 101 781
rect 67 679 101 713
rect 67 611 101 645
rect 67 543 101 577
rect 67 475 101 509
rect 67 407 101 441
rect 67 339 101 373
rect 67 271 101 305
rect 67 203 101 237
rect 67 135 101 169
rect 223 1019 257 1053
rect 223 951 257 985
rect 223 883 257 917
rect 223 815 257 849
rect 223 747 257 781
rect 223 679 257 713
rect 223 611 257 645
rect 223 543 257 577
rect 223 475 257 509
rect 223 407 257 441
rect 223 339 257 373
rect 223 271 257 305
rect 223 203 257 237
rect 223 135 257 169
rect 379 1019 413 1053
rect 379 951 413 985
rect 379 883 413 917
rect 379 815 413 849
rect 379 747 413 781
rect 379 679 413 713
rect 379 611 413 645
rect 379 543 413 577
rect 379 475 413 509
rect 379 407 413 441
rect 379 339 413 373
rect 379 271 413 305
rect 379 203 413 237
rect 379 135 413 169
rect 535 1019 569 1053
rect 535 951 569 985
rect 535 883 569 917
rect 535 815 569 849
rect 535 747 569 781
rect 535 679 569 713
rect 535 611 569 645
rect 535 543 569 577
rect 535 475 569 509
rect 535 407 569 441
rect 535 339 569 373
rect 535 271 569 305
rect 535 203 569 237
rect 535 135 569 169
<< nsubdiff >>
rect 67 2575 101 2609
rect 135 2575 169 2609
rect 203 2575 237 2609
rect 271 2575 305 2609
rect 339 2575 373 2609
rect 407 2575 441 2609
rect 475 2575 509 2609
rect 543 2575 603 2609
<< mvpsubdiff >>
rect 1305 1082 1339 1116
rect 1305 971 1339 1048
rect 1305 859 1339 937
rect 1305 747 1339 825
rect 1305 635 1339 713
rect 1305 523 1339 601
rect 1305 411 1339 489
rect 1305 299 1339 377
rect 1305 187 1339 265
rect 1305 119 1339 153
<< mvnsubdiff >>
rect 59 15 83 49
rect 117 15 171 49
rect 205 15 258 49
rect 292 15 345 49
rect 379 15 432 49
rect 466 15 519 49
rect 553 15 577 49
<< nsubdiffcont >>
rect 101 2575 135 2609
rect 169 2575 203 2609
rect 237 2575 271 2609
rect 305 2575 339 2609
rect 373 2575 407 2609
rect 441 2575 475 2609
rect 509 2575 543 2609
<< mvpsubdiffcont >>
rect 1305 1048 1339 1082
rect 1305 937 1339 971
rect 1305 825 1339 859
rect 1305 713 1339 747
rect 1305 601 1339 635
rect 1305 489 1339 523
rect 1305 377 1339 411
rect 1305 265 1339 299
rect 1305 153 1339 187
<< mvnsubdiffcont >>
rect 83 15 117 49
rect 171 15 205 49
rect 258 15 292 49
rect 345 15 379 49
rect 432 15 466 49
rect 519 15 553 49
<< poly >>
rect 84 2501 134 2533
rect 190 2501 240 2533
rect 407 2501 457 2533
rect 513 2501 563 2533
rect 879 2182 929 2214
rect 985 2182 1035 2214
rect 1201 2182 1251 2214
rect 1307 2182 1357 2214
rect 879 1550 929 1582
rect 863 1534 929 1550
rect 84 1469 134 1501
rect 190 1469 240 1501
rect 84 1453 240 1469
rect 407 1460 457 1501
rect 513 1460 563 1501
rect 863 1500 879 1534
rect 913 1500 929 1534
rect 84 1419 100 1453
rect 134 1419 190 1453
rect 224 1419 240 1453
rect 84 1403 240 1419
rect 398 1444 464 1460
rect 398 1410 414 1444
rect 448 1410 464 1444
rect 398 1354 464 1410
rect 398 1320 414 1354
rect 448 1320 464 1354
rect 398 1304 464 1320
rect 513 1444 579 1460
rect 513 1410 529 1444
rect 563 1410 579 1444
rect 513 1354 579 1410
rect 863 1444 929 1500
rect 863 1410 879 1444
rect 913 1410 929 1444
rect 863 1394 929 1410
rect 985 1550 1035 1582
rect 1201 1550 1251 1582
rect 1307 1550 1357 1582
rect 985 1534 1051 1550
rect 985 1500 1001 1534
rect 1035 1500 1051 1534
rect 985 1444 1051 1500
rect 1201 1534 1357 1550
rect 1201 1500 1217 1534
rect 1251 1500 1307 1534
rect 1341 1500 1357 1534
rect 1201 1484 1357 1500
rect 985 1410 1001 1444
rect 1035 1410 1051 1444
rect 985 1394 1051 1410
rect 513 1320 529 1354
rect 563 1320 579 1354
rect 513 1304 579 1320
rect 914 1273 1014 1289
rect 914 1239 946 1273
rect 980 1239 1014 1273
rect 75 1205 212 1221
rect 75 1171 91 1205
rect 125 1171 162 1205
rect 196 1171 212 1205
rect 75 1155 212 1171
rect 112 1123 212 1155
rect 268 1205 524 1221
rect 268 1171 284 1205
rect 318 1171 379 1205
rect 413 1171 474 1205
rect 508 1171 524 1205
rect 268 1155 524 1171
rect 268 1123 368 1155
rect 424 1123 524 1155
rect 914 1205 1014 1239
rect 914 1171 946 1205
rect 980 1171 1014 1205
rect 914 1123 1014 1171
rect 1070 1273 1170 1289
rect 1070 1239 1102 1273
rect 1136 1239 1170 1273
rect 1070 1205 1170 1239
rect 1070 1171 1102 1205
rect 1136 1171 1170 1205
rect 1070 1123 1170 1171
rect 112 91 212 123
rect 268 91 368 123
rect 424 91 524 123
rect 914 91 1014 123
rect 1070 91 1170 123
<< polycont >>
rect 879 1500 913 1534
rect 100 1419 134 1453
rect 190 1419 224 1453
rect 414 1410 448 1444
rect 414 1320 448 1354
rect 529 1410 563 1444
rect 879 1410 913 1444
rect 1001 1500 1035 1534
rect 1217 1500 1251 1534
rect 1307 1500 1341 1534
rect 1001 1410 1035 1444
rect 529 1320 563 1354
rect 946 1239 980 1273
rect 91 1171 125 1205
rect 162 1171 196 1205
rect 284 1171 318 1205
rect 379 1171 413 1205
rect 474 1171 508 1205
rect 946 1171 980 1205
rect 1102 1239 1136 1273
rect 1102 1171 1136 1205
<< locali >>
rect 135 2575 149 2609
rect 203 2575 231 2609
rect 271 2575 305 2609
rect 347 2575 373 2609
rect 429 2575 441 2609
rect 475 2575 476 2609
rect 543 2575 557 2609
rect 591 2575 603 2609
rect 39 2431 73 2455
rect 39 2363 73 2381
rect 39 2295 73 2307
rect 39 2227 73 2233
rect 39 2119 73 2125
rect 39 2045 73 2057
rect 39 1971 73 1989
rect 39 1898 73 1921
rect 39 1825 73 1853
rect 39 1752 73 1785
rect 39 1683 73 1717
rect 39 1615 73 1645
rect 39 1547 73 1581
rect 39 1497 73 1513
rect 145 2435 179 2447
rect 145 2363 179 2397
rect 145 2295 179 2326
rect 145 2227 179 2251
rect 145 2159 179 2176
rect 145 2091 179 2101
rect 145 2023 179 2026
rect 145 1985 179 1989
rect 145 1910 179 1921
rect 145 1835 179 1853
rect 145 1759 179 1785
rect 145 1683 179 1717
rect 145 1615 179 1649
rect 145 1547 179 1581
rect 145 1497 179 1513
rect 251 2431 285 2455
rect 251 2363 285 2381
rect 251 2295 285 2307
rect 251 2227 285 2233
rect 251 2119 285 2125
rect 251 2045 285 2057
rect 251 1971 285 1989
rect 251 1898 285 1921
rect 251 1825 285 1853
rect 251 1752 285 1785
rect 251 1683 285 1717
rect 251 1615 285 1645
rect 251 1547 285 1581
rect 251 1497 285 1513
rect 362 2435 396 2447
rect 362 2363 396 2397
rect 362 2295 396 2326
rect 362 2227 396 2251
rect 362 2159 396 2176
rect 362 2091 396 2101
rect 362 2023 396 2026
rect 362 1985 396 1989
rect 362 1910 396 1921
rect 362 1835 396 1853
rect 362 1760 396 1785
rect 362 1685 396 1717
rect 362 1615 396 1649
rect 362 1547 396 1581
rect 362 1497 396 1513
rect 468 2431 502 2455
rect 468 2363 502 2381
rect 468 2295 502 2307
rect 468 2227 502 2233
rect 468 2119 502 2125
rect 468 2045 502 2057
rect 468 1971 502 1989
rect 468 1898 502 1921
rect 468 1825 502 1853
rect 468 1752 502 1785
rect 468 1683 502 1717
rect 468 1615 502 1645
rect 468 1547 502 1581
rect 468 1497 502 1513
rect 574 2435 608 2447
rect 574 2363 608 2397
rect 574 2295 608 2326
rect 574 2227 608 2251
rect 574 2159 608 2176
rect 574 2091 608 2101
rect 574 2023 608 2026
rect 574 1984 608 1989
rect 574 1908 608 1921
rect 574 1832 608 1853
rect 574 1756 608 1785
rect 574 1683 608 1717
rect 574 1615 608 1646
rect 834 2174 868 2186
rect 834 2102 868 2136
rect 834 2034 868 2060
rect 834 1966 868 1980
rect 834 1898 868 1900
rect 834 1853 868 1864
rect 834 1772 868 1796
rect 834 1694 868 1728
rect 834 1644 868 1657
rect 940 2174 974 2186
rect 940 2102 974 2136
rect 940 2034 974 2060
rect 940 1966 974 1980
rect 940 1898 974 1900
rect 940 1853 974 1864
rect 940 1772 974 1796
rect 940 1694 974 1728
rect 940 1644 974 1657
rect 1046 2174 1080 2186
rect 1046 2102 1080 2136
rect 1046 2034 1080 2060
rect 1046 1966 1080 1980
rect 1046 1898 1080 1900
rect 1046 1853 1080 1864
rect 1046 1772 1080 1796
rect 1046 1694 1080 1728
rect 1046 1644 1080 1657
rect 1156 2174 1190 2186
rect 1156 2102 1190 2136
rect 1156 2034 1190 2060
rect 1156 1966 1190 1980
rect 1156 1898 1190 1900
rect 1156 1853 1190 1864
rect 1156 1772 1190 1796
rect 1156 1694 1190 1728
rect 1156 1644 1190 1657
rect 1262 2174 1296 2186
rect 1262 2102 1296 2136
rect 1262 2034 1296 2060
rect 1262 1966 1296 1980
rect 1262 1898 1296 1900
rect 1262 1853 1296 1864
rect 1262 1772 1296 1796
rect 1262 1694 1296 1728
rect 1262 1644 1296 1657
rect 1368 2174 1402 2186
rect 1368 2102 1402 2136
rect 1368 2034 1402 2060
rect 1368 1966 1402 1980
rect 1368 1898 1402 1900
rect 1368 1853 1402 1864
rect 1368 1772 1402 1796
rect 1368 1694 1402 1728
rect 1368 1644 1402 1657
rect 574 1547 608 1581
rect 574 1497 608 1513
rect 879 1534 913 1550
rect 414 1457 448 1460
rect 84 1419 97 1453
rect 134 1419 190 1453
rect 228 1419 240 1453
rect 414 1385 448 1410
rect 414 1304 448 1320
rect 529 1457 563 1460
rect 529 1385 563 1410
rect 879 1444 913 1476
rect 879 1394 913 1404
rect 1001 1538 1035 1550
rect 1201 1500 1213 1534
rect 1251 1500 1297 1534
rect 1341 1500 1357 1534
rect 1001 1466 1035 1500
rect 1001 1394 1035 1410
rect 529 1304 563 1320
rect 1272 1387 1370 1421
rect 1238 1339 1404 1387
rect 1272 1305 1370 1339
rect 946 1274 980 1289
rect 1102 1274 1136 1289
rect 946 1273 949 1274
rect 980 1239 983 1240
rect 946 1205 983 1239
rect 75 1171 87 1205
rect 125 1171 162 1205
rect 200 1171 212 1205
rect 268 1171 280 1205
rect 318 1171 379 1205
rect 413 1171 474 1205
rect 512 1171 524 1205
rect 980 1202 983 1205
rect 946 1168 949 1171
rect 1102 1205 1136 1239
rect 946 1155 980 1168
rect 1102 1155 1136 1168
rect 1238 1257 1404 1305
rect 1272 1223 1370 1257
rect 1238 1175 1404 1223
rect 1272 1141 1370 1175
rect 1238 1092 1404 1141
rect 1238 1069 1305 1092
rect 67 1053 101 1069
rect 67 941 101 951
rect 67 863 101 883
rect 67 785 101 815
rect 67 713 101 747
rect 67 645 101 673
rect 67 577 101 595
rect 67 509 101 517
rect 67 473 101 475
rect 67 396 101 407
rect 67 319 101 339
rect 67 242 101 271
rect 67 169 101 203
rect 67 119 101 131
rect 223 1053 257 1069
rect 223 941 257 951
rect 223 863 257 883
rect 223 785 257 815
rect 223 713 257 747
rect 223 645 257 673
rect 223 577 257 595
rect 223 509 257 517
rect 223 473 257 475
rect 223 396 257 407
rect 223 319 257 339
rect 223 242 257 271
rect 223 169 257 203
rect 223 119 257 131
rect 379 1053 413 1069
rect 379 941 413 951
rect 379 863 413 883
rect 379 785 413 815
rect 379 713 413 747
rect 379 645 413 673
rect 379 577 413 595
rect 379 509 413 517
rect 379 473 413 475
rect 379 396 413 407
rect 379 319 413 339
rect 379 242 413 271
rect 379 169 413 203
rect 379 119 413 131
rect 535 1053 569 1069
rect 535 941 569 951
rect 535 863 569 883
rect 535 785 569 815
rect 535 713 569 747
rect 535 645 569 673
rect 535 577 569 595
rect 535 509 569 517
rect 535 473 569 475
rect 535 396 569 407
rect 535 319 569 339
rect 535 242 569 271
rect 535 169 569 203
rect 535 119 569 131
rect 869 1053 903 1069
rect 869 941 903 951
rect 869 863 903 883
rect 869 785 903 815
rect 869 713 903 747
rect 869 645 903 673
rect 869 577 903 595
rect 869 509 903 517
rect 869 473 903 475
rect 869 396 903 407
rect 869 319 903 339
rect 869 242 903 271
rect 869 169 903 203
rect 869 119 903 131
rect 1025 1053 1059 1069
rect 1025 941 1059 951
rect 1025 863 1059 883
rect 1025 785 1059 815
rect 1025 713 1059 747
rect 1025 645 1059 673
rect 1025 577 1059 595
rect 1025 509 1059 517
rect 1025 473 1059 475
rect 1025 396 1059 407
rect 1025 319 1059 339
rect 1025 242 1059 271
rect 1025 169 1059 203
rect 1025 119 1059 131
rect 1181 1053 1305 1069
rect 1215 1048 1305 1053
rect 1339 1048 1404 1092
rect 1215 1015 1404 1048
rect 1215 981 1305 1015
rect 1339 981 1404 1015
rect 1215 971 1404 981
rect 1215 951 1305 971
rect 1181 941 1305 951
rect 1215 904 1305 941
rect 1339 904 1404 971
rect 1215 883 1404 904
rect 1181 863 1404 883
rect 1215 861 1404 863
rect 1215 825 1305 861
rect 1339 825 1404 861
rect 1215 815 1404 825
rect 1181 785 1404 815
rect 1215 784 1404 785
rect 1215 750 1305 784
rect 1339 750 1404 784
rect 1215 747 1404 750
rect 1181 713 1305 747
rect 1339 713 1404 747
rect 1215 707 1404 713
rect 1215 673 1305 707
rect 1339 673 1404 707
rect 1181 645 1404 673
rect 1215 635 1404 645
rect 1215 596 1305 635
rect 1339 596 1404 635
rect 1215 595 1404 596
rect 1181 577 1404 595
rect 1215 553 1404 577
rect 1215 517 1305 553
rect 1181 509 1305 517
rect 1215 489 1305 509
rect 1339 489 1404 553
rect 1215 476 1404 489
rect 1215 475 1305 476
rect 1181 473 1305 475
rect 1215 442 1305 473
rect 1339 442 1404 476
rect 1215 411 1404 442
rect 1215 407 1305 411
rect 1181 396 1305 407
rect 1215 365 1305 396
rect 1339 365 1404 411
rect 1215 339 1404 365
rect 1181 321 1404 339
rect 1181 319 1305 321
rect 1215 271 1305 319
rect 1181 265 1305 271
rect 1339 265 1404 321
rect 1181 243 1404 265
rect 1181 242 1305 243
rect 1215 209 1305 242
rect 1339 209 1404 243
rect 1215 203 1404 209
rect 1181 187 1404 203
rect 1181 169 1305 187
rect 1215 131 1305 169
rect 1339 131 1404 187
rect 1181 119 1404 131
rect 117 15 141 49
rect 205 15 224 49
rect 292 15 307 49
rect 341 15 345 49
rect 379 15 390 49
rect 424 15 432 49
rect 466 15 473 49
rect 507 15 519 49
rect 553 15 556 49
<< viali >>
rect 67 2575 101 2609
rect 149 2575 169 2609
rect 169 2575 183 2609
rect 231 2575 237 2609
rect 237 2575 265 2609
rect 313 2575 339 2609
rect 339 2575 347 2609
rect 395 2575 407 2609
rect 407 2575 429 2609
rect 476 2575 509 2609
rect 509 2575 510 2609
rect 557 2575 591 2609
rect 39 2455 73 2489
rect 251 2455 285 2489
rect 39 2397 73 2415
rect 39 2381 73 2397
rect 39 2329 73 2341
rect 39 2307 73 2329
rect 39 2261 73 2267
rect 39 2233 73 2261
rect 39 2159 73 2193
rect 39 2091 73 2119
rect 39 2085 73 2091
rect 39 2023 73 2045
rect 39 2011 73 2023
rect 39 1955 73 1971
rect 39 1937 73 1955
rect 39 1887 73 1898
rect 39 1864 73 1887
rect 39 1819 73 1825
rect 39 1791 73 1819
rect 39 1751 73 1752
rect 39 1718 73 1751
rect 39 1649 73 1679
rect 39 1645 73 1649
rect 145 2431 179 2435
rect 145 2401 179 2431
rect 145 2329 179 2360
rect 145 2326 179 2329
rect 145 2261 179 2285
rect 145 2251 179 2261
rect 145 2193 179 2210
rect 145 2176 179 2193
rect 145 2125 179 2135
rect 145 2101 179 2125
rect 145 2057 179 2060
rect 145 2026 179 2057
rect 145 1955 179 1985
rect 145 1951 179 1955
rect 145 1887 179 1910
rect 145 1876 179 1887
rect 145 1819 179 1835
rect 145 1801 179 1819
rect 145 1751 179 1759
rect 145 1725 179 1751
rect 145 1649 179 1683
rect 468 2455 502 2489
rect 251 2397 285 2415
rect 251 2381 285 2397
rect 251 2329 285 2341
rect 251 2307 285 2329
rect 251 2261 285 2267
rect 251 2233 285 2261
rect 251 2159 285 2193
rect 251 2091 285 2119
rect 251 2085 285 2091
rect 251 2023 285 2045
rect 251 2011 285 2023
rect 251 1955 285 1971
rect 251 1937 285 1955
rect 251 1887 285 1898
rect 251 1864 285 1887
rect 251 1819 285 1825
rect 251 1791 285 1819
rect 251 1751 285 1752
rect 251 1718 285 1751
rect 251 1649 285 1679
rect 251 1645 285 1649
rect 362 2431 396 2435
rect 362 2401 396 2431
rect 362 2329 396 2360
rect 362 2326 396 2329
rect 362 2261 396 2285
rect 362 2251 396 2261
rect 362 2193 396 2210
rect 362 2176 396 2193
rect 362 2125 396 2135
rect 362 2101 396 2125
rect 362 2057 396 2060
rect 362 2026 396 2057
rect 362 1955 396 1985
rect 362 1951 396 1955
rect 362 1887 396 1910
rect 362 1876 396 1887
rect 362 1819 396 1835
rect 362 1801 396 1819
rect 362 1751 396 1760
rect 362 1726 396 1751
rect 362 1683 396 1685
rect 362 1651 396 1683
rect 468 2397 502 2415
rect 468 2381 502 2397
rect 468 2329 502 2341
rect 468 2307 502 2329
rect 468 2261 502 2267
rect 468 2233 502 2261
rect 468 2159 502 2193
rect 468 2091 502 2119
rect 468 2085 502 2091
rect 468 2023 502 2045
rect 468 2011 502 2023
rect 468 1955 502 1971
rect 468 1937 502 1955
rect 468 1887 502 1898
rect 468 1864 502 1887
rect 468 1819 502 1825
rect 468 1791 502 1819
rect 468 1751 502 1752
rect 468 1718 502 1751
rect 468 1649 502 1679
rect 468 1645 502 1649
rect 574 2431 608 2435
rect 574 2401 608 2431
rect 574 2329 608 2360
rect 574 2326 608 2329
rect 574 2261 608 2285
rect 574 2251 608 2261
rect 574 2193 608 2210
rect 574 2176 608 2193
rect 574 2125 608 2135
rect 574 2101 608 2125
rect 574 2057 608 2060
rect 574 2026 608 2057
rect 574 1955 608 1984
rect 574 1950 608 1955
rect 574 1887 608 1908
rect 574 1874 608 1887
rect 574 1819 608 1832
rect 574 1798 608 1819
rect 574 1751 608 1756
rect 574 1722 608 1751
rect 574 1649 608 1680
rect 574 1646 608 1649
rect 834 2170 868 2174
rect 834 2140 868 2170
rect 834 2068 868 2094
rect 834 2060 868 2068
rect 834 2000 868 2014
rect 834 1980 868 2000
rect 834 1932 868 1934
rect 834 1900 868 1932
rect 834 1830 868 1853
rect 834 1819 868 1830
rect 834 1762 868 1772
rect 834 1738 868 1762
rect 834 1660 868 1691
rect 834 1657 868 1660
rect 940 2170 974 2174
rect 940 2140 974 2170
rect 940 2068 974 2094
rect 940 2060 974 2068
rect 940 2000 974 2014
rect 940 1980 974 2000
rect 940 1932 974 1934
rect 940 1900 974 1932
rect 940 1830 974 1853
rect 940 1819 974 1830
rect 940 1762 974 1772
rect 940 1738 974 1762
rect 940 1660 974 1691
rect 940 1657 974 1660
rect 1046 2170 1080 2174
rect 1046 2140 1080 2170
rect 1046 2068 1080 2094
rect 1046 2060 1080 2068
rect 1046 2000 1080 2014
rect 1046 1980 1080 2000
rect 1046 1932 1080 1934
rect 1046 1900 1080 1932
rect 1046 1830 1080 1853
rect 1046 1819 1080 1830
rect 1046 1762 1080 1772
rect 1046 1738 1080 1762
rect 1046 1660 1080 1691
rect 1046 1657 1080 1660
rect 1156 2170 1190 2174
rect 1156 2140 1190 2170
rect 1156 2068 1190 2094
rect 1156 2060 1190 2068
rect 1156 2000 1190 2014
rect 1156 1980 1190 2000
rect 1156 1932 1190 1934
rect 1156 1900 1190 1932
rect 1156 1830 1190 1853
rect 1156 1819 1190 1830
rect 1156 1762 1190 1772
rect 1156 1738 1190 1762
rect 1156 1660 1190 1691
rect 1156 1657 1190 1660
rect 1262 2170 1296 2174
rect 1262 2140 1296 2170
rect 1262 2068 1296 2094
rect 1262 2060 1296 2068
rect 1262 2000 1296 2014
rect 1262 1980 1296 2000
rect 1262 1932 1296 1934
rect 1262 1900 1296 1932
rect 1262 1830 1296 1853
rect 1262 1819 1296 1830
rect 1262 1762 1296 1772
rect 1262 1738 1296 1762
rect 1262 1660 1296 1691
rect 1262 1657 1296 1660
rect 1368 2170 1402 2174
rect 1368 2140 1402 2170
rect 1368 2068 1402 2094
rect 1368 2060 1402 2068
rect 1368 2000 1402 2014
rect 1368 1980 1402 2000
rect 1368 1932 1402 1934
rect 1368 1900 1402 1932
rect 1368 1830 1402 1853
rect 1368 1819 1402 1830
rect 1368 1762 1402 1772
rect 1368 1738 1402 1762
rect 1368 1660 1402 1691
rect 1368 1657 1402 1660
rect 879 1500 913 1510
rect 879 1476 913 1500
rect 97 1419 100 1453
rect 100 1419 131 1453
rect 194 1419 224 1453
rect 224 1419 228 1453
rect 414 1444 448 1457
rect 414 1423 448 1444
rect 414 1354 448 1385
rect 414 1351 448 1354
rect 529 1444 563 1457
rect 529 1423 563 1444
rect 879 1410 913 1438
rect 879 1404 913 1410
rect 1001 1534 1035 1538
rect 1001 1504 1035 1534
rect 1213 1500 1217 1534
rect 1217 1500 1247 1534
rect 1297 1500 1307 1534
rect 1307 1500 1331 1534
rect 1001 1444 1035 1466
rect 1001 1432 1035 1444
rect 529 1354 563 1385
rect 529 1351 563 1354
rect 1238 1387 1272 1421
rect 1370 1387 1404 1421
rect 1238 1305 1272 1339
rect 1370 1305 1404 1339
rect 949 1273 983 1274
rect 949 1240 980 1273
rect 980 1240 983 1273
rect 87 1171 91 1205
rect 91 1171 121 1205
rect 166 1171 196 1205
rect 196 1171 200 1205
rect 280 1171 284 1205
rect 284 1171 314 1205
rect 379 1171 413 1205
rect 478 1171 508 1205
rect 508 1171 512 1205
rect 949 1171 980 1202
rect 980 1171 983 1202
rect 949 1168 983 1171
rect 1102 1273 1136 1274
rect 1102 1240 1136 1273
rect 1102 1171 1136 1202
rect 1102 1168 1136 1171
rect 1238 1223 1272 1257
rect 1370 1223 1404 1257
rect 1238 1141 1272 1175
rect 1370 1141 1404 1175
rect 1305 1082 1339 1092
rect 67 985 101 1019
rect 67 917 101 941
rect 67 907 101 917
rect 67 849 101 863
rect 67 829 101 849
rect 67 781 101 785
rect 67 751 101 781
rect 67 679 101 707
rect 67 673 101 679
rect 67 611 101 629
rect 67 595 101 611
rect 67 543 101 551
rect 67 517 101 543
rect 67 441 101 473
rect 67 439 101 441
rect 67 373 101 396
rect 67 362 101 373
rect 67 305 101 319
rect 67 285 101 305
rect 67 237 101 242
rect 67 208 101 237
rect 67 135 101 165
rect 67 131 101 135
rect 223 985 257 1019
rect 223 917 257 941
rect 223 907 257 917
rect 223 849 257 863
rect 223 829 257 849
rect 223 781 257 785
rect 223 751 257 781
rect 223 679 257 707
rect 223 673 257 679
rect 223 611 257 629
rect 223 595 257 611
rect 223 543 257 551
rect 223 517 257 543
rect 223 441 257 473
rect 223 439 257 441
rect 223 373 257 396
rect 223 362 257 373
rect 223 305 257 319
rect 223 285 257 305
rect 223 237 257 242
rect 223 208 257 237
rect 223 135 257 165
rect 223 131 257 135
rect 379 985 413 1019
rect 379 917 413 941
rect 379 907 413 917
rect 379 849 413 863
rect 379 829 413 849
rect 379 781 413 785
rect 379 751 413 781
rect 379 679 413 707
rect 379 673 413 679
rect 379 611 413 629
rect 379 595 413 611
rect 379 543 413 551
rect 379 517 413 543
rect 379 441 413 473
rect 379 439 413 441
rect 379 373 413 396
rect 379 362 413 373
rect 379 305 413 319
rect 379 285 413 305
rect 379 237 413 242
rect 379 208 413 237
rect 379 135 413 165
rect 379 131 413 135
rect 535 985 569 1019
rect 535 917 569 941
rect 535 907 569 917
rect 535 849 569 863
rect 535 829 569 849
rect 535 781 569 785
rect 535 751 569 781
rect 535 679 569 707
rect 535 673 569 679
rect 535 611 569 629
rect 535 595 569 611
rect 535 543 569 551
rect 535 517 569 543
rect 535 441 569 473
rect 535 439 569 441
rect 535 373 569 396
rect 535 362 569 373
rect 535 305 569 319
rect 535 285 569 305
rect 535 237 569 242
rect 535 208 569 237
rect 535 135 569 165
rect 535 131 569 135
rect 869 985 903 1019
rect 869 917 903 941
rect 869 907 903 917
rect 869 849 903 863
rect 869 829 903 849
rect 869 781 903 785
rect 869 751 903 781
rect 869 679 903 707
rect 869 673 903 679
rect 869 611 903 629
rect 869 595 903 611
rect 869 543 903 551
rect 869 517 903 543
rect 869 441 903 473
rect 869 439 903 441
rect 869 373 903 396
rect 869 362 903 373
rect 869 305 903 319
rect 869 285 903 305
rect 869 237 903 242
rect 869 208 903 237
rect 869 135 903 165
rect 869 131 903 135
rect 1025 985 1059 1019
rect 1025 917 1059 941
rect 1025 907 1059 917
rect 1025 849 1059 863
rect 1025 829 1059 849
rect 1025 781 1059 785
rect 1025 751 1059 781
rect 1025 679 1059 707
rect 1025 673 1059 679
rect 1025 611 1059 629
rect 1025 595 1059 611
rect 1025 543 1059 551
rect 1025 517 1059 543
rect 1025 441 1059 473
rect 1025 439 1059 441
rect 1025 373 1059 396
rect 1025 362 1059 373
rect 1025 305 1059 319
rect 1025 285 1059 305
rect 1025 237 1059 242
rect 1025 208 1059 237
rect 1025 135 1059 165
rect 1025 131 1059 135
rect 1305 1058 1339 1082
rect 1181 985 1215 1019
rect 1305 981 1339 1015
rect 1181 917 1215 941
rect 1181 907 1215 917
rect 1305 937 1339 938
rect 1305 904 1339 937
rect 1181 849 1215 863
rect 1181 829 1215 849
rect 1305 859 1339 861
rect 1305 827 1339 859
rect 1181 781 1215 785
rect 1181 751 1215 781
rect 1305 750 1339 784
rect 1181 679 1215 707
rect 1181 673 1215 679
rect 1305 673 1339 707
rect 1181 611 1215 629
rect 1181 595 1215 611
rect 1305 601 1339 630
rect 1305 596 1339 601
rect 1181 543 1215 551
rect 1181 517 1215 543
rect 1305 523 1339 553
rect 1305 519 1339 523
rect 1181 441 1215 473
rect 1305 442 1339 476
rect 1181 439 1215 441
rect 1181 373 1215 396
rect 1181 362 1215 373
rect 1305 377 1339 399
rect 1305 365 1339 377
rect 1181 305 1215 319
rect 1181 285 1215 305
rect 1305 299 1339 321
rect 1305 287 1339 299
rect 1181 237 1215 242
rect 1181 208 1215 237
rect 1305 209 1339 243
rect 1181 135 1215 165
rect 1181 131 1215 135
rect 1305 153 1339 165
rect 1305 131 1339 153
rect 57 15 83 49
rect 83 15 91 49
rect 141 15 171 49
rect 171 15 175 49
rect 224 15 258 49
rect 307 15 341 49
rect 390 15 424 49
rect 473 15 507 49
rect 556 15 590 49
<< metal1 >>
rect 55 2609 774 2615
rect 55 2575 67 2609
rect 101 2575 149 2609
rect 183 2575 231 2609
rect 265 2575 313 2609
rect 347 2575 395 2609
rect 429 2575 476 2609
rect 510 2575 557 2609
rect 591 2575 774 2609
tri 33 2517 55 2539 se
rect 55 2517 774 2575
rect 33 2489 89 2517
tri 89 2489 117 2517 nw
tri 209 2501 225 2517 ne
rect 225 2501 301 2517
tri 225 2489 237 2501 ne
rect 237 2489 301 2501
tri 301 2489 329 2517 nw
tri 424 2489 452 2517 ne
rect 452 2501 528 2517
tri 528 2501 544 2517 nw
tri 618 2501 634 2517 ne
rect 634 2501 774 2517
rect 452 2489 508 2501
rect 33 2455 39 2489
rect 73 2455 79 2489
tri 79 2479 89 2489 nw
tri 237 2481 245 2489 ne
rect 33 2415 79 2455
rect 245 2455 251 2489
rect 285 2455 291 2489
tri 291 2479 301 2489 nw
tri 452 2479 462 2489 ne
rect 33 2381 39 2415
rect 73 2381 79 2415
rect 33 2341 79 2381
rect 33 2307 39 2341
rect 73 2307 79 2341
rect 33 2267 79 2307
rect 33 2233 39 2267
rect 73 2233 79 2267
rect 33 2193 79 2233
rect 33 2159 39 2193
rect 73 2159 79 2193
rect 33 2119 79 2159
rect 33 2085 39 2119
rect 73 2085 79 2119
rect 33 2045 79 2085
rect 33 2011 39 2045
rect 73 2011 79 2045
rect 33 1971 79 2011
rect 33 1937 39 1971
rect 73 1937 79 1971
rect 33 1898 79 1937
rect 33 1864 39 1898
rect 73 1864 79 1898
rect 33 1825 79 1864
rect 33 1791 39 1825
rect 73 1791 79 1825
rect 33 1752 79 1791
rect 33 1718 39 1752
rect 73 1718 79 1752
rect 33 1679 79 1718
rect 33 1645 39 1679
rect 73 1645 79 1679
rect 33 1633 79 1645
rect 136 2435 188 2447
rect 136 2401 145 2435
rect 179 2401 188 2435
rect 136 2360 188 2401
rect 136 2326 145 2360
rect 179 2326 188 2360
rect 136 2285 188 2326
rect 136 2251 145 2285
rect 179 2251 188 2285
rect 136 2210 188 2251
rect 136 2176 145 2210
rect 179 2176 188 2210
rect 136 2135 188 2176
rect 136 2101 145 2135
rect 179 2101 188 2135
rect 136 2092 188 2101
rect 136 2028 145 2040
rect 179 2028 188 2040
rect 136 1951 145 1976
rect 179 1951 188 1976
rect 136 1910 188 1951
rect 136 1876 145 1910
rect 179 1876 188 1910
rect 136 1835 188 1876
rect 136 1801 145 1835
rect 179 1801 188 1835
rect 136 1759 188 1801
rect 136 1725 145 1759
rect 179 1725 188 1759
rect 136 1683 188 1725
rect 136 1649 145 1683
rect 179 1649 188 1683
rect 136 1637 188 1649
rect 245 2415 291 2455
rect 462 2455 468 2489
rect 502 2455 508 2489
tri 508 2481 528 2501 nw
tri 634 2481 654 2501 ne
rect 654 2481 774 2501
tri 654 2479 656 2481 ne
rect 656 2479 774 2481
tri 656 2477 658 2479 ne
rect 245 2381 251 2415
rect 285 2381 291 2415
rect 245 2341 291 2381
rect 245 2307 251 2341
rect 285 2307 291 2341
rect 245 2267 291 2307
rect 245 2233 251 2267
rect 285 2233 291 2267
rect 245 2193 291 2233
rect 245 2159 251 2193
rect 285 2159 291 2193
rect 245 2119 291 2159
rect 245 2085 251 2119
rect 285 2085 291 2119
rect 245 2045 291 2085
rect 245 2011 251 2045
rect 285 2011 291 2045
rect 245 1971 291 2011
rect 245 1937 251 1971
rect 285 1937 291 1971
rect 245 1898 291 1937
rect 245 1864 251 1898
rect 285 1864 291 1898
rect 245 1825 291 1864
rect 245 1791 251 1825
rect 285 1791 291 1825
rect 245 1752 291 1791
rect 245 1718 251 1752
rect 285 1718 291 1752
rect 245 1679 291 1718
rect 245 1645 251 1679
rect 285 1645 291 1679
rect 245 1633 291 1645
rect 353 2435 405 2447
rect 353 2401 362 2435
rect 396 2401 405 2435
rect 353 2360 405 2401
rect 353 2326 362 2360
rect 396 2326 405 2360
rect 353 2285 405 2326
rect 353 2251 362 2285
rect 396 2251 405 2285
rect 353 2210 405 2251
rect 353 2176 362 2210
rect 396 2176 405 2210
rect 353 2135 405 2176
rect 353 2101 362 2135
rect 396 2101 405 2135
rect 353 2060 405 2101
rect 353 2026 362 2060
rect 396 2026 405 2060
rect 353 1985 405 2026
rect 353 1951 362 1985
rect 396 1951 405 1985
rect 353 1934 405 1951
rect 353 1876 362 1882
rect 396 1876 405 1882
rect 353 1870 405 1876
rect 353 1801 362 1818
rect 396 1801 405 1818
rect 353 1760 405 1801
rect 353 1726 362 1760
rect 396 1726 405 1760
rect 353 1685 405 1726
rect 353 1651 362 1685
rect 396 1651 405 1685
rect 353 1497 405 1651
rect 462 2415 508 2455
rect 462 2381 468 2415
rect 502 2381 508 2415
rect 462 2341 508 2381
rect 462 2307 468 2341
rect 502 2307 508 2341
rect 462 2267 508 2307
rect 462 2233 468 2267
rect 502 2233 508 2267
rect 462 2193 508 2233
rect 462 2159 468 2193
rect 502 2159 508 2193
rect 462 2119 508 2159
rect 462 2085 468 2119
rect 502 2085 508 2119
rect 462 2045 508 2085
rect 462 2011 468 2045
rect 502 2011 508 2045
rect 462 1971 508 2011
rect 462 1937 468 1971
rect 502 1937 508 1971
rect 462 1898 508 1937
rect 462 1864 468 1898
rect 502 1864 508 1898
rect 462 1825 508 1864
rect 462 1791 468 1825
rect 502 1791 508 1825
rect 462 1752 508 1791
rect 462 1718 468 1752
rect 502 1718 508 1752
rect 462 1679 508 1718
rect 462 1645 468 1679
rect 502 1645 508 1679
rect 462 1633 508 1645
rect 565 2435 617 2447
rect 565 2401 574 2435
rect 608 2401 617 2435
rect 565 2360 617 2401
rect 565 2326 574 2360
rect 608 2326 617 2360
rect 565 2285 617 2326
rect 565 2251 574 2285
rect 608 2251 617 2285
rect 565 2210 617 2251
rect 565 2176 574 2210
rect 608 2176 617 2210
rect 565 2135 617 2176
rect 565 2101 574 2135
rect 608 2101 617 2135
rect 565 2060 617 2101
rect 565 2026 574 2060
rect 608 2026 617 2060
rect 565 1984 617 2026
rect 565 1950 574 1984
rect 608 1950 617 1984
rect 565 1908 617 1950
rect 565 1874 574 1908
rect 608 1874 617 1908
rect 565 1832 617 1874
rect 565 1798 574 1832
rect 608 1798 617 1832
rect 565 1766 617 1798
rect 565 1702 617 1714
rect 565 1646 574 1650
rect 608 1646 617 1650
rect 565 1634 617 1646
rect 405 1463 457 1469
rect 85 1410 91 1462
rect 143 1410 183 1462
rect 235 1410 241 1462
rect 405 1399 457 1411
rect 405 1339 457 1347
rect 520 1457 572 1469
rect 520 1435 529 1457
rect 563 1435 572 1457
rect 520 1371 529 1383
rect 563 1371 572 1383
rect 520 1313 572 1319
rect 75 1162 81 1214
rect 133 1162 154 1214
rect 206 1162 212 1214
rect 268 1162 274 1214
rect 326 1162 338 1214
rect 390 1205 402 1214
rect 390 1162 402 1171
rect 454 1162 466 1214
rect 518 1162 524 1214
rect 58 1019 110 1031
rect 58 985 67 1019
rect 101 985 110 1019
rect 58 941 110 985
rect 58 907 67 941
rect 101 907 110 941
rect 58 863 110 907
rect 214 1026 266 1032
rect 214 941 266 974
rect 214 938 223 941
rect 257 938 266 941
tri 110 863 112 865 sw
rect 214 863 266 886
rect 58 829 67 863
rect 101 831 112 863
tri 112 831 144 863 sw
rect 101 829 173 831
rect 58 825 173 829
rect 58 785 121 825
rect 58 751 67 785
rect 101 773 121 785
rect 101 751 173 773
rect 58 737 173 751
rect 58 707 121 737
rect 58 673 67 707
rect 101 685 121 707
rect 101 679 173 685
rect 214 829 223 863
rect 257 829 266 863
rect 214 785 266 829
rect 214 751 223 785
rect 257 751 266 785
rect 214 707 266 751
rect 101 673 131 679
tri 131 673 137 679 nw
rect 214 673 223 707
rect 257 673 266 707
rect 58 629 110 673
tri 110 652 131 673 nw
rect 58 595 67 629
rect 101 595 110 629
rect 58 551 110 595
rect 58 517 67 551
rect 101 517 110 551
rect 58 473 110 517
rect 58 439 67 473
rect 101 439 110 473
rect 58 396 110 439
rect 58 362 67 396
rect 101 362 110 396
rect 58 319 110 362
rect 58 285 67 319
rect 101 285 110 319
rect 58 242 110 285
rect 58 208 67 242
rect 101 208 110 242
rect 58 165 110 208
rect 58 131 67 165
rect 101 131 110 165
rect 58 119 110 131
rect 214 629 266 673
rect 214 595 223 629
rect 257 595 266 629
rect 214 551 266 595
rect 214 517 223 551
rect 257 517 266 551
rect 214 473 266 517
rect 214 439 223 473
rect 257 439 266 473
rect 214 396 266 439
rect 214 362 223 396
rect 257 362 266 396
rect 214 319 266 362
rect 214 285 223 319
rect 257 285 266 319
rect 214 242 266 285
rect 214 208 223 242
rect 257 208 266 242
rect 214 165 266 208
rect 214 131 223 165
rect 257 131 266 165
rect 214 119 266 131
rect 370 1019 422 1031
rect 370 985 379 1019
rect 413 985 422 1019
rect 370 941 422 985
rect 370 907 379 941
rect 413 907 422 941
rect 370 863 422 907
rect 370 829 379 863
rect 413 829 422 863
rect 370 825 422 829
rect 370 751 379 773
rect 413 751 422 773
rect 370 737 422 751
rect 370 673 379 685
rect 413 673 422 685
rect 370 629 422 673
rect 370 595 379 629
rect 413 595 422 629
rect 370 551 422 595
rect 370 517 379 551
rect 413 517 422 551
rect 370 473 422 517
rect 370 439 379 473
rect 413 439 422 473
rect 370 396 422 439
rect 370 362 379 396
rect 413 362 422 396
rect 370 319 422 362
rect 370 285 379 319
rect 413 285 422 319
rect 370 242 422 285
rect 370 208 379 242
rect 413 208 422 242
rect 370 165 422 208
rect 370 131 379 165
rect 413 131 422 165
rect 370 119 422 131
rect 526 1026 578 1032
rect 526 941 578 974
rect 526 938 535 941
rect 569 938 578 941
rect 526 863 578 886
rect 526 829 535 863
rect 569 829 578 863
rect 526 785 578 829
rect 526 751 535 785
rect 569 751 578 785
rect 526 707 578 751
rect 526 673 535 707
rect 569 673 578 707
rect 526 629 578 673
rect 526 595 535 629
rect 569 595 578 629
rect 526 551 578 595
rect 526 517 535 551
rect 569 517 578 551
rect 526 473 578 517
rect 526 439 535 473
rect 569 439 578 473
rect 526 396 578 439
rect 526 362 535 396
rect 569 362 578 396
rect 526 319 578 362
rect 526 285 535 319
rect 569 285 578 319
rect 526 242 578 285
rect 526 208 535 242
rect 569 208 578 242
rect 526 165 578 208
rect 526 131 535 165
rect 569 131 578 165
rect 526 119 578 131
rect 658 825 774 2479
rect 934 2240 1518 2330
rect 934 2223 1218 2240
tri 1218 2223 1235 2240 nw
tri 1314 2223 1331 2240 ne
rect 1331 2223 1518 2240
rect 825 2174 877 2186
rect 825 2140 834 2174
rect 868 2140 877 2174
rect 825 2094 877 2140
rect 825 2060 834 2094
rect 868 2060 877 2094
rect 825 2014 877 2060
rect 825 1980 834 2014
rect 868 1980 877 2014
rect 825 1934 877 1980
rect 825 1900 834 1934
rect 868 1900 877 1934
rect 825 1853 877 1900
rect 825 1819 834 1853
rect 868 1819 877 1853
rect 825 1772 877 1819
rect 825 1766 834 1772
rect 868 1766 877 1772
rect 825 1702 877 1714
rect 825 1644 877 1650
rect 934 2174 980 2223
tri 980 2187 1016 2223 nw
tri 1122 2195 1150 2223 ne
rect 934 2140 940 2174
rect 974 2140 980 2174
rect 934 2094 980 2140
rect 934 2060 940 2094
rect 974 2060 980 2094
rect 934 2014 980 2060
rect 934 1980 940 2014
rect 974 1980 980 2014
rect 934 1934 980 1980
rect 934 1900 940 1934
rect 974 1900 980 1934
rect 934 1853 980 1900
rect 934 1819 940 1853
rect 974 1819 980 1853
rect 934 1772 980 1819
rect 934 1738 940 1772
rect 974 1738 980 1772
rect 934 1691 980 1738
rect 934 1657 940 1691
rect 974 1657 980 1691
rect 934 1645 980 1657
rect 1037 2174 1089 2186
rect 1037 2140 1046 2174
rect 1080 2140 1089 2174
rect 1037 2094 1089 2140
rect 1037 2060 1046 2094
rect 1080 2060 1089 2094
rect 1037 2014 1089 2060
rect 1037 1980 1046 2014
rect 1080 1980 1089 2014
rect 1037 1934 1089 1980
rect 1037 1870 1089 1882
rect 1037 1772 1089 1818
rect 1037 1738 1046 1772
rect 1080 1738 1089 1772
rect 1037 1691 1089 1738
rect 1037 1657 1046 1691
rect 1080 1657 1089 1691
rect 1037 1634 1089 1657
rect 1150 2174 1196 2223
tri 1196 2201 1218 2223 nw
tri 1331 2201 1353 2223 ne
rect 1353 2201 1518 2223
tri 1353 2195 1359 2201 ne
rect 1359 2195 1518 2201
tri 1359 2192 1362 2195 ne
rect 1150 2140 1156 2174
rect 1190 2140 1196 2174
rect 1150 2094 1196 2140
rect 1150 2060 1156 2094
rect 1190 2060 1196 2094
rect 1150 2014 1196 2060
rect 1150 1980 1156 2014
rect 1190 1980 1196 2014
rect 1150 1934 1196 1980
rect 1150 1900 1156 1934
rect 1190 1900 1196 1934
rect 1150 1853 1196 1900
rect 1150 1819 1156 1853
rect 1190 1819 1196 1853
rect 1150 1772 1196 1819
rect 1150 1738 1156 1772
rect 1190 1738 1196 1772
rect 1150 1691 1196 1738
rect 1150 1657 1156 1691
rect 1190 1657 1196 1691
rect 1150 1645 1196 1657
rect 1253 2174 1305 2186
rect 1253 2140 1262 2174
rect 1296 2140 1305 2174
rect 1253 2094 1305 2140
rect 1253 2092 1262 2094
rect 1296 2092 1305 2094
rect 1253 2028 1305 2040
rect 1253 1934 1305 1976
rect 1253 1900 1262 1934
rect 1296 1900 1305 1934
rect 1253 1853 1305 1900
rect 1253 1819 1262 1853
rect 1296 1819 1305 1853
rect 1253 1772 1305 1819
rect 1253 1738 1262 1772
rect 1296 1738 1305 1772
rect 1253 1691 1305 1738
rect 1253 1657 1262 1691
rect 1296 1657 1305 1691
rect 1253 1645 1305 1657
rect 1362 2174 1518 2195
rect 1362 2140 1368 2174
rect 1402 2140 1518 2174
rect 1362 2094 1518 2140
rect 1362 2060 1368 2094
rect 1402 2060 1518 2094
rect 1362 2014 1518 2060
rect 1362 1980 1368 2014
rect 1402 1980 1518 2014
rect 1362 1934 1518 1980
rect 1362 1900 1368 1934
rect 1402 1900 1518 1934
rect 1362 1853 1518 1900
rect 1362 1819 1368 1853
rect 1402 1819 1518 1853
rect 1362 1772 1518 1819
rect 1362 1738 1368 1772
rect 1402 1738 1518 1772
rect 1362 1691 1518 1738
rect 1362 1657 1368 1691
rect 1402 1657 1518 1691
rect 1362 1645 1518 1657
tri 1388 1634 1399 1645 ne
rect 1399 1634 1518 1645
tri 1399 1609 1424 1634 ne
rect 992 1544 1044 1550
rect 710 773 722 825
rect 658 737 774 773
rect 710 685 722 737
tri 618 55 658 95 se
rect 658 55 774 685
rect 814 1516 922 1522
rect 814 1464 870 1516
rect 814 1452 922 1464
rect 814 1400 870 1452
rect 992 1480 1044 1492
rect 1201 1491 1207 1543
rect 1259 1534 1299 1543
rect 1259 1500 1297 1534
rect 1259 1491 1299 1500
rect 1351 1491 1357 1543
tri 1399 1433 1424 1458 se
rect 1424 1433 1518 1634
rect 992 1420 1044 1428
rect 1232 1421 1518 1433
rect 814 1394 922 1400
rect 814 1392 920 1394
tri 920 1392 922 1394 nw
rect 814 1387 915 1392
tri 915 1387 920 1392 nw
rect 1232 1387 1238 1421
rect 1272 1387 1370 1421
rect 1404 1387 1518 1421
rect 814 1058 868 1387
tri 868 1340 915 1387 nw
rect 1232 1339 1518 1387
rect 1232 1305 1238 1339
rect 1272 1305 1370 1339
rect 1404 1305 1518 1339
rect 940 1280 992 1286
rect 940 1214 992 1228
rect 940 1156 992 1162
rect 1090 1280 1142 1286
rect 1090 1214 1142 1228
rect 1090 1156 1142 1162
rect 1232 1257 1518 1305
rect 1232 1223 1238 1257
rect 1272 1223 1370 1257
rect 1404 1223 1518 1257
rect 1232 1175 1518 1223
rect 1232 1141 1238 1175
rect 1272 1141 1370 1175
rect 1404 1141 1518 1175
rect 1232 1092 1518 1141
tri 1205 1061 1232 1088 se
rect 1232 1061 1305 1092
tri 868 1058 871 1061 sw
tri 1202 1058 1205 1061 se
rect 1205 1058 1305 1061
rect 1339 1058 1518 1092
rect 814 1032 871 1058
tri 871 1032 897 1058 sw
tri 1176 1032 1202 1058 se
rect 1202 1032 1518 1058
rect 814 1026 930 1032
tri 1175 1031 1176 1032 se
rect 1176 1031 1518 1032
rect 866 1019 878 1026
rect 866 985 869 1019
rect 866 974 878 985
rect 814 941 930 974
rect 814 938 869 941
rect 903 938 930 941
rect 866 907 869 938
rect 866 886 878 907
rect 814 880 930 886
rect 814 863 913 880
tri 913 863 930 880 nw
rect 1019 1019 1065 1031
rect 1019 985 1025 1019
rect 1059 985 1065 1019
rect 1019 941 1065 985
rect 1019 907 1025 941
rect 1059 907 1065 941
rect 1019 863 1065 907
rect 814 829 869 863
rect 903 829 912 863
tri 912 862 913 863 nw
rect 814 785 912 829
rect 814 751 869 785
rect 903 751 912 785
rect 814 707 912 751
rect 814 673 869 707
rect 903 673 912 707
rect 814 629 912 673
rect 814 595 869 629
rect 903 595 912 629
rect 814 551 912 595
rect 814 517 869 551
rect 903 517 912 551
rect 814 473 912 517
rect 814 439 869 473
rect 903 439 912 473
rect 814 396 912 439
rect 814 362 869 396
rect 903 362 912 396
rect 814 319 912 362
rect 814 285 869 319
rect 903 285 912 319
rect 814 242 912 285
rect 814 208 869 242
rect 903 208 912 242
rect 814 165 912 208
rect 814 131 869 165
rect 903 131 912 165
rect 814 119 912 131
rect 1019 829 1025 863
rect 1059 829 1065 863
rect 1019 785 1065 829
rect 1019 751 1025 785
rect 1059 751 1065 785
rect 1019 707 1065 751
rect 1019 673 1025 707
rect 1059 673 1065 707
rect 1019 629 1065 673
rect 1019 595 1025 629
rect 1059 595 1065 629
rect 1019 551 1065 595
rect 1019 517 1025 551
rect 1059 517 1065 551
rect 1019 473 1065 517
rect 1019 439 1025 473
rect 1059 439 1065 473
rect 1019 396 1065 439
rect 1019 362 1025 396
rect 1059 362 1065 396
rect 1019 319 1065 362
rect 1019 285 1025 319
rect 1059 285 1065 319
rect 1019 242 1065 285
rect 1019 208 1025 242
rect 1059 208 1065 242
rect 1019 165 1065 208
rect 1019 131 1025 165
rect 1059 131 1065 165
rect 1019 119 1065 131
rect 1175 1019 1518 1031
rect 1175 985 1181 1019
rect 1215 1015 1518 1019
rect 1215 985 1305 1015
rect 1175 981 1305 985
rect 1339 981 1518 1015
rect 1175 941 1518 981
rect 1175 907 1181 941
rect 1215 938 1518 941
rect 1215 907 1305 938
rect 1175 904 1305 907
rect 1339 904 1518 938
rect 1175 863 1518 904
rect 1175 829 1181 863
rect 1215 861 1518 863
rect 1215 829 1305 861
rect 1175 827 1305 829
rect 1339 827 1518 861
rect 1175 785 1518 827
rect 1175 751 1181 785
rect 1215 784 1518 785
rect 1215 751 1305 784
rect 1175 750 1305 751
rect 1339 750 1518 784
rect 1175 707 1518 750
rect 1175 673 1181 707
rect 1215 673 1305 707
rect 1339 673 1518 707
rect 1175 630 1518 673
rect 1175 629 1305 630
rect 1175 595 1181 629
rect 1215 596 1305 629
rect 1339 596 1518 630
rect 1215 595 1518 596
rect 1175 553 1518 595
rect 1175 551 1305 553
rect 1175 517 1181 551
rect 1215 519 1305 551
rect 1339 519 1518 553
rect 1215 517 1518 519
rect 1175 476 1518 517
rect 1175 473 1305 476
rect 1175 439 1181 473
rect 1215 442 1305 473
rect 1339 442 1518 476
rect 1215 439 1518 442
rect 1175 399 1518 439
rect 1175 396 1305 399
rect 1175 362 1181 396
rect 1215 365 1305 396
rect 1339 365 1518 399
rect 1215 362 1518 365
rect 1175 321 1518 362
rect 1175 319 1305 321
rect 1175 285 1181 319
rect 1215 287 1305 319
rect 1339 287 1518 321
rect 1215 285 1518 287
rect 1175 243 1518 285
rect 1175 242 1305 243
rect 1175 208 1181 242
rect 1215 209 1305 242
rect 1339 209 1518 243
rect 1215 208 1518 209
rect 1175 165 1518 208
rect 1175 131 1181 165
rect 1215 131 1305 165
rect 1339 131 1518 165
rect 1175 119 1518 131
rect 1175 105 1504 119
tri 1504 105 1518 119 nw
rect 45 49 774 55
rect 45 15 57 49
rect 91 15 141 49
rect 175 15 224 49
rect 258 15 307 49
rect 341 15 390 49
rect 424 15 473 49
rect 507 15 556 49
rect 590 15 774 49
rect 45 9 774 15
tri 1079 9 1175 105 se
rect 1175 9 1467 105
tri 1467 68 1504 105 nw
tri 1043 -27 1079 9 se
rect 1079 -27 1467 9
rect 448 -228 1467 -27
tri 1467 -228 1476 -219 sw
<< via1 >>
rect 136 2060 188 2092
rect 136 2040 145 2060
rect 145 2040 179 2060
rect 179 2040 188 2060
rect 136 2026 145 2028
rect 145 2026 179 2028
rect 179 2026 188 2028
rect 136 1985 188 2026
rect 136 1976 145 1985
rect 145 1976 179 1985
rect 179 1976 188 1985
rect 353 1910 405 1934
rect 353 1882 362 1910
rect 362 1882 396 1910
rect 396 1882 405 1910
rect 353 1835 405 1870
rect 353 1818 362 1835
rect 362 1818 396 1835
rect 396 1818 405 1835
rect 565 1756 617 1766
rect 565 1722 574 1756
rect 574 1722 608 1756
rect 608 1722 617 1756
rect 565 1714 617 1722
rect 565 1680 617 1702
rect 565 1650 574 1680
rect 574 1650 608 1680
rect 608 1650 617 1680
rect 91 1453 143 1462
rect 91 1419 97 1453
rect 97 1419 131 1453
rect 131 1419 143 1453
rect 91 1410 143 1419
rect 183 1453 235 1462
rect 183 1419 194 1453
rect 194 1419 228 1453
rect 228 1419 235 1453
rect 183 1410 235 1419
rect 405 1457 457 1463
rect 405 1423 414 1457
rect 414 1423 448 1457
rect 448 1423 457 1457
rect 405 1411 457 1423
rect 405 1385 457 1399
rect 405 1351 414 1385
rect 414 1351 448 1385
rect 448 1351 457 1385
rect 405 1347 457 1351
rect 520 1423 529 1435
rect 529 1423 563 1435
rect 563 1423 572 1435
rect 520 1385 572 1423
rect 520 1383 529 1385
rect 529 1383 563 1385
rect 563 1383 572 1385
rect 520 1351 529 1371
rect 529 1351 563 1371
rect 563 1351 572 1371
rect 520 1319 572 1351
rect 81 1205 133 1214
rect 81 1171 87 1205
rect 87 1171 121 1205
rect 121 1171 133 1205
rect 81 1162 133 1171
rect 154 1205 206 1214
rect 154 1171 166 1205
rect 166 1171 200 1205
rect 200 1171 206 1205
rect 154 1162 206 1171
rect 274 1205 326 1214
rect 274 1171 280 1205
rect 280 1171 314 1205
rect 314 1171 326 1205
rect 274 1162 326 1171
rect 338 1205 390 1214
rect 402 1205 454 1214
rect 338 1171 379 1205
rect 379 1171 390 1205
rect 402 1171 413 1205
rect 413 1171 454 1205
rect 338 1162 390 1171
rect 402 1162 454 1171
rect 466 1205 518 1214
rect 466 1171 478 1205
rect 478 1171 512 1205
rect 512 1171 518 1205
rect 466 1162 518 1171
rect 214 1019 266 1026
rect 214 985 223 1019
rect 223 985 257 1019
rect 257 985 266 1019
rect 214 974 266 985
rect 214 907 223 938
rect 223 907 257 938
rect 257 907 266 938
rect 214 886 266 907
rect 121 773 173 825
rect 121 685 173 737
rect 370 785 422 825
rect 370 773 379 785
rect 379 773 413 785
rect 413 773 422 785
rect 370 707 422 737
rect 370 685 379 707
rect 379 685 413 707
rect 413 685 422 707
rect 526 1019 578 1026
rect 526 985 535 1019
rect 535 985 569 1019
rect 569 985 578 1019
rect 526 974 578 985
rect 526 907 535 938
rect 535 907 569 938
rect 569 907 578 938
rect 526 886 578 907
rect 825 1738 834 1766
rect 834 1738 868 1766
rect 868 1738 877 1766
rect 825 1714 877 1738
rect 825 1691 877 1702
rect 825 1657 834 1691
rect 834 1657 868 1691
rect 868 1657 877 1691
rect 825 1650 877 1657
rect 1037 1900 1046 1934
rect 1046 1900 1080 1934
rect 1080 1900 1089 1934
rect 1037 1882 1089 1900
rect 1037 1853 1089 1870
rect 1037 1819 1046 1853
rect 1046 1819 1080 1853
rect 1080 1819 1089 1853
rect 1037 1818 1089 1819
rect 1253 2060 1262 2092
rect 1262 2060 1296 2092
rect 1296 2060 1305 2092
rect 1253 2040 1305 2060
rect 1253 2014 1305 2028
rect 1253 1980 1262 2014
rect 1262 1980 1296 2014
rect 1296 1980 1305 2014
rect 1253 1976 1305 1980
rect 992 1538 1044 1544
rect 658 773 710 825
rect 722 773 774 825
rect 658 685 710 737
rect 722 685 774 737
rect 870 1510 922 1516
rect 870 1476 879 1510
rect 879 1476 913 1510
rect 913 1476 922 1510
rect 870 1464 922 1476
rect 870 1438 922 1452
rect 870 1404 879 1438
rect 879 1404 913 1438
rect 913 1404 922 1438
rect 992 1504 1001 1538
rect 1001 1504 1035 1538
rect 1035 1504 1044 1538
rect 992 1492 1044 1504
rect 1207 1534 1259 1543
rect 1299 1534 1351 1543
rect 1207 1500 1213 1534
rect 1213 1500 1247 1534
rect 1247 1500 1259 1534
rect 1299 1500 1331 1534
rect 1331 1500 1351 1534
rect 1207 1491 1259 1500
rect 1299 1491 1351 1500
rect 992 1466 1044 1480
rect 992 1432 1001 1466
rect 1001 1432 1035 1466
rect 1035 1432 1044 1466
rect 992 1428 1044 1432
rect 870 1400 922 1404
rect 940 1274 992 1280
rect 940 1240 949 1274
rect 949 1240 983 1274
rect 983 1240 992 1274
rect 940 1228 992 1240
rect 940 1202 992 1214
rect 940 1168 949 1202
rect 949 1168 983 1202
rect 983 1168 992 1202
rect 940 1162 992 1168
rect 1090 1274 1142 1280
rect 1090 1240 1102 1274
rect 1102 1240 1136 1274
rect 1136 1240 1142 1274
rect 1090 1228 1142 1240
rect 1090 1202 1142 1214
rect 1090 1168 1102 1202
rect 1102 1168 1136 1202
rect 1136 1168 1142 1202
rect 1090 1162 1142 1168
rect 814 974 866 1026
rect 878 1019 930 1026
rect 878 985 903 1019
rect 903 985 930 1019
rect 878 974 930 985
rect 814 886 866 938
rect 878 907 903 938
rect 903 907 930 938
rect 878 886 930 907
<< metal2 >>
rect 136 2092 1305 2098
rect 188 2040 1253 2092
rect 136 2028 1305 2040
rect 188 1976 1253 2028
rect 136 1970 1305 1976
rect 85 1934 1357 1940
rect 85 1882 353 1934
rect 405 1882 1037 1934
rect 1089 1882 1357 1934
rect 85 1870 1357 1882
rect 85 1818 353 1870
rect 405 1818 1037 1870
rect 1089 1818 1357 1870
rect 85 1812 1357 1818
rect 85 1462 241 1812
tri 241 1783 270 1812 nw
tri 1171 1783 1200 1812 ne
rect 1200 1783 1357 1812
tri 1200 1782 1201 1783 ne
tri 558 1766 564 1772 se
rect 564 1766 1044 1772
tri 533 1741 558 1766 se
rect 558 1741 565 1766
rect 533 1714 565 1741
rect 617 1714 825 1766
rect 877 1714 1044 1766
rect 533 1702 1044 1714
rect 533 1650 565 1702
rect 617 1650 825 1702
rect 877 1650 1044 1702
rect 533 1644 1044 1650
tri 490 1566 533 1609 se
rect 533 1566 622 1644
tri 622 1616 650 1644 nw
tri 951 1616 979 1644 ne
rect 979 1616 1044 1644
tri 979 1609 986 1616 ne
rect 986 1609 1044 1616
tri 986 1603 992 1609 ne
rect 85 1410 91 1462
rect 143 1410 183 1462
rect 235 1410 241 1462
rect 405 1494 622 1566
rect 992 1544 1044 1609
rect 405 1472 600 1494
tri 600 1472 622 1494 nw
rect 870 1516 922 1522
tri 855 1472 870 1487 se
rect 405 1469 483 1472
tri 483 1469 486 1472 nw
tri 852 1469 855 1472 se
rect 855 1469 870 1472
rect 405 1464 478 1469
tri 478 1464 483 1469 nw
tri 847 1464 852 1469 se
rect 852 1464 870 1469
rect 405 1463 466 1464
rect 457 1452 466 1463
tri 466 1452 478 1464 nw
tri 835 1452 847 1464 se
rect 847 1452 922 1464
tri 457 1443 466 1452 nw
tri 826 1443 835 1452 se
rect 835 1443 870 1452
tri 825 1442 826 1443 se
rect 826 1442 870 1443
tri 824 1441 825 1442 se
rect 825 1441 870 1442
rect 405 1399 457 1411
rect 405 1341 457 1347
rect 520 1435 870 1441
rect 572 1400 870 1435
rect 992 1480 1044 1492
rect 1201 1543 1357 1783
rect 1201 1491 1207 1543
rect 1259 1491 1299 1543
rect 1351 1491 1357 1543
rect 992 1422 1044 1428
rect 572 1394 922 1400
rect 520 1371 572 1383
tri 572 1349 617 1394 nw
rect 520 1313 572 1319
rect 940 1280 992 1286
tri 908 1228 940 1260 se
tri 894 1214 908 1228 se
rect 908 1214 992 1228
rect 75 1162 81 1214
rect 133 1162 154 1214
rect 206 1162 212 1214
rect 268 1162 274 1214
rect 326 1162 338 1214
rect 390 1162 402 1214
rect 454 1162 466 1214
rect 518 1211 524 1214
tri 524 1211 527 1214 sw
tri 891 1211 894 1214 se
rect 894 1211 940 1214
rect 518 1165 940 1211
rect 518 1162 524 1165
tri 524 1162 527 1165 nw
tri 931 1162 934 1165 ne
rect 934 1162 940 1165
tri 44 1131 75 1162 se
rect 75 1156 212 1162
tri 212 1156 218 1162 sw
tri 934 1156 940 1162 ne
rect 940 1156 992 1162
rect 1090 1280 1142 1286
rect 1090 1214 1142 1228
rect 75 1131 218 1156
rect 44 1130 218 1131
tri 218 1130 244 1156 sw
tri 1064 1130 1090 1156 se
rect 1090 1130 1142 1162
rect 44 1128 894 1130
tri 894 1128 896 1130 sw
tri 1062 1128 1064 1130 se
rect 1064 1128 1142 1130
rect 44 1079 1142 1128
rect 44 53 82 1079
tri 82 1042 119 1079 nw
rect 214 1026 930 1032
rect 266 974 526 1026
rect 578 974 814 1026
rect 866 974 878 1026
rect 214 938 930 974
rect 266 886 526 938
rect 578 886 814 938
rect 866 886 878 938
rect 214 880 930 886
rect 121 825 774 831
rect 173 773 370 825
rect 422 773 658 825
rect 710 773 722 825
rect 121 737 774 773
rect 173 685 370 737
rect 422 685 658 737
rect 710 685 722 737
rect 121 679 774 685
use sky130_fd_pr__nfet_01v8__example_55959141808546  sky130_fd_pr__nfet_01v8__example_55959141808546_1
timestamp 1619862920
transform -1 0 1035 0 -1 2182
box -28 0 78 267
use sky130_fd_pr__nfet_01v8__example_55959141808546  sky130_fd_pr__nfet_01v8__example_55959141808546_0
timestamp 1619862920
transform -1 0 929 0 -1 2182
box -28 0 78 267
use sky130_fd_pr__nfet_01v8__example_55959141808547  sky130_fd_pr__nfet_01v8__example_55959141808547_0
timestamp 1619862920
transform -1 0 1357 0 -1 2182
box -28 0 184 267
use sky130_fd_pr__pfet_01v8__example_55959141808545  sky130_fd_pr__pfet_01v8__example_55959141808545_0
timestamp 1619862920
transform 1 0 112 0 1 123
box -28 0 440 471
use sky130_fd_pr__pfet_01v8__example_55959141808543  sky130_fd_pr__pfet_01v8__example_55959141808543_0
timestamp 1619862920
transform 1 0 84 0 1 1501
box -28 0 184 471
use sky130_fd_pr__pfet_01v8__example_55959141808544  sky130_fd_pr__pfet_01v8__example_55959141808544_1
timestamp 1619862920
transform 1 0 407 0 1 1501
box -28 0 78 471
use sky130_fd_pr__pfet_01v8__example_55959141808544  sky130_fd_pr__pfet_01v8__example_55959141808544_0
timestamp 1619862920
transform 1 0 513 0 1 1501
box -28 0 78 471
use sky130_fd_pr__nfet_01v8__example_55959141808533  sky130_fd_pr__nfet_01v8__example_55959141808533_1
timestamp 1619862920
transform -1 0 1014 0 1 123
box -28 0 128 471
use sky130_fd_pr__nfet_01v8__example_55959141808533  sky130_fd_pr__nfet_01v8__example_55959141808533_0
timestamp 1619862920
transform -1 0 1170 0 1 123
box -28 0 128 471
<< labels >>
flabel metal2 s 983 1844 1106 1920 3 FreeSans 520 0 0 0 OUT_B
port 1 nsew
flabel metal2 s 1008 1992 1118 2067 3 FreeSans 520 0 0 0 OUT
port 2 nsew
flabel metal2 s 89 1150 183 1201 3 FreeSans 520 0 0 0 ENABLE_VDDIO_LV
port 3 nsew
flabel comment s 783 1702 783 1702 0 FreeSans 200 0 0 0 FBK
flabel comment s 837 1298 837 1298 0 FreeSans 200 90 0 0 FBK_N
flabel comment s 381 2593 381 2593 0 FreeSans 600 0 0 0 LV_NET
flabel metal1 s 1399 1064 1483 1129 3 FreeSans 520 0 0 0 VSSD
port 4 nsew
flabel metal1 s 258 2538 420 2602 3 FreeSans 200 0 0 0 VCCHIB
port 5 nsew
flabel metal1 s 955 1180 980 1265 3 FreeSans 200 0 0 0 IN
port 6 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 36200652
string GDS_START 36163832
<< end >>
