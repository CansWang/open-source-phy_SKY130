module term_res_flat (
    input IN,
    output OUT
);
    
endmodule