**** Created by MC2: Version 2013.12.00.f on 2020/05/11, 12:57:43 

************************************************************************
* auCdl Netlist:
* 
* Library Name:  N16_HDSPSB_LEAFCELL
* Top Cell Name: LEAFCELL_TILING
* View Name:     schematic
* Netlisted on:  Oct  2 11:11:16 2014
************************************************************************

*.BIPOLAR
*.CAPA
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.PARAM

.SUBCKT ndio_mac PLUS MINUS 
*.PININFO 
.ENDS

*.PIN vss

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    DIODE
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_DIODE TSMC_1 TSMC_2 VSS 
*.PININFO  TSMC_1:I TSMC_2:B VSS:B 
MMDIODE TSMC_1 TSMC_2 TSMC_1 VSS nch_lvt_mac l=20n nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: simLib

* View Name:    schematic
************************************************************************



************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    XDRV_LA512_884_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_XDRV_LA512_884_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 
*.PININFO  TSMC_30:I TSMC_31:I TSMC_22:O TSMC_23:O TSMC_24:O TSMC_25:O 
*.PININFO  TSMC_26:O TSMC_27:O TSMC_28:O TSMC_29:O TSMC_1:B 
*.PININFO  TSMC_2:B TSMC_3:B TSMC_4:B TSMC_5:B TSMC_6:B 
*.PININFO  TSMC_7:B TSMC_8:B TSMC_9:B TSMC_10:B TSMC_11:B 
*.PININFO  TSMC_12:B TSMC_13:B TSMC_14:B TSMC_15:B TSMC_16:B 
*.PININFO  TSMC_17:B TSMC_18:B TSMC_19:B TSMC_20:B TSMC_21:B 
MM37 TSMC_28 TSMC_32 TSMC_20 TSMC_20 pch_svt_mac l=20n nfin=8 m=8 
MM36 TSMC_32 TSMC_30 TSMC_20 TSMC_20 pch_lvt_mac l=20n nfin=7 m=1 
MM35 TSMC_24 TSMC_32 TSMC_20 TSMC_20 pch_svt_mac l=20n nfin=8 m=8 
MM34 TSMC_32 TSMC_33 TSMC_20 TSMC_20 pch_lvt_mac l=20n nfin=7 m=1 
MM33 TSMC_33 TSMC_3 TSMC_34 TSMC_20 pch_lvt_mac l=20n nfin=7 m=1 
MM21 TSMC_29 TSMC_35 TSMC_20 TSMC_20 pch_svt_mac l=20n nfin=8 m=8 
MM16 TSMC_35 TSMC_30 TSMC_20 TSMC_20 pch_lvt_mac l=20n nfin=7 m=1 
MM13 TSMC_25 TSMC_35 TSMC_20 TSMC_20 pch_svt_mac l=20n nfin=8 m=8 
MM11 TSMC_35 TSMC_36 TSMC_20 TSMC_20 pch_lvt_mac l=20n nfin=7 m=1 
MM10 TSMC_36 TSMC_4 TSMC_34 TSMC_20 pch_lvt_mac l=20n nfin=7 m=1 
MM3 TSMC_27 TSMC_37 TSMC_20 TSMC_20 pch_svt_mac l=20n nfin=8 m=8 
MM2 TSMC_26 TSMC_38 TSMC_20 TSMC_20 pch_svt_mac l=20n nfin=8 m=8 
MM23 TSMC_23 TSMC_37 TSMC_20 TSMC_20 pch_svt_mac l=20n nfin=8 m=8 
MM20 TSMC_22 TSMC_38 TSMC_20 TSMC_20 pch_svt_mac l=20n nfin=8 m=8 
MM28 TSMC_37 TSMC_30 TSMC_20 TSMC_20 pch_lvt_mac l=20n nfin=7 m=1 
MM27 TSMC_38 TSMC_30 TSMC_20 TSMC_20 pch_lvt_mac l=20n nfin=7 m=1 
MM26 TSMC_37 TSMC_39 TSMC_20 TSMC_20 pch_lvt_mac l=20n nfin=7 m=1 
MM18 TSMC_38 TSMC_40 TSMC_20 TSMC_20 pch_lvt_mac l=20n nfin=7 m=1 
MM12 TSMC_39 TSMC_2 TSMC_34 TSMC_20 pch_lvt_mac l=20n nfin=7 m=1 
MP6 TSMC_40 TSMC_1 TSMC_34 TSMC_20 pch_lvt_mac l=20n nfin=7 m=1 
MM39 TSMC_34 TSMC_9 TSMC_20 TSMC_20 pch_lvt_mac l=20n nfin=7 m=4 
MM32 TSMC_28 TSMC_32 TSMC_21 TSMC_21 nch_lvt_mac l=20n nfin=10 m=4 
MM31 TSMC_24 TSMC_32 TSMC_21 TSMC_21 nch_lvt_mac l=20n nfin=10 m=4 
MM30 TSMC_32 TSMC_33 TSMC_31 TSMC_21 nch_lvt_mac l=20n nfin=12 m=1 
MM29 TSMC_33 TSMC_9 TSMC_21 TSMC_21 nch_lvt_mac l=20n nfin=3 m=1 
MM22 TSMC_33 TSMC_3 TSMC_21 TSMC_21 nch_lvt_mac l=20n nfin=3 m=1 
MM9 TSMC_29 TSMC_35 TSMC_21 TSMC_21 nch_lvt_mac l=20n nfin=10 m=4 
MM8 TSMC_25 TSMC_35 TSMC_21 TSMC_21 nch_lvt_mac l=20n nfin=10 m=4 
MM7 TSMC_35 TSMC_36 TSMC_31 TSMC_21 nch_lvt_mac l=20n nfin=12 m=1 
MM5 TSMC_36 TSMC_9 TSMC_21 TSMC_21 nch_lvt_mac l=20n nfin=3 m=1 
MM4 TSMC_36 TSMC_4 TSMC_21 TSMC_21 nch_lvt_mac l=20n nfin=3 m=1 
MM1 TSMC_27 TSMC_37 TSMC_21 TSMC_21 nch_lvt_mac l=20n nfin=10 m=4 
MM0 TSMC_26 TSMC_38 TSMC_21 TSMC_21 nch_lvt_mac l=20n nfin=10 m=4 
MM24 TSMC_23 TSMC_37 TSMC_21 TSMC_21 nch_lvt_mac l=20n nfin=10 m=4 
MM19 TSMC_22 TSMC_38 TSMC_21 TSMC_21 nch_lvt_mac l=20n nfin=10 m=4 
MM25 TSMC_37 TSMC_39 TSMC_31 TSMC_21 nch_lvt_mac l=20n nfin=12 m=1 
MM17 TSMC_38 TSMC_40 TSMC_31 TSMC_21 nch_lvt_mac l=20n nfin=12 m=1 
MM14 TSMC_39 TSMC_9 TSMC_21 TSMC_21 nch_lvt_mac l=20n nfin=3 m=1 
MM6 TSMC_40 TSMC_9 TSMC_21 TSMC_21 nch_lvt_mac l=20n nfin=3 m=1 
MM15 TSMC_39 TSMC_2 TSMC_21 TSMC_21 nch_lvt_mac l=20n nfin=3 m=1 
MP9 TSMC_40 TSMC_1 TSMC_21 TSMC_21 nch_lvt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    BCELL_SD_HD
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_BCELL_SD_HD TSMC_1 TSMC_2 VDDAI TSMC_3 TSMC_4 TSMC_5 
*.PININFO  TSMC_1:B TSMC_2:B VDDAI:B TSMC_3:B TSMC_4:B TSMC_5:B 
MM5 TSMC_2 TSMC_5 TSMC_6 TSMC_4 nchpg_hdsr_mac l=20n nfin=1 m=1 
MM0 TSMC_1 TSMC_5 TSMC_7 TSMC_4 nchpg_hdsr_mac l=20n nfin=1 m=1 
MM2 TSMC_6 TSMC_7 TSMC_4 TSMC_4 nchpd_hdsr_mac l=20n nfin=1 m=1 
MM1 TSMC_7 TSMC_6 TSMC_4 TSMC_4 nchpd_hdsr_mac l=20n nfin=1 m=1 
MM6 TSMC_7 TSMC_6 VDDAI TSMC_3 pchpu_hdsr_mac l=20n nfin=1 m=1 
MM4 TSMC_6 TSMC_7 VDDAI TSMC_3 pchpu_hdsr_mac l=20n nfin=1 m=1 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    MCB_2X4_SD_HD
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_MCB_2X4_SD_HD TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
*.PININFO  TSMC_1:B TSMC_2:B TSMC_3:B TSMC_4:B TSMC_5:B TSMC_6:B TSMC_7:B 
*.PININFO  TSMC_8:B 
*.PININFO  TSMC_9:B TSMC_10:B TSMC_11:B TSMC_12:B TSMC_13:B TSMC_14:B TSMC_15:B 
*.PININFO  TSMC_16:B 
XMCB_0[0] TSMC_1 TSMC_5 TSMC_9 TSMC_13 TSMC_14 TSMC_15 
+ S1CSLVTSW400W90_BCELL_SD_HD 
XMCB_0[1] TSMC_2 TSMC_6 TSMC_10 TSMC_13 TSMC_14 TSMC_15 
+ S1CSLVTSW400W90_BCELL_SD_HD 
XMCB_0[2] TSMC_3 TSMC_7 TSMC_11 TSMC_13 TSMC_14 TSMC_15 
+ S1CSLVTSW400W90_BCELL_SD_HD 
XMCB_0[3] TSMC_4 TSMC_8 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ S1CSLVTSW400W90_BCELL_SD_HD 
XMCB_1[0] TSMC_1 TSMC_5 TSMC_9 TSMC_13 TSMC_14 TSMC_16 
+ S1CSLVTSW400W90_BCELL_SD_HD 
XMCB_1[1] TSMC_2 TSMC_6 TSMC_10 TSMC_13 TSMC_14 TSMC_16 
+ S1CSLVTSW400W90_BCELL_SD_HD 
XMCB_1[2] TSMC_3 TSMC_7 TSMC_11 TSMC_13 TSMC_14 TSMC_16 
+ S1CSLVTSW400W90_BCELL_SD_HD 
XMCB_1[3] TSMC_4 TSMC_8 TSMC_12 TSMC_13 TSMC_14 TSMC_16 
+ S1CSLVTSW400W90_BCELL_SD_HD 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    inv_lvt_mac_pcell_0
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_inv_lvt_mac_pcell_0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_5:I TSMC_6:I TSMC_4:O 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    inv_svt_mac_pcell_0
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_inv_svt_mac_pcell_0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_5:I TSMC_6:I TSMC_4:O 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand2_lvt_mac_pcell_1
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:O 
MM2 TSMC_7 TSMC_2 TSMC_5 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_7 TSMC_1 TSMC_5 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_8 TSMC_2 TSMC_3 TSMC_4 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_8 TSMC_4 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand2_svt_mac_pcell_1
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_nand2_svt_mac_pcell_1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:O 
MM2 TSMC_7 TSMC_2 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_7 TSMC_1 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_8 TSMC_2 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_8 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand3_lvt_mac_pcell_2
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_nand3_lvt_mac_pcell_2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:I 
*.PININFO  TSMC_8:O 
MM3 TSMC_8 TSMC_3 TSMC_6 TSMC_7 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_8 TSMC_2 TSMC_6 TSMC_7 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_6 TSMC_7 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM6 TSMC_9 TSMC_3 TSMC_4 TSMC_5 nch_lvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM5 TSMC_10 TSMC_2 TSMC_9 TSMC_5 nch_lvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM4 TSMC_8 TSMC_1 TSMC_10 TSMC_5 nch_lvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    WEBBUF_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_WEBBUF_SB_BASE TSMC_1 TSMC_2 VDDHD TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_5:I TSMC_6:O TSMC_7:O VDDHD:B TSMC_3:B 
*.PININFO  TSMC_4:B 
MM36 TSMC_8 TSMC_9 TSMC_4 TSMC_4 nch_lvt_mac l=20n nfin=3 m=1 
MM35 TSMC_10 TSMC_2 TSMC_8 TSMC_4 nch_lvt_mac l=20n nfin=3 m=1 
MM31 TSMC_11 TSMC_1 TSMC_4 TSMC_4 nch_lvt_mac l=20n nfin=5 m=2 
MM30 TSMC_10 TSMC_5 TSMC_11 TSMC_4 nch_lvt_mac l=20n nfin=5 m=1 
MM34 TSMC_12 TSMC_9 VDDHD TSMC_3 pch_lvt_mac l=20n nfin=3 m=1 
MM33 TSMC_10 TSMC_1 TSMC_12 TSMC_3 pch_lvt_mac l=20n nfin=3 m=1 
MM6 TSMC_10 TSMC_5 TSMC_13 TSMC_3 pch_lvt_mac l=20n nfin=5 m=1 
MM32 TSMC_13 TSMC_2 VDDHD TSMC_3 pch_lvt_mac l=20n nfin=5 m=2 
XI25 TSMC_4 TSMC_4 TSMC_10 TSMC_9 VDDHD TSMC_3 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI32 TSMC_4 TSMC_4 TSMC_10 TSMC_7 VDDHD TSMC_3 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=2 n_nfin=4 n_l=20n p_totalM=2 
+ p_nfin=7 p_l=20n 
XI33 TSMC_4 TSMC_4 TSMC_7 TSMC_6 VDDHD TSMC_3 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=7 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    RESETD_TSEL
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_RESETD_TSEL TSMC_1 TSMC_2 TSMC_3 VDDHD TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_6:O TSMC_7:O VDDHD:B TSMC_4:B 
*.PININFO  TSMC_5:B 
MM15 TSMC_8 TSMC_1 TSMC_9 TSMC_4 pch_svt_mac l=20n nfin=3 m=1 
MM14 TSMC_9 TSMC_1 VDDHD TSMC_4 pch_svt_mac l=20n nfin=3 m=1 
MM25 TSMC_6 TSMC_2 VDDHD TSMC_4 pch_lvt_mac l=20n nfin=3 m=1 
MM23 TSMC_6 TSMC_10 VDDHD TSMC_4 pch_lvt_mac l=20n nfin=3 m=1 
MM18 TSMC_8 TSMC_1 TSMC_11 TSMC_5 nch_svt_mac l=20n nfin=3 m=1 
MM19 TSMC_11 TSMC_1 TSMC_5 TSMC_5 nch_svt_mac l=20n nfin=3 m=1 
MM24 TSMC_12 TSMC_10 TSMC_5 TSMC_5 nch_lvt_mac l=20n nfin=3 m=1 
MM21 TSMC_6 TSMC_2 TSMC_12 TSMC_5 nch_lvt_mac l=20n nfin=3 m=1 
XI737 TSMC_5 TSMC_5 TSMC_13 TSMC_7 VDDHD TSMC_4 
+ S1CSLVTSW400W90_inv_svt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI736 TSMC_5 TSMC_5 TSMC_14 TSMC_13 VDDHD TSMC_4 
+ S1CSLVTSW400W90_inv_svt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XND0 TSMC_1 TSMC_7 TSMC_5 TSMC_5 VDDHD TSMC_4 TSMC_10 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI91 TSMC_3 TSMC_8 TSMC_5 TSMC_5 VDDHD TSMC_4 TSMC_14 
+ S1CSLVTSW400W90_nand2_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    RESETD_WTSEL_SB_NEW
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_RESETD_WTSEL_SB_NEW TSMC_1 TSMC_2 VDDHD TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 
*.PININFO  TSMC_1:I TSMC_5:I TSMC_6:I TSMC_2:O VDDHD:B TSMC_3:B TSMC_4:B 
XI87 TSMC_7 TSMC_8 TSMC_4 TSMC_4 VDDHD TSMC_3 TSMC_9 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XND5 TSMC_6 TSMC_10 TSMC_4 TSMC_4 VDDHD TSMC_3 TSMC_7 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI84 TSMC_5 TSMC_11 TSMC_4 TSMC_4 VDDHD TSMC_3 TSMC_8 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XND0 TSMC_7 TSMC_1 TSMC_4 TSMC_4 VDDHD TSMC_3 TSMC_11 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI89 TSMC_4 TSMC_4 TSMC_9 TSMC_2 VDDHD TSMC_3 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI65 TSMC_4 TSMC_4 TSMC_12 TSMC_13 VDDHD TSMC_3 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI83 TSMC_4 TSMC_4 TSMC_13 TSMC_10 VDDHD TSMC_3 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI64 TSMC_4 TSMC_4 TSMC_1 TSMC_12 VDDHD TSMC_3 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    DECB1_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_DECB1_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 VDDHD TSMC_8 TSMC_9 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:I TSMC_3:O 
*.PININFO  VDDHD:B TSMC_8:B TSMC_9:B 
MTN1 TSMC_10 TSMC_1 TSMC_11 TSMC_9 nch_lvt_mac l=20n nfin=3 m=1 
MTN2 TSMC_11 TSMC_7 TSMC_5 TSMC_9 nch_lvt_mac l=20n nfin=7 m=2 
MM0 TSMC_10 TSMC_2 TSMC_11 TSMC_9 nch_lvt_mac l=20n nfin=7 m=2 
MN0 TSMC_3 TSMC_10 TSMC_9 TSMC_9 nch_lvt_mac l=20n nfin=8 m=4 
MM1 TSMC_12 TSMC_2 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=1 
MM3 TSMC_10 TSMC_7 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=1 
MP0 TSMC_3 TSMC_10 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=8 m=6 
MP5 TSMC_10 TSMC_4 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=2 
MM2 TSMC_10 TSMC_1 TSMC_12 TSMC_8 pch_lvt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    DECB1_BLEQ_SB_M4
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_DECB1_BLEQ_SB_M4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 VDDHD TSMC_7 TSMC_8 
*.PININFO  TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_1:O TSMC_2:O VDDHD:B 
*.PININFO  TSMC_7:B TSMC_8:B 
MN0 TSMC_1 TSMC_9 TSMC_8 TSMC_8 nch_lvt_mac l=20n nfin=8 m=4 
MTN1 TSMC_9 TSMC_3 TSMC_6 TSMC_8 nch_lvt_mac l=20n nfin=3 m=1 
MM0 TSMC_9 TSMC_4 TSMC_6 TSMC_8 nch_lvt_mac l=20n nfin=6 m=2 
MM2 TSMC_2 TSMC_9 TSMC_8 TSMC_8 nch_lvt_mac l=20n nfin=8 m=4 
MP0 TSMC_1 TSMC_9 VDDHD TSMC_7 pch_lvt_mac l=20n nfin=8 m=6 
MM4 TSMC_9 TSMC_5 VDDHD TSMC_7 pch_lvt_mac l=20n nfin=3 m=2 
MM3 TSMC_9 TSMC_3 TSMC_10 TSMC_7 pch_lvt_mac l=20n nfin=3 m=1 
MM1 TSMC_10 TSMC_4 VDDHD TSMC_7 pch_lvt_mac l=20n nfin=3 m=1 
MM5 TSMC_2 TSMC_9 VDDHD TSMC_7 pch_lvt_mac l=20n nfin=8 m=6 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    DECB1_WLNAD2_SB_X0
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_DECB1_WLNAD2_SB_X0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 VDDHD TSMC_8 TSMC_9 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:I TSMC_3:O 
*.PININFO  VDDHD:B TSMC_8:B TSMC_9:B 
MM5 TSMC_10 TSMC_11 TSMC_9 TSMC_9 nch_lvt_mac l=20n nfin=6 m=1 
MTN1 TSMC_11 TSMC_1 TSMC_12 TSMC_9 nch_lvt_mac l=20n nfin=3 m=1 
MTN2 TSMC_12 TSMC_7 TSMC_5 TSMC_9 nch_lvt_mac l=20n nfin=6 m=2 
MM0 TSMC_11 TSMC_2 TSMC_12 TSMC_9 nch_lvt_mac l=20n nfin=6 m=2 
MN0 TSMC_3 TSMC_10 TSMC_9 TSMC_9 nch_lvt_mac l=20n nfin=8 m=6 
MM4 TSMC_10 TSMC_11 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=4 
MM1 TSMC_13 TSMC_2 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=1 
MM3 TSMC_11 TSMC_7 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=1 
MP0 TSMC_3 TSMC_10 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=8 m=3 
MP5 TSMC_11 TSMC_4 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=2 
MM2 TSMC_11 TSMC_1 TSMC_13 TSMC_8 pch_lvt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    CKBUF_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_CKBUF_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDDHD TSMC_5 
+ TSMC_6 
*.PININFO  TSMC_3:I TSMC_4:I TSMC_1:O TSMC_2:O VDDHD:B TSMC_5:B TSMC_6:B 
XINV0 TSMC_6 TSMC_6 TSMC_1 TSMC_2 VDDHD TSMC_5 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=2 n_nfin=7 n_l=20n p_totalM=3 
+ p_nfin=9 p_l=20n 
MM1 TSMC_1 TSMC_3 TSMC_6 TSMC_6 nch_lvt_mac l=20n nfin=3 m=1 
MM34 TSMC_1 TSMC_4 TSMC_6 TSMC_6 nch_lvt_mac l=20n nfin=7 m=2 
MM26 TSMC_7 TSMC_3 VDDHD TSMC_5 pch_lvt_mac l=20n nfin=9 m=2 
MM0 TSMC_1 TSMC_4 TSMC_7 TSMC_5 pch_lvt_mac l=20n nfin=9 m=2 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    ABUF_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_ABUF_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDDM 
+ VDDMHD TSMC_6 
*.PININFO  TSMC_1:I TSMC_4:I TSMC_5:I TSMC_2:O TSMC_3:O VDDM:B VDDMHD:B 
*.PININFO  TSMC_6:B 
MM15 TSMC_7 TSMC_8 TSMC_6 TSMC_6 nch_lvt_mac l=20n nfin=3 m=1 
MM14 TSMC_3 TSMC_5 TSMC_7 TSMC_6 nch_lvt_mac l=20n nfin=3 m=1 
MM9 TSMC_9 TSMC_4 TSMC_6 TSMC_6 nch_lvt_mac l=20n nfin=4 m=1 
MM8 TSMC_3 TSMC_1 TSMC_9 TSMC_6 nch_lvt_mac l=20n nfin=4 m=1 
MM13 TSMC_10 TSMC_8 VDDMHD VDDM pch_lvt_mac l=20n nfin=3 m=1 
MM12 TSMC_3 TSMC_4 TSMC_10 VDDM pch_lvt_mac l=20n nfin=3 m=1 
MM11 TSMC_3 TSMC_1 TSMC_11 VDDM pch_lvt_mac l=20n nfin=5 m=1 
MM10 TSMC_11 TSMC_5 VDDMHD VDDM pch_lvt_mac l=20n nfin=5 m=2 
XI34 TSMC_6 TSMC_6 TSMC_3 TSMC_8 VDDMHD VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI35 TSMC_6 TSMC_6 TSMC_3 TSMC_2 VDDMHD VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nor2_lvt_mac_pcell_4
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_nor2_lvt_mac_pcell_4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:O 
MM2 TSMC_7 TSMC_2 TSMC_8 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_5 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_7 TSMC_2 TSMC_3 TSMC_4 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_3 TSMC_4 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    ENBUFB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_ENBUFB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDDHD TSMC_9 TSMC_10 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_8:I TSMC_4:O TSMC_5:O TSMC_6:O 
*.PININFO  TSMC_7:O VDDHD:B TSMC_9:B 
*.PININFO  TSMC_10:B 
XI158 TSMC_11 TSMC_11 TSMC_10 TSMC_10 VDDHD TSMC_9 TSMC_12 
+ S1CSLVTSW400W90_nor2_lvt_mac_pcell_4 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
MM19 TSMC_13 TSMC_3 TSMC_9 TSMC_9 pch_lvt_mac l=20n nfin=6 m=1 
MM2 TSMC_14 TSMC_4 TSMC_9 TSMC_9 pch_lvt_mac l=20n nfin=3 m=1 
MM7 TSMC_15 TSMC_8 TSMC_9 TSMC_9 pch_lvt_mac l=20n nfin=5 m=1 
MM16 TSMC_15 TSMC_1 TSMC_13 TSMC_9 pch_lvt_mac l=20n nfin=6 m=1 
MM1 TSMC_15 TSMC_2 TSMC_14 TSMC_9 pch_lvt_mac l=20n nfin=3 m=1 
MM5 TSMC_16 TSMC_8 TSMC_10 TSMC_10 nch_lvt_mac l=20n nfin=3 m=1 
MN200 TSMC_6 TSMC_4 TSMC_10 TSMC_10 nch_lvt_mac l=20n nfin=7 m=2 
MM4 TSMC_17 TSMC_4 TSMC_16 TSMC_10 nch_lvt_mac l=20n nfin=3 m=1 
MM3 TSMC_15 TSMC_3 TSMC_17 TSMC_10 nch_lvt_mac l=20n nfin=3 m=1 
MM20 TSMC_18 TSMC_8 TSMC_10 TSMC_10 nch_lvt_mac l=20n nfin=7 m=1 
MM17 TSMC_15 TSMC_1 TSMC_19 TSMC_10 nch_lvt_mac l=20n nfin=4 m=1 
MM18 TSMC_19 TSMC_2 TSMC_18 TSMC_10 nch_lvt_mac l=20n nfin=4 m=1 
MN300 TSMC_5 TSMC_4 TSMC_10 TSMC_10 nch_lvt_mac l=20n nfin=11 m=6 
XI166 TSMC_10 TSMC_10 TSMC_20 TSMC_11 VDDHD TSMC_9 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI148 TSMC_10 TSMC_10 TSMC_4 TSMC_20 VDDHD TSMC_9 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI152 TSMC_10 TSMC_10 TSMC_21 TSMC_7 VDDHD TSMC_9 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=4 n_nfin=4 n_l=20n p_totalM=4 
+ p_nfin=8 p_l=20n 
XINV5 TSMC_10 TSMC_10 TSMC_4 TSMC_21 TSMC_9 TSMC_9 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=3 
+ p_nfin=3 p_l=20n 
XINV4 TSMC_10 TSMC_10 TSMC_12 TSMC_22 VDDHD TSMC_9 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI141 TSMC_10 TSMC_10 TSMC_15 TSMC_4 TSMC_9 TSMC_9 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=2 n_nfin=7 n_l=20n p_totalM=3 
+ p_nfin=9 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    DECB4_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_DECB4_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 VDDHD TSMC_10 TSMC_11 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:O TSMC_7:O 
*.PININFO  TSMC_8:O 
*.PININFO  TSMC_9:O VDDHD:B TSMC_10:B TSMC_11:B 
MM15 TSMC_12 TSMC_4 VDDHD TSMC_10 pch_lvt_mac l=20n nfin=3 m=1 
MM16 TSMC_12 TSMC_2 VDDHD TSMC_10 pch_lvt_mac l=20n nfin=3 m=1 
MM17 TSMC_13 TSMC_4 VDDHD TSMC_10 pch_lvt_mac l=20n nfin=3 m=1 
MM18 TSMC_13 TSMC_1 VDDHD TSMC_10 pch_lvt_mac l=20n nfin=3 m=1 
MM22 TSMC_13 TSMC_5 VDDHD TSMC_10 pch_lvt_mac l=20n nfin=3 m=1 
MM23 TSMC_12 TSMC_5 VDDHD TSMC_10 pch_lvt_mac l=20n nfin=3 m=1 
MM24 TSMC_14 TSMC_5 VDDHD TSMC_10 pch_lvt_mac l=20n nfin=3 m=1 
MM25 TSMC_15 TSMC_5 VDDHD TSMC_10 pch_lvt_mac l=20n nfin=3 m=1 
MM5 TSMC_14 TSMC_3 VDDHD TSMC_10 pch_lvt_mac l=20n nfin=3 m=1 
MM4 TSMC_14 TSMC_2 VDDHD TSMC_10 pch_lvt_mac l=20n nfin=3 m=1 
MM2 TSMC_15 TSMC_3 VDDHD TSMC_10 pch_lvt_mac l=20n nfin=3 m=1 
MM1 TSMC_15 TSMC_1 VDDHD TSMC_10 pch_lvt_mac l=20n nfin=3 m=1 
MM19 TSMC_16 TSMC_4 TSMC_17 TSMC_11 nch_lvt_mac l=20n nfin=3 m=2 
MM20 TSMC_12 TSMC_2 TSMC_16 TSMC_11 nch_lvt_mac l=20n nfin=3 m=1 
MM21 TSMC_13 TSMC_1 TSMC_16 TSMC_11 nch_lvt_mac l=20n nfin=3 m=1 
MM26 TSMC_17 TSMC_5 TSMC_11 TSMC_11 nch_lvt_mac l=20n nfin=3 m=4 
MM8 TSMC_18 TSMC_3 TSMC_17 TSMC_11 nch_lvt_mac l=20n nfin=3 m=2 
MM7 TSMC_14 TSMC_2 TSMC_18 TSMC_11 nch_lvt_mac l=20n nfin=3 m=1 
MM0 TSMC_15 TSMC_1 TSMC_18 TSMC_11 nch_lvt_mac l=20n nfin=3 m=1 
XINV3 TSMC_11 TSMC_11 TSMC_12 TSMC_9 VDDHD TSMC_10 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XINV2 TSMC_11 TSMC_11 TSMC_13 TSMC_8 VDDHD TSMC_10 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XINV1 TSMC_11 TSMC_11 TSMC_14 TSMC_7 VDDHD TSMC_10 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XINV0 TSMC_11 TSMC_11 TSMC_15 TSMC_6 VDDHD TSMC_10 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    DECB1_WLNAD2_SB_X1
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_DECB1_WLNAD2_SB_X1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 VDDHD TSMC_8 TSMC_9 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:I TSMC_3:O 
*.PININFO  VDDHD:B TSMC_8:B TSMC_9:B 
MM5 TSMC_10 TSMC_11 TSMC_9 TSMC_9 nch_lvt_mac l=20n nfin=6 m=1 
MTN1 TSMC_11 TSMC_1 TSMC_12 TSMC_9 nch_lvt_mac l=20n nfin=3 m=1 
MTN2 TSMC_12 TSMC_7 TSMC_5 TSMC_9 nch_lvt_mac l=20n nfin=6 m=2 
MM0 TSMC_11 TSMC_2 TSMC_12 TSMC_9 nch_lvt_mac l=20n nfin=6 m=2 
MN0 TSMC_3 TSMC_10 TSMC_9 TSMC_9 nch_lvt_mac l=20n nfin=8 m=6 
MM4 TSMC_10 TSMC_11 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=4 
MM1 TSMC_13 TSMC_2 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=1 
MM3 TSMC_11 TSMC_7 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=1 
MP0 TSMC_3 TSMC_10 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=8 m=3 
MP5 TSMC_11 TSMC_4 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=2 
MM2 TSMC_11 TSMC_1 TSMC_13 TSMC_8 pch_lvt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    DECB2_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_DECB2_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDDHD 
+ TSMC_6 TSMC_7 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:O TSMC_5:O VDDHD:B TSMC_6:B 
*.PININFO  TSMC_7:B 
MM2 TSMC_8 TSMC_3 VDDHD TSMC_6 pch_lvt_mac l=20n nfin=3 m=1 
MM1 TSMC_8 TSMC_1 VDDHD TSMC_6 pch_lvt_mac l=20n nfin=3 m=1 
MM5 TSMC_9 TSMC_3 VDDHD TSMC_6 pch_lvt_mac l=20n nfin=3 m=1 
MM4 TSMC_9 TSMC_2 VDDHD TSMC_6 pch_lvt_mac l=20n nfin=3 m=1 
MM0 TSMC_8 TSMC_1 TSMC_10 TSMC_7 nch_lvt_mac l=20n nfin=3 m=1 
MM7 TSMC_9 TSMC_2 TSMC_10 TSMC_7 nch_lvt_mac l=20n nfin=3 m=1 
MM8 TSMC_10 TSMC_3 TSMC_7 TSMC_7 nch_lvt_mac l=20n nfin=3 m=2 
XINV0 TSMC_7 TSMC_7 TSMC_9 TSMC_5 VDDHD TSMC_6 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XINV1 TSMC_7 TSMC_7 TSMC_8 TSMC_4 VDDHD TSMC_6 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    PRECHARGE_SB_SD
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_PRECHARGE_SB_SD TSMC_1 TSMC_2 TSMC_3 VDDAI TSMC_4 
*.PININFO  TSMC_3:I TSMC_1:B TSMC_2:B VDDAI:B TSMC_4:B 
MMPBLPRE VDDAI TSMC_3 TSMC_1 TSMC_4 pch_lvt_mac l=20n nfin=5 m=2 
MMPBLEQ TSMC_1 TSMC_3 TSMC_2 TSMC_4 pch_lvt_mac l=20n nfin=5 m=1 
MMPBLBPRE TSMC_2 TSMC_3 VDDAI TSMC_4 pch_lvt_mac l=20n nfin=5 m=2 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    MIO_M4_SB_NBL_S
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_MIO_M4_SB_NBL_S TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 VDDM VDDMHD TSMC_7 
*.PININFO  TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_1:B 
*.PININFO  TSMC_6:B VDDM:B VDDMHD:B TSMC_7:B 
MM12 TSMC_8 TSMC_6 TSMC_8 VDDM pch_lvt_mac l=20n nfin=11 m=4 
MM13 TSMC_9 TSMC_6 TSMC_9 VDDM pch_lvt_mac l=20n nfin=10 m=5 
MM14 TSMC_9 TSMC_6 TSMC_9 VDDM pch_lvt_mac l=20n nfin=10 m=4 
MM11 TSMC_8 TSMC_6 TSMC_8 VDDM pch_lvt_mac l=20n nfin=11 m=5 
MN34 TSMC_6 TSMC_10 TSMC_7 TSMC_7 nch_lvt_mac l=20n nfin=12 m=3 
MN33 TSMC_6 TSMC_10 TSMC_7 TSMC_7 nch_lvt_mac l=20n nfin=12 m=3 
XI8 TSMC_7 TSMC_7 TSMC_11 TSMC_8 VDDMHD VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=2 n_nfin=5 n_l=20n p_totalM=2 
+ p_nfin=5 p_l=20n 
XI16 TSMC_7 TSMC_7 TSMC_12 TSMC_10 VDDM VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=5 n_l=20n p_totalM=1 
+ p_nfin=5 p_l=20n 
XI1 TSMC_7 TSMC_7 TSMC_13 TSMC_14 VDDM VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
XI7 TSMC_7 TSMC_7 TSMC_14 TSMC_11 VDDMHD VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI17 TSMC_7 TSMC_7 TSMC_14 TSMC_12 VDDMHD VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
XI11 TSMC_7 TSMC_7 TSMC_14 TSMC_15 VDDMHD VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI9 TSMC_7 TSMC_7 TSMC_15 TSMC_9 VDDMHD VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=2 n_nfin=5 n_l=20n p_totalM=2 
+ p_nfin=5 p_l=20n 
XLD01 TSMC_7 TSMC_7 TSMC_2 TSMC_13 VDDMHD VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    LOGIC_D0734_TRKWL
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_LOGIC_D0734_TRKWL VSS TSMC_1 TSMC_2 
*.PININFO  VSS:B TSMC_1:B TSMC_2:B 
MMTRKWL1_PG VSS TSMC_1 VSS VSS nch_lvt_mac l=20n nfin=4 m=1 
MMTRKWL_PG VSS TSMC_1 VSS VSS nch_lvt_mac l=20n nfin=4 m=1 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    DECB1_DCLK_M4_SB_V2
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_DECB1_DCLK_M4_SB_V2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 VDDHD TSMC_8 TSMC_9 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_5:I TSMC_6:I TSMC_7:I TSMC_3:O TSMC_4:O 
*.PININFO  VDDHD:B TSMC_8:B TSMC_9:B 
MM2 TSMC_4 TSMC_10 TSMC_9 TSMC_9 nch_lvt_mac l=20n nfin=8 m=5 
MTN1 TSMC_10 TSMC_1 TSMC_11 TSMC_9 nch_lvt_mac l=20n nfin=3 m=1 
MTN2 TSMC_11 TSMC_7 TSMC_6 TSMC_9 nch_lvt_mac l=20n nfin=6 m=4 
MM0 TSMC_10 TSMC_2 TSMC_11 TSMC_9 nch_lvt_mac l=20n nfin=6 m=4 
MN0 TSMC_3 TSMC_10 TSMC_9 TSMC_9 nch_lvt_mac l=20n nfin=8 m=5 
MM4 TSMC_4 TSMC_10 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=8 m=8 
MM1 TSMC_12 TSMC_2 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=1 
MM3 TSMC_10 TSMC_7 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=1 
MP0 TSMC_3 TSMC_10 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=8 m=8 
MP5 TSMC_10 TSMC_5 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=2 
MM5 TSMC_10 TSMC_1 TSMC_12 TSMC_8 pch_lvt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    DECB1_Y_M4_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_DECB1_Y_M4_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 VDDHD TSMC_8 TSMC_9 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:I TSMC_3:O 
*.PININFO  VDDHD:B TSMC_8:B TSMC_9:B 
MM6 TSMC_10 TSMC_11 TSMC_9 TSMC_9 nch_lvt_mac l=20n nfin=6 m=1 
MN0 TSMC_3 TSMC_10 TSMC_9 TSMC_9 nch_lvt_mac l=20n nfin=9 m=9 
MTN1 TSMC_11 TSMC_1 TSMC_12 TSMC_9 nch_lvt_mac l=20n nfin=3 m=1 
MTN2 TSMC_12 TSMC_7 TSMC_5 TSMC_9 nch_lvt_mac l=20n nfin=6 m=2 
MM0 TSMC_11 TSMC_2 TSMC_12 TSMC_9 nch_lvt_mac l=20n nfin=6 m=2 
MM7 TSMC_10 TSMC_11 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=4 
MP0 TSMC_3 TSMC_10 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=7 m=6 
MM3 TSMC_11 TSMC_7 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=1 
MP5 TSMC_11 TSMC_4 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=2 
MM1 TSMC_13 TSMC_2 VDDHD TSMC_8 pch_lvt_mac l=20n nfin=3 m=1 
MM2 TSMC_11 TSMC_1 TSMC_13 TSMC_8 pch_lvt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    CDEC_M4_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_CDEC_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 VDDM VDDMHD TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 
+ TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 
+ TSMC_60 TSMC_61 
*.PININFO  TSMC_3:I TSMC_8:I TSMC_9:I TSMC_10:I TSMC_11:I TSMC_41:I TSMC_43:I 
*.PININFO  TSMC_46:I TSMC_47:I 
*.PININFO  TSMC_48:I TSMC_49:I TSMC_50:I TSMC_51:I TSMC_52:I TSMC_53:I 
*.PININFO  TSMC_54:I TSMC_55:I 
*.PININFO  TSMC_56:I TSMC_57:I TSMC_58:I TSMC_59:I TSMC_1:O TSMC_2:O TSMC_4:O 
*.PININFO  TSMC_5:O 
*.PININFO  TSMC_6:O TSMC_7:O TSMC_12:O TSMC_13:O TSMC_14:O TSMC_15:O 
*.PININFO  TSMC_16:O TSMC_17:O TSMC_18:O TSMC_19:O TSMC_20:O 
*.PININFO  TSMC_21:O TSMC_22:O TSMC_23:O TSMC_24:O TSMC_25:O 
*.PININFO  TSMC_26:O TSMC_27:O TSMC_28:O TSMC_29:O TSMC_30:O 
*.PININFO  TSMC_31:O TSMC_32:O TSMC_33:O TSMC_34:O TSMC_35:O 
*.PININFO  TSMC_36:O TSMC_37:O TSMC_38:O TSMC_39:O TSMC_40:O TSMC_42:O 
*.PININFO  TSMC_45:O 
*.PININFO  TSMC_60:O TSMC_61:O VDDM:B VDDMHD:B TSMC_44:B 
XIDEC_X2[0] TSMC_8 TSMC_10 TSMC_28 TSMC_40 TSMC_62 TSMC_41 TSMC_63 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_SB 
XIDEC_X2[1] TSMC_8 TSMC_10 TSMC_29 TSMC_40 TSMC_62 TSMC_41 TSMC_64 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_SB 
XIDEC_X2[2] TSMC_8 TSMC_10 TSMC_30 TSMC_40 TSMC_62 TSMC_41 TSMC_65 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_SB 
XIDEC_X2[3] TSMC_8 TSMC_10 TSMC_31 TSMC_40 TSMC_62 TSMC_41 TSMC_66 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_SB 
XDECB1_BLEQ TSMC_1 TSMC_2 TSMC_9 TSMC_10 TSMC_67 TSMC_68 VDDMHD VDDM TSMC_44 
+ S1CSLVTSW400W90_DECB1_BLEQ_SB_M4 
XIDEC_X0[0] TSMC_9 TSMC_10 TSMC_12 TSMC_67 TSMC_68 TSMC_41 TSMC_69 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_WLNAD2_SB_X0 
XIDEC_X0[1] TSMC_9 TSMC_10 TSMC_13 TSMC_67 TSMC_68 TSMC_41 TSMC_70 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_WLNAD2_SB_X0 
XIDEC_X0[2] TSMC_9 TSMC_10 TSMC_14 TSMC_67 TSMC_68 TSMC_41 TSMC_71 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_WLNAD2_SB_X0 
XIDEC_X0[3] TSMC_9 TSMC_10 TSMC_15 TSMC_67 TSMC_68 TSMC_41 TSMC_72 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_WLNAD2_SB_X0 
XIDEC_X0[4] TSMC_9 TSMC_10 TSMC_16 TSMC_67 TSMC_68 TSMC_41 TSMC_73 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_WLNAD2_SB_X0 
XIDEC_X0[5] TSMC_9 TSMC_10 TSMC_17 TSMC_67 TSMC_68 TSMC_41 TSMC_74 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_WLNAD2_SB_X0 
XIDEC_X0[6] TSMC_9 TSMC_10 TSMC_18 TSMC_67 TSMC_68 TSMC_41 TSMC_75 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_WLNAD2_SB_X0 
XIDEC_X0[7] TSMC_9 TSMC_10 TSMC_19 TSMC_67 TSMC_68 TSMC_41 TSMC_76 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_WLNAD2_SB_X0 
XPREDEC_Y[0] TSMC_77 TSMC_78 TSMC_79 TSMC_80 TSMC_46 TSMC_81 TSMC_82 TSMC_83 
+ TSMC_84 VDDMHD VDDM TSMC_44 S1CSLVTSW400W90_DECB4_SB 
XPREDEC_Y[1] TSMC_77 TSMC_78 TSMC_79 TSMC_80 TSMC_47 TSMC_85 TSMC_86 TSMC_87 
+ TSMC_88 VDDMHD VDDM TSMC_44 S1CSLVTSW400W90_DECB4_SB 
XIPDEC_X1[0] TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 
+ TSMC_97 VDDMHD VDDM TSMC_44 S1CSLVTSW400W90_DECB4_SB 
XIPDEC_X1[1] TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_98 TSMC_99 TSMC_100 TSMC_101 
+ TSMC_102 VDDMHD VDDM TSMC_44 S1CSLVTSW400W90_DECB4_SB 
XIPDEC_X0[0] TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 VDDMHD VDDM TSMC_44 S1CSLVTSW400W90_DECB4_SB 
XIPDEC_X0[1] TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_108 TSMC_73 TSMC_74 
+ TSMC_75 TSMC_76 VDDMHD VDDM TSMC_44 S1CSLVTSW400W90_DECB4_SB 
XCKBUF TSMC_4 TSMC_5 TSMC_9 TSMC_11 VDDMHD VDDM TSMC_44 
+ S1CSLVTSW400W90_CKBUF_SB 
XABUF_Y[0] TSMC_56 TSMC_77 TSMC_78 TSMC_4 TSMC_5 VDDM VDDMHD TSMC_44 
+ S1CSLVTSW400W90_ABUF_SB_BASE 
XABUF_Y[1] TSMC_57 TSMC_79 TSMC_80 TSMC_4 TSMC_5 VDDM VDDMHD TSMC_44 
+ S1CSLVTSW400W90_ABUF_SB_BASE 
XABUF_X[3] TSMC_51 TSMC_89 TSMC_90 TSMC_4 TSMC_5 VDDM VDDMHD TSMC_44 
+ S1CSLVTSW400W90_ABUF_SB_BASE 
XABUF_X[4] TSMC_52 TSMC_91 TSMC_92 TSMC_4 TSMC_5 VDDM VDDMHD TSMC_44 
+ S1CSLVTSW400W90_ABUF_SB_BASE 
XABUF_X[5] TSMC_53 TSMC_93 TSMC_98 TSMC_4 TSMC_5 VDDM VDDMHD TSMC_44 
+ S1CSLVTSW400W90_ABUF_SB_BASE 
XABUF_X[6] TSMC_54 TSMC_109 TSMC_110 TSMC_4 TSMC_5 VDDM VDDMHD TSMC_44 
+ S1CSLVTSW400W90_ABUF_SB_BASE 
XABUF_X[7] TSMC_55 TSMC_111 TSMC_112 TSMC_4 TSMC_5 VDDM VDDMHD TSMC_44 
+ S1CSLVTSW400W90_ABUF_SB_BASE 
XABUF_X[0] TSMC_48 TSMC_103 TSMC_104 TSMC_4 TSMC_5 VDDM VDDMHD TSMC_44 
+ S1CSLVTSW400W90_ABUF_SB_BASE 
XABUF_X[1] TSMC_49 TSMC_105 TSMC_106 TSMC_4 TSMC_5 VDDM VDDMHD TSMC_44 
+ S1CSLVTSW400W90_ABUF_SB_BASE 
XABUF_X[2] TSMC_50 TSMC_107 TSMC_108 TSMC_4 TSMC_5 VDDM VDDMHD TSMC_44 
+ S1CSLVTSW400W90_ABUF_SB_BASE 
XIDEC_Y[0] TSMC_9 TSMC_10 TSMC_32 TSMC_67 TSMC_68 TSMC_41 TSMC_81 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_Y_M4_SB 
XIDEC_Y[1] TSMC_9 TSMC_10 TSMC_33 TSMC_67 TSMC_68 TSMC_41 TSMC_82 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_Y_M4_SB 
XIDEC_Y[2] TSMC_9 TSMC_10 TSMC_34 TSMC_67 TSMC_68 TSMC_41 TSMC_83 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_Y_M4_SB 
XIDEC_Y[3] TSMC_9 TSMC_10 TSMC_35 TSMC_67 TSMC_68 TSMC_41 TSMC_84 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_Y_M4_SB 
XIDEC_Y[4] TSMC_9 TSMC_11 TSMC_36 TSMC_67 TSMC_68 TSMC_41 TSMC_85 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_Y_M4_SB 
XIDEC_Y[5] TSMC_9 TSMC_11 TSMC_37 TSMC_67 TSMC_68 TSMC_41 TSMC_86 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_Y_M4_SB 
XIDEC_Y[6] TSMC_9 TSMC_11 TSMC_38 TSMC_67 TSMC_68 TSMC_41 TSMC_87 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_Y_M4_SB 
XIDEC_Y[7] TSMC_9 TSMC_11 TSMC_39 TSMC_67 TSMC_68 TSMC_41 TSMC_88 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_Y_M4_SB 
XIDEC_CKD TSMC_9 TSMC_10 TSMC_6 TSMC_7 TSMC_67 TSMC_68 TSMC_47 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_DCLK_M4_SB_V2 
XIDEC_X1[0] TSMC_9 TSMC_10 TSMC_20 TSMC_67 TSMC_68 TSMC_41 TSMC_94 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_WLNAD2_SB_X1 
XIDEC_X1[1] TSMC_9 TSMC_10 TSMC_21 TSMC_67 TSMC_68 TSMC_41 TSMC_95 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_WLNAD2_SB_X1 
XIDEC_X1[2] TSMC_9 TSMC_10 TSMC_22 TSMC_67 TSMC_68 TSMC_41 TSMC_96 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_WLNAD2_SB_X1 
XIDEC_X1[3] TSMC_9 TSMC_10 TSMC_23 TSMC_67 TSMC_68 TSMC_41 TSMC_97 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_WLNAD2_SB_X1 
XIDEC_X1[4] TSMC_9 TSMC_10 TSMC_24 TSMC_67 TSMC_68 TSMC_41 TSMC_99 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_WLNAD2_SB_X1 
XIDEC_X1[5] TSMC_9 TSMC_10 TSMC_25 TSMC_67 TSMC_68 TSMC_41 TSMC_100 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_WLNAD2_SB_X1 
XIDEC_X1[6] TSMC_9 TSMC_10 TSMC_26 TSMC_67 TSMC_68 TSMC_41 TSMC_101 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_WLNAD2_SB_X1 
XIDEC_X1[7] TSMC_9 TSMC_10 TSMC_27 TSMC_67 TSMC_68 TSMC_41 TSMC_102 VDDMHD VDDM 
+ TSMC_44 S1CSLVTSW400W90_DECB1_WLNAD2_SB_X1 
XCEBBUF TSMC_3 TSMC_4 TSMC_5 TSMC_40 TSMC_68 TSMC_62 TSMC_67 TSMC_43 VDDMHD 
+ VDDM TSMC_44 S1CSLVTSW400W90_ENBUFB_BASE 
XI381[0] TSMC_109 TSMC_110 TSMC_111 TSMC_63 TSMC_64 VDDMHD VDDM TSMC_44 
+ S1CSLVTSW400W90_DECB2_SB 
XI381[1] TSMC_109 TSMC_110 TSMC_112 TSMC_65 TSMC_66 VDDMHD VDDM TSMC_44 
+ S1CSLVTSW400W90_DECB2_SB 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    RESETD_884_M4_SB_NBL
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_RESETD_884_M4_SB_NBL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 VDDHD TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 
*.PININFO  TSMC_2:I TSMC_3:I TSMC_6:I TSMC_9:I TSMC_10:I TSMC_14:I TSMC_16:I 
*.PININFO  TSMC_17:I 
*.PININFO  TSMC_18:I TSMC_19:I TSMC_20:I TSMC_1:O TSMC_4:O TSMC_5:O TSMC_7:O 
*.PININFO  TSMC_8:O TSMC_15:O TSMC_11:B VDDHD:B TSMC_12:B TSMC_13:B 
XTSEL_READ TSMC_3 TSMC_16 TSMC_17 VDDHD TSMC_12 TSMC_13 TSMC_21 TSMC_22 
+ S1CSLVTSW400W90_RESETD_TSEL 
MM10 TSMC_23 TSMC_9 TSMC_11 TSMC_12 pch_lvt_mac l=16.0n nfin=3 m=1 
MP0 TSMC_11 TSMC_1 TSMC_12 TSMC_12 pch_lvt_mac l=20n nfin=4 m=3 
MM0 TSMC_24 TSMC_25 VDDHD TSMC_12 pch_lvt_mac l=20n nfin=5 m=1 
MI537 TSMC_1 TSMC_25 VDDHD TSMC_12 pch_svt_mac l=16.0n nfin=8 m=4 
MM5 TSMC_23 TSMC_26 TSMC_27 TSMC_12 pch_lvt_mac l=20n nfin=3 m=1 
MM12 TSMC_23 TSMC_26 TSMC_11 TSMC_13 nch_lvt_mac l=16.0n nfin=4 m=2 
MM11 TSMC_1 TSMC_25 TSMC_13 TSMC_13 nch_lvt_mac l=16.0n nfin=5 m=4 
MM4 TSMC_23 TSMC_9 TSMC_27 TSMC_13 nch_lvt_mac l=20n nfin=4 m=2 
MM1 TSMC_8 TSMC_25 TSMC_13 TSMC_13 nch_lvt_mac l=20n nfin=5 m=1 
XTSEL_WT TSMC_28 TSMC_29 VDDHD TSMC_12 TSMC_13 TSMC_18 TSMC_19 
+ S1CSLVTSW400W90_RESETD_WTSEL_SB_NEW 
XNAND3 TSMC_22 TSMC_21 TSMC_3 TSMC_13 TSMC_13 TSMC_12 TSMC_12 TSMC_25 
+ S1CSLVTSW400W90_nand3_lvt_mac_pcell_2 n_totalM=2 n_nfin=9 n_l=16.0n 
+ p_totalM=2 p_nfin=3 p_l=16.0n 
XI667 TSMC_28 TSMC_2 TSMC_30 TSMC_13 TSMC_13 VDDHD TSMC_12 TSMC_31 
+ S1CSLVTSW400W90_nand3_lvt_mac_pcell_2 n_totalM=1 n_nfin=9 n_l=16.0n 
+ p_totalM=1 p_nfin=3 p_l=16.0n 
XI696 TSMC_28 TSMC_29 TSMC_13 TSMC_13 VDDHD TSMC_12 TSMC_32 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI658 TSMC_20 TSMC_1 TSMC_13 TSMC_13 VDDHD TSMC_12 TSMC_33 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI728 TSMC_1 TSMC_34 TSMC_13 TSMC_13 VDDHD TSMC_12 TSMC_27 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI666 TSMC_31 TSMC_35 TSMC_13 TSMC_13 VDDHD TSMC_12 TSMC_36 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=16.0n 
+ p_totalM=1 p_nfin=3 p_l=16.0n 
XI654 TSMC_33 TSMC_32 TSMC_13 TSMC_13 TSMC_24 TSMC_12 TSMC_8 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=5 n_l=20n p_totalM=1 
+ p_nfin=5 p_l=20n 
XI725 TSMC_13 TSMC_13 TSMC_9 TSMC_26 VDDHD TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI730 TSMC_13 TSMC_13 TSMC_37 TSMC_38 VDDHD TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI731 TSMC_13 TSMC_13 TSMC_38 TSMC_39 VDDHD TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI732 TSMC_13 TSMC_13 TSMC_39 TSMC_40 VDDHD TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI733 TSMC_13 TSMC_13 TSMC_40 TSMC_30 VDDHD TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI703 TSMC_13 TSMC_13 TSMC_14 TSMC_37 VDDHD TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI695 TSMC_13 TSMC_13 TSMC_41 TSMC_4 VDDHD TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=3 n_nfin=6 n_l=20n p_totalM=4 
+ p_nfin=7 p_l=20n 
XI679 TSMC_13 TSMC_13 TSMC_36 TSMC_42 TSMC_12 TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=9 n_l=16.0n p_totalM=1 
+ p_nfin=8 p_l=16.0n 
XI693 TSMC_13 TSMC_13 TSMC_3 TSMC_41 VDDHD TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=2 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=4 p_l=20n 
XI713 TSMC_13 TSMC_13 TSMC_23 TSMC_28 VDDHD TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=16.0n p_totalM=2 
+ p_nfin=3 p_l=16.0n 
XI718 TSMC_13 TSMC_13 TSMC_6 TSMC_34 VDDHD TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=5 p_l=20n 
XI533 TSMC_13 TSMC_13 TSMC_25 TSMC_43 VDDHD TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI686 TSMC_13 TSMC_13 TSMC_44 TSMC_35 VDDHD TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI687 TSMC_13 TSMC_13 TSMC_42 TSMC_15 VDDHD TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=8 n_nfin=7 n_l=16.0n p_totalM=8 
+ p_nfin=10 p_l=16.0n 
XI534 TSMC_13 TSMC_13 TSMC_43 TSMC_45 TSMC_12 TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI535 TSMC_13 TSMC_13 TSMC_45 TSMC_46 VDDHD TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI536 TSMC_13 TSMC_13 TSMC_46 TSMC_47 TSMC_12 TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI685 TSMC_13 TSMC_13 TSMC_33 TSMC_44 VDDHD TSMC_12 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    CKG_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_CKG_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDDHD TSMC_6 
+ TSMC_7 
*.PININFO  TSMC_2:I TSMC_3:I TSMC_5:I TSMC_1:O TSMC_4:O VDDHD:B TSMC_6:B 
*.PININFO  TSMC_7:B 
XI58 TSMC_7 TSMC_7 TSMC_8 TSMC_4 VDDHD TSMC_6 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=2 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
MM0 TSMC_1 TSMC_9 VDDHD TSMC_6 pch_lvt_mac l=16.0n nfin=4 m=1 
MM26 TSMC_1 TSMC_10 VDDHD TSMC_6 pch_lvt_mac l=16.0n nfin=4 m=4 
MM1 TSMC_11 TSMC_10 TSMC_7 TSMC_7 nch_lvt_mac l=16.0n nfin=8 m=3 
MM34 TSMC_1 TSMC_9 TSMC_11 TSMC_7 nch_lvt_mac l=16.0n nfin=8 m=3 
XNAND2 TSMC_2 TSMC_8 TSMC_7 TSMC_7 VDDHD TSMC_6 TSMC_12 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XNAND5 TSMC_4 TSMC_1 TSMC_7 TSMC_7 TSMC_6 TSMC_6 TSMC_9 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XNAND0 TSMC_1 TSMC_5 TSMC_7 TSMC_7 VDDHD TSMC_6 TSMC_13 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XNAND3 TSMC_12 TSMC_13 TSMC_7 TSMC_7 VDDHD TSMC_6 TSMC_8 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XNAND12 TSMC_2 TSMC_3 TSMC_4 TSMC_7 TSMC_7 TSMC_6 TSMC_6 TSMC_10 
+ S1CSLVTSW400W90_nand3_lvt_mac_pcell_2 n_totalM=1 n_nfin=10 n_l=16.0n 
+ p_totalM=1 p_nfin=4 p_l=16.0n 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    COTH_M4_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_COTH_M4_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 VDDM VDDMHD 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
*.PININFO  TSMC_3:I TSMC_4:I TSMC_7:I TSMC_8:I TSMC_10:I TSMC_11:I TSMC_12:I 
*.PININFO  TSMC_13:I TSMC_16:I 
*.PININFO  TSMC_21:I TSMC_22:I TSMC_23:I TSMC_1:O TSMC_5:O TSMC_6:O TSMC_9:O 
*.PININFO  TSMC_17:O TSMC_18:O TSMC_19:O TSMC_20:O TSMC_2:B TSMC_14:B VDDM:B 
*.PININFO  VDDMHD:B TSMC_15:B 
XRESETD TSMC_1 TSMC_2 TSMC_5 TSMC_6 TSMC_24 TSMC_7 TSMC_20 TSMC_25 TSMC_12 
+ TSMC_13 TSMC_14 VDDMHD VDDM TSMC_15 TSMC_18 TSMC_19 TSMC_10 TSMC_11 
+ TSMC_21 TSMC_22 TSMC_23 S1CSLVTSW400W90_RESETD_884_M4_SB_NBL 
XWEBBUF TSMC_3 TSMC_4 VDDMHD VDDM TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ S1CSLVTSW400W90_WEBBUF_SB_BASE 
XCKG TSMC_5 TSMC_7 TSMC_8 TSMC_9 TSMC_25 VDDMHD VDDM TSMC_15 
+ S1CSLVTSW400W90_CKG_SB 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    CNT_M4_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_CNT_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 VDD TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 
*.PININFO  TSMC_4:I TSMC_8:I TSMC_9:I TSMC_42:I TSMC_43:I TSMC_45:I TSMC_48:I 
*.PININFO  TSMC_50:I 
*.PININFO  TSMC_51:I TSMC_52:I TSMC_53:I TSMC_54:I TSMC_55:I TSMC_56:I 
*.PININFO  TSMC_57:I 
*.PININFO  TSMC_58:I TSMC_59:I TSMC_60:I TSMC_61:I TSMC_62:I TSMC_63:I 
*.PININFO  TSMC_64:I TSMC_1:O 
*.PININFO  TSMC_2:O TSMC_3:O TSMC_5:O TSMC_6:O TSMC_7:O TSMC_10:O TSMC_11:O 
*.PININFO  TSMC_12:O TSMC_13:O TSMC_14:O TSMC_15:O TSMC_16:O 
*.PININFO  TSMC_17:O TSMC_18:O TSMC_19:O TSMC_20:O TSMC_21:O 
*.PININFO  TSMC_22:O TSMC_23:O TSMC_24:O TSMC_25:O TSMC_26:O 
*.PININFO  TSMC_27:O TSMC_28:O TSMC_29:O TSMC_30:O TSMC_31:O 
*.PININFO  TSMC_32:O TSMC_33:O TSMC_34:O TSMC_35:O TSMC_36:O 
*.PININFO  TSMC_37:O TSMC_38:O TSMC_39:O TSMC_40:O TSMC_41:O TSMC_44:O 
*.PININFO  TSMC_49:O TSMC_46:B VDD:B TSMC_47:B 
Xcdec TSMC_1 TSMC_2 TSMC_4 TSMC_65 TSMC_66 TSMC_5 TSMC_6 TSMC_7 TSMC_67 TSMC_9 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_34 TSMC_35 
+ TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 VDD VDD TSMC_47 TSMC_72 TSMC_73 TSMC_49 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_74 TSMC_75 S1CSLVTSW400W90_CDEC_M4_SB_BASE 
XCOTHERS TSMC_3 TSMC_3 TSMC_65 TSMC_66 TSMC_7 TSMC_67 TSMC_9 TSMC_68 TSMC_71 
+ TSMC_42 TSMC_43 TSMC_45 TSMC_76 TSMC_46 VDD VDD TSMC_47 TSMC_48 
+ TSMC_73 TSMC_49 TSMC_44 TSMC_77 TSMC_50 TSMC_51 TSMC_52 
+ S1CSLVTSW400W90_COTH_M4_BASE 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    DIN_M4_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_DIN_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDDHD TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_7:O TSMC_8:O TSMC_4:B VDDHD:B 
*.PININFO  TSMC_5:B TSMC_6:B 
MMNCKGW TSMC_9 TSMC_10 TSMC_6 TSMC_6 nch_lvt_mac l=20n nfin=4 m=1 
MMNLCHDXCLK TSMC_11 TSMC_12 TSMC_13 TSMC_6 nch_lvt_mac l=20n nfin=2 m=1 
MM35 TSMC_14 TSMC_15 TSMC_6 TSMC_6 nch_lvt_mac l=20n nfin=2 m=2 
MMNLCHBXIN TSMC_16 TSMC_15 TSMC_6 TSMC_6 nch_lvt_mac l=20n nfin=2 m=1 
MMNGW TSMC_9 TSMC_17 TSMC_6 TSMC_6 nch_lvt_mac l=20n nfin=4 m=1 
MMNLCHBWIN TSMC_18 TSMC_1 TSMC_19 TSMC_6 nch_lvt_mac l=20n nfin=2 m=1 
MMNLCHDCLK TSMC_6 TSMC_10 TSMC_20 TSMC_6 nch_lvt_mac l=20n nfin=2 m=1 
MMNLCHBXCLK TSMC_18 TSMC_12 TSMC_16 TSMC_6 nch_lvt_mac l=20n nfin=2 m=1 
MMNLCHDXIN TSMC_6 TSMC_21 TSMC_13 TSMC_6 nch_lvt_mac l=20n nfin=2 m=1 
MMNCKGWB TSMC_22 TSMC_10 TSMC_6 TSMC_6 nch_lvt_mac l=20n nfin=4 m=1 
MMNLCHBWCLK TSMC_19 TSMC_10 TSMC_6 TSMC_6 nch_lvt_mac l=20n nfin=2 m=1 
MMNLCHDIN TSMC_11 TSMC_3 TSMC_20 TSMC_6 nch_lvt_mac l=20n nfin=2 m=1 
MMNGWB TSMC_22 TSMC_23 TSMC_6 TSMC_6 nch_lvt_mac l=20n nfin=4 m=1 
MMPLCHBWCLK TSMC_24 TSMC_12 VDDHD TSMC_5 pch_lvt_mac l=20n nfin=2 m=1 
MMPLCHDCLK VDDHD TSMC_12 TSMC_25 TSMC_5 pch_lvt_mac l=20n nfin=2 m=1 
MMPCKGW TSMC_26 TSMC_10 VDDHD TSMC_5 pch_lvt_mac l=20n nfin=6 m=2 
MMPLCHDXIN VDDHD TSMC_21 TSMC_27 TSMC_5 pch_lvt_mac l=20n nfin=2 m=1 
MM33 TSMC_23 TSMC_15 VDDHD TSMC_5 pch_lvt_mac l=20n nfin=2 m=1 
MM36 TSMC_17 TSMC_15 VDDHD TSMC_5 pch_lvt_mac l=20n nfin=2 m=1 
MMPLCHDXCLK TSMC_11 TSMC_10 TSMC_27 TSMC_5 pch_lvt_mac l=20n nfin=2 m=1 
MMPGWB TSMC_22 TSMC_23 TSMC_26 TSMC_5 pch_lvt_mac l=20n nfin=6 m=1 
MMPLCHDIN TSMC_11 TSMC_3 TSMC_25 TSMC_5 pch_lvt_mac l=20n nfin=2 m=1 
MMPGW TSMC_9 TSMC_17 TSMC_26 TSMC_5 pch_lvt_mac l=20n nfin=6 m=1 
MMPLCHBXCLK TSMC_18 TSMC_10 TSMC_28 TSMC_5 pch_lvt_mac l=20n nfin=2 m=1 
MMPLCHBWIN TSMC_18 TSMC_1 TSMC_24 TSMC_5 pch_lvt_mac l=20n nfin=2 m=1 
MMPLCHBXIN TSMC_28 TSMC_15 VDDHD TSMC_5 pch_lvt_mac l=20n nfin=2 m=1 
XI395 TSMC_14 TSMC_6 TSMC_11 TSMC_23 VDDHD TSMC_5 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XIWT TSMC_4 TSMC_6 TSMC_9 TSMC_8 VDDHD TSMC_5 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=3 n_nfin=9 n_l=20n p_totalM=3 
+ p_nfin=2 p_l=20n 
XICKD1D TSMC_6 TSMC_6 TSMC_2 TSMC_10 VDDHD TSMC_5 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI396 TSMC_14 TSMC_6 TSMC_21 TSMC_17 VDDHD TSMC_5 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XIBXL1B TSMC_6 TSMC_6 TSMC_18 TSMC_15 VDDHD TSMC_5 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XIWC TSMC_4 TSMC_6 TSMC_22 TSMC_7 VDDHD TSMC_5 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=3 n_nfin=9 n_l=20n p_totalM=3 
+ p_nfin=2 p_l=20n 
XICKD2 TSMC_6 TSMC_6 TSMC_10 TSMC_12 VDDHD TSMC_5 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XIDXL1B TSMC_6 TSMC_6 TSMC_11 TSMC_21 VDDHD TSMC_5 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    YPASS_M4_SB_NBL_V2
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_YPASS_M4_SB_NBL_V2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 
*.PININFO  TSMC_9:I TSMC_18:I TSMC_19:I TSMC_20:I TSMC_21:I TSMC_22:I TSMC_23:I 
*.PININFO  TSMC_24:I 
*.PININFO  TSMC_25:I TSMC_10:O TSMC_1:B TSMC_2:B TSMC_3:B TSMC_4:B TSMC_5:B 
*.PININFO  TSMC_6:B 
*.PININFO  TSMC_7:B TSMC_8:B TSMC_11:B TSMC_12:B TSMC_13:B TSMC_14:B TSMC_15:B 
*.PININFO  TSMC_16:B TSMC_17:B 
XIWCS[4] TSMC_13 TSMC_15 TSMC_22 TSMC_26 TSMC_14 TSMC_14 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XIWCS[5] TSMC_13 TSMC_15 TSMC_23 TSMC_27 TSMC_14 TSMC_14 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XIWCS[6] TSMC_13 TSMC_15 TSMC_24 TSMC_28 TSMC_14 TSMC_14 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XIWCS[7] TSMC_13 TSMC_15 TSMC_25 TSMC_29 TSMC_14 TSMC_14 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
MMNWCS_BLB[0] TSMC_5 TSMC_26 TSMC_16 TSMC_15 nch_ulvt_mac l=20n nfin=5 
+ m=2 
MMNWCS_BLB[1] TSMC_6 TSMC_27 TSMC_16 TSMC_15 nch_ulvt_mac l=20n nfin=5 
+ m=2 
MMNWCS_BLB[2] TSMC_7 TSMC_28 TSMC_16 TSMC_15 nch_ulvt_mac l=20n nfin=5 
+ m=2 
MMNWCS_BLB[3] TSMC_8 TSMC_29 TSMC_16 TSMC_15 nch_ulvt_mac l=20n nfin=5 
+ m=2 
MMNWCS_BL[0] TSMC_1 TSMC_26 TSMC_17 TSMC_15 nch_ulvt_mac l=20n nfin=5 
+ m=2 
MMNWCS_BL[1] TSMC_2 TSMC_27 TSMC_17 TSMC_15 nch_ulvt_mac l=20n nfin=5 
+ m=2 
MMNWCS_BL[2] TSMC_3 TSMC_28 TSMC_17 TSMC_15 nch_ulvt_mac l=20n nfin=5 
+ m=2 
MMNWCS_BL[3] TSMC_4 TSMC_29 TSMC_17 TSMC_15 nch_ulvt_mac l=20n nfin=5 
+ m=2 
MMNBLEQB TSMC_10 TSMC_9 TSMC_15 TSMC_15 nch_lvt_mac l=20n nfin=4 m=1 
MMNBLEQT TSMC_30 TSMC_10 TSMC_15 TSMC_15 nch_lvt_mac l=20n nfin=2 m=2 
MMPBLEQB TSMC_10 TSMC_9 TSMC_14 TSMC_14 pch_lvt_mac l=20n nfin=4 m=1 
MMPRCS_BLB[0] TSMC_12 TSMC_18 TSMC_5 TSMC_14 pch_lvt_mac l=20n nfin=3 
+ m=1 
MMPRCS_BLB[1] TSMC_12 TSMC_19 TSMC_6 TSMC_14 pch_lvt_mac l=20n nfin=3 
+ m=1 
MMPRCS_BLB[2] TSMC_12 TSMC_20 TSMC_7 TSMC_14 pch_lvt_mac l=20n nfin=3 
+ m=1 
MMPRCS_BLB[3] TSMC_12 TSMC_21 TSMC_8 TSMC_14 pch_lvt_mac l=20n nfin=3 
+ m=1 
MMPDLBPRE TSMC_12 TSMC_30 TSMC_14 TSMC_14 pch_lvt_mac l=20n nfin=2 m=2 
MMPDLPRE TSMC_14 TSMC_30 TSMC_11 TSMC_14 pch_lvt_mac l=20n nfin=2 m=2 
MMPRCS_BL[0] TSMC_11 TSMC_18 TSMC_1 TSMC_14 pch_lvt_mac l=20n nfin=3 
+ m=1 
MMPRCS_BL[1] TSMC_11 TSMC_19 TSMC_2 TSMC_14 pch_lvt_mac l=20n nfin=3 
+ m=1 
MMPRCS_BL[2] TSMC_11 TSMC_20 TSMC_3 TSMC_14 pch_lvt_mac l=20n nfin=3 
+ m=1 
MMPRCS_BL[3] TSMC_11 TSMC_21 TSMC_4 TSMC_14 pch_lvt_mac l=20n nfin=3 
+ m=1 
MMPBLEQT TSMC_30 TSMC_10 TSMC_14 TSMC_14 pch_lvt_mac l=20n nfin=5 m=2 
MMPXBL[0] TSMC_1 TSMC_5 TSMC_14 TSMC_14 pch_lvt_mac l=20n nfin=3 m=1 
MMPXBL[1] TSMC_2 TSMC_6 TSMC_14 TSMC_14 pch_lvt_mac l=20n nfin=3 m=1 
MMPXBL[2] TSMC_3 TSMC_7 TSMC_14 TSMC_14 pch_lvt_mac l=20n nfin=3 m=1 
MMPXBL[3] TSMC_4 TSMC_8 TSMC_14 TSMC_14 pch_lvt_mac l=20n nfin=3 m=1 
MMPXBLB[0] TSMC_5 TSMC_1 TSMC_14 TSMC_14 pch_lvt_mac l=20n nfin=3 m=1 
MMPXBLB[1] TSMC_6 TSMC_2 TSMC_14 TSMC_14 pch_lvt_mac l=20n nfin=3 m=1 
MMPXBLB[2] TSMC_7 TSMC_3 TSMC_14 TSMC_14 pch_lvt_mac l=20n nfin=3 m=1 
MMPXBLB[3] TSMC_8 TSMC_4 TSMC_14 TSMC_14 pch_lvt_mac l=20n nfin=3 m=1 
XPRECHARGE[0] TSMC_1 TSMC_5 TSMC_30 TSMC_14 TSMC_14 
+ S1CSLVTSW400W90_PRECHARGE_SB_SD 
XPRECHARGE[1] TSMC_2 TSMC_6 TSMC_30 TSMC_14 TSMC_14 
+ S1CSLVTSW400W90_PRECHARGE_SB_SD 
XPRECHARGE[2] TSMC_3 TSMC_7 TSMC_30 TSMC_14 TSMC_14 
+ S1CSLVTSW400W90_PRECHARGE_SB_SD 
XPRECHARGE[3] TSMC_4 TSMC_8 TSMC_30 TSMC_14 TSMC_14 
+ S1CSLVTSW400W90_PRECHARGE_SB_SD 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    DOUT_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_DOUT_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDDHD TSMC_6 
+ TSMC_7 
*.PININFO  TSMC_1:I TSMC_5:I TSMC_4:O TSMC_2:B TSMC_3:B VDDHD:B TSMC_6:B 
*.PININFO  TSMC_7:B 
MMPSA[0] TSMC_8 TSMC_9 VDDHD TSMC_6 pch_lvt_mac l=20n nfin=5 m=1 
MMPSAEQ TSMC_8 TSMC_10 TSMC_9 TSMC_6 pch_lvt_mac l=20n nfin=5 m=2 
MMPLCHQBCLK TSMC_11 TSMC_12 TSMC_13 TSMC_6 pch_lvt_mac l=20n nfin=3 m=1 
MMPSAPRE[1] TSMC_9 TSMC_10 VDDHD TSMC_6 pch_lvt_mac l=20n nfin=5 m=1 
MMPLCHSAIN[1] TSMC_14 TSMC_9 VDDHD TSMC_6 pch_lvt_mac l=16n nfin=6 m=1 
MMPSAPGB[0] TSMC_8 TSMC_15 TSMC_2 TSMC_6 pch_lvt_mac l=20n nfin=5 m=1 
MMPSAPGB[1] TSMC_9 TSMC_15 TSMC_3 TSMC_6 pch_lvt_mac l=20n nfin=5 m=1 
MMPLCHSACLK[0] TSMC_11 TSMC_16 TSMC_17 TSMC_6 pch_lvt_mac l=16n nfin=6 
+ m=1 
MMPSAPRE[0] TSMC_8 TSMC_10 VDDHD TSMC_6 pch_lvt_mac l=20n nfin=5 m=1 
MMPSA[1] TSMC_9 TSMC_8 VDDHD TSMC_6 pch_lvt_mac l=20n nfin=5 m=1 
MMPQ TSMC_4 TSMC_11 VDDHD TSMC_6 pch_lvt_mac l=20n nfin=4 m=4 
MMPLCHSACLK[1] TSMC_18 TSMC_16 TSMC_14 TSMC_6 pch_lvt_mac l=16n nfin=6 
+ m=1 
MMPLCHSAIN[0] TSMC_17 TSMC_8 VDDHD TSMC_6 pch_lvt_mac l=16n nfin=6 m=1 
MMPLCHQBIN TSMC_13 TSMC_19 VDDHD TSMC_6 pch_lvt_mac l=20n nfin=3 m=1 
MMNSA[0] TSMC_8 TSMC_9 TSMC_20 TSMC_7 nch_lvt_mac l=20n nfin=10 m=4 
MMNLCHSACLK[1] TSMC_18 TSMC_12 TSMC_21 TSMC_7 nch_lvt_mac l=16n nfin=3 
+ m=1 
MMNSAEN TSMC_20 TSMC_12 TSMC_7 TSMC_7 nch_lvt_mac l=20n nfin=10 m=4 
MMNSA[1] TSMC_9 TSMC_8 TSMC_20 TSMC_7 nch_lvt_mac l=20n nfin=10 m=4 
MMNLCHSAIN[1] TSMC_21 TSMC_9 TSMC_7 TSMC_7 nch_lvt_mac l=16n nfin=3 m=1 
MMNLCHSAIN[0] TSMC_22 TSMC_8 TSMC_7 TSMC_7 nch_lvt_mac l=16n nfin=3 m=1 
MMNLCHQBCLK TSMC_11 TSMC_16 TSMC_23 TSMC_7 nch_lvt_mac l=20n nfin=3 m=1 
MMNQ TSMC_4 TSMC_11 TSMC_7 TSMC_7 nch_lvt_mac l=20n nfin=4 m=4 
MMNLCHQBIN TSMC_23 TSMC_19 TSMC_7 TSMC_7 nch_lvt_mac l=20n nfin=3 m=1 
MMNLCHSACLK[0] TSMC_11 TSMC_12 TSMC_22 TSMC_7 nch_lvt_mac l=16n nfin=3 
+ m=1 
XIPGB TSMC_24 TSMC_16 TSMC_10 TSMC_7 TSMC_7 VDDHD TSMC_6 TSMC_15 
+ S1CSLVTSW400W90_nand3_lvt_mac_pcell_2 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI202 TSMC_1 TSMC_25 TSMC_7 TSMC_7 VDDHD TSMC_6 TSMC_26 
+ S1CSLVTSW400W90_nor2_lvt_mac_pcell_4 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XIPREB TSMC_16 TSMC_27 TSMC_7 TSMC_7 VDDHD TSMC_6 TSMC_10 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI185 TSMC_7 TSMC_7 TSMC_16 TSMC_28 VDDHD TSMC_6 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XIBLEQB TSMC_7 TSMC_7 TSMC_26 TSMC_27 VDDHD TSMC_6 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XISAEB TSMC_7 TSMC_7 TSMC_12 TSMC_16 VDDHD TSMC_6 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=2 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XISAE TSMC_7 TSMC_7 TSMC_29 TSMC_12 VDDHD TSMC_6 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=2 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XISAEC TSMC_7 TSMC_7 TSMC_5 TSMC_29 VDDHD TSMC_6 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI186 TSMC_7 TSMC_7 TSMC_28 TSMC_24 VDDHD TSMC_6 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI201 TSMC_7 TSMC_7 TSMC_1 TSMC_30 VDDHD TSMC_6 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI207 TSMC_7 TSMC_7 TSMC_30 TSMC_31 VDDHD TSMC_6 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XIQF TSMC_7 TSMC_7 TSMC_11 TSMC_19 VDDHD TSMC_6 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
XI209 TSMC_7 TSMC_7 TSMC_32 TSMC_25 VDDHD TSMC_6 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI208 TSMC_7 TSMC_7 TSMC_31 TSMC_32 VDDHD TSMC_6 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    MIO_M4_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_MIO_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ VDD TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
*.PININFO  TSMC_9:I TSMC_10:I TSMC_11:I TSMC_12:I TSMC_15:I TSMC_17:I TSMC_18:I 
*.PININFO  TSMC_19:I TSMC_20:I 
*.PININFO  TSMC_21:I TSMC_22:I TSMC_23:I TSMC_24:I TSMC_14:O TSMC_1:B TSMC_2:B 
*.PININFO  TSMC_3:B TSMC_4:B 
*.PININFO  TSMC_5:B TSMC_6:B TSMC_7:B TSMC_8:B TSMC_13:B VDD:B TSMC_16:B 
XDIN TSMC_10 TSMC_11 TSMC_12 TSMC_13 VDD VDD TSMC_16 TSMC_25 TSMC_26 
+ S1CSLVTSW400W90_DIN_M4_SB_BASE 
XYPASS TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_27 
+ TSMC_28 TSMC_29 TSMC_13 VDD TSMC_16 TSMC_25 TSMC_26 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ S1CSLVTSW400W90_YPASS_M4_SB_NBL_V2 
XDOUT TSMC_27 TSMC_28 TSMC_29 TSMC_14 TSMC_15 VDD VDD TSMC_16 
+ S1CSLVTSW400W90_DOUT_SB 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    XDRV_STRAP_BT_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_XDRV_STRAP_BT_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 
*.PININFO  TSMC_1:B TSMC_2:B TSMC_3:B TSMC_4:B 
MM0 TSMC_2 TSMC_1 TSMC_4 TSMC_4 nch_lvt_mac l=20n nfin=12 m=4 
MM10 TSMC_2 TSMC_1 TSMC_4 TSMC_4 nch_lvt_mac l=20n nfin=6 m=12 
MM1 TSMC_2 TSMC_1 TSMC_3 TSMC_3 pch_lvt_mac l=20n nfin=3 m=10 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    MIO_M4_SB_BUF
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_MIO_M4_SB_BUF TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD TSMC_5 
*.PININFO  TSMC_1:I TSMC_3:I TSMC_2:O TSMC_4:O VDD:B TSMC_5:B 
XI8 TSMC_5 TSMC_5 TSMC_6 TSMC_7 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI9 TSMC_5 TSMC_5 TSMC_7 TSMC_4 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI15 TSMC_5 TSMC_5 TSMC_8 TSMC_2 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI14 TSMC_5 TSMC_5 TSMC_9 TSMC_8 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI16 TSMC_5 TSMC_5 TSMC_3 TSMC_6 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI17 TSMC_5 TSMC_5 TSMC_1 TSMC_9 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    DIO_TALL
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_DIO_TALL TSMC_1 VSS 
*.PININFO  TSMC_1:B VSS:B 
XDDIO_TALL VSS TSMC_1 ndio_mac nfin=2 l=2e-07 m=1 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    CNT_M4_SB_BUF
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_CNT_M4_SB_BUF TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 
*.PININFO  TSMC_1:I TSMC_3:I VDD:I TSMC_6:I TSMC_8:I TSMC_9:I TSMC_10:I 
*.PININFO  TSMC_11:I TSMC_12:I TSMC_13:I 
*.PININFO  TSMC_14:I TSMC_15:I TSMC_24:I TSMC_25:I TSMC_26:I TSMC_27:I TSMC_2:B 
*.PININFO  TSMC_4:B TSMC_5:B 
*.PININFO  TSMC_7:B TSMC_16:B TSMC_17:B TSMC_18:B TSMC_19:B TSMC_20:B TSMC_21:B 
*.PININFO  TSMC_22:B 
*.PININFO  TSMC_23:B TSMC_28:B TSMC_29:B TSMC_30:B TSMC_31:B 
XI32 TSMC_5 TSMC_5 TSMC_32 TSMC_4 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=2 n_nfin=10 n_l=20n p_totalM=2 
+ p_nfin=10 p_l=20n 
XI31 TSMC_5 TSMC_5 TSMC_3 TSMC_32 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=10 n_l=20n p_totalM=1 
+ p_nfin=10 p_l=20n 
XWEB_INV TSMC_5 TSMC_5 TSMC_6 TSMC_7 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI29[0] TSMC_5 TSMC_5 TSMC_24 TSMC_28 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI29[1] TSMC_5 TSMC_5 TSMC_25 TSMC_29 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI30 TSMC_5 TSMC_5 TSMC_1 TSMC_2 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=5 n_l=20n p_totalM=1 
+ p_nfin=7 p_l=20n 
XI28[0] TSMC_5 TSMC_5 TSMC_8 TSMC_16 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28[1] TSMC_5 TSMC_5 TSMC_9 TSMC_17 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28[2] TSMC_5 TSMC_5 TSMC_10 TSMC_18 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28[3] TSMC_5 TSMC_5 TSMC_11 TSMC_19 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28[4] TSMC_5 TSMC_5 TSMC_12 TSMC_20 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28[5] TSMC_5 TSMC_5 TSMC_13 TSMC_21 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28[6] TSMC_5 TSMC_5 TSMC_14 TSMC_22 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28[7] TSMC_5 TSMC_5 TSMC_15 TSMC_23 VDD VDD 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    DECB1_WAS
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_DECB1_WAS TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
*.PININFO  TSMC_1:I TSMC_6:I TSMC_4:O TSMC_2:B TSMC_3:B TSMC_5:B 
MMN0 TSMC_7 TSMC_1 TSMC_8 TSMC_5 nch_lvt_mac l=20n nfin=6 m=1 
MMN1 TSMC_8 TSMC_6 TSMC_5 TSMC_5 nch_lvt_mac l=20n nfin=6 m=1 
MMN2 TSMC_4 TSMC_7 TSMC_5 TSMC_5 nch_lvt_mac l=20n nfin=5 m=2 
MMP1 TSMC_7 TSMC_6 TSMC_3 TSMC_3 pch_lvt_mac l=20n nfin=3 m=1 
MMP2 TSMC_4 TSMC_7 TSMC_2 TSMC_3 pch_lvt_mac l=20n nfin=5 m=2 
MMP0 TSMC_7 TSMC_1 TSMC_3 TSMC_3 pch_lvt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    RESETD_TSEL_NBL
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_RESETD_TSEL_NBL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
*.PININFO  TSMC_1:I TSMC_4:I TSMC_5:I TSMC_7:O TSMC_8:O TSMC_2:B TSMC_3:B 
*.PININFO  TSMC_6:B 
CC2 TSMC_9 TSMC_6 600.0a $[CP] 
CC3 TSMC_10 TSMC_6 600.0a $[CP] 
CC0 TSMC_11 TSMC_6 600.0a $[CP] 
CC4 TSMC_12 TSMC_6 600.0a $[CP] 
MM16 TSMC_10 TSMC_1 TSMC_13 TSMC_6 nch_lvt_mac l=20n nfin=2 m=1 
MM10 TSMC_14 TSMC_9 TSMC_6 TSMC_6 nch_lvt_mac l=20n nfin=2 m=1 
MM9 TSMC_12 TSMC_9 TSMC_14 TSMC_6 nch_lvt_mac l=20n nfin=2 m=1 
MM3 TSMC_15 TSMC_10 TSMC_6 TSMC_6 nch_lvt_mac l=20n nfin=2 m=1 
MM2 TSMC_9 TSMC_10 TSMC_15 TSMC_6 nch_lvt_mac l=20n nfin=2 m=1 
MM22 TSMC_13 TSMC_1 TSMC_6 TSMC_6 nch_lvt_mac l=20n nfin=2 m=1 
MM6 TSMC_16 TSMC_9 TSMC_2 TSMC_3 pch_lvt_mac l=20n nfin=2 m=1 
MM1 TSMC_17 TSMC_10 TSMC_2 TSMC_3 pch_lvt_mac l=20n nfin=2 m=1 
MM31 TSMC_18 TSMC_1 TSMC_2 TSMC_3 pch_lvt_mac l=20n nfin=2 m=1 
MM7 TSMC_12 TSMC_9 TSMC_16 TSMC_3 pch_lvt_mac l=20n nfin=2 m=1 
MM30 TSMC_10 TSMC_1 TSMC_18 TSMC_3 pch_lvt_mac l=20n nfin=2 m=1 
MM0 TSMC_9 TSMC_10 TSMC_17 TSMC_3 pch_lvt_mac l=20n nfin=2 m=1 
XI92 TSMC_4 TSMC_11 TSMC_6 TSMC_6 TSMC_2 TSMC_3 TSMC_7 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI93 TSMC_8 TSMC_1 TSMC_6 TSMC_6 TSMC_2 TSMC_3 TSMC_11 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI91 TSMC_5 TSMC_12 TSMC_6 TSMC_6 TSMC_2 TSMC_3 TSMC_8 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    MIO_SB_EDGE
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_MIO_SB_EDGE TSMC_1 TSMC_2 TSMC_3 TSMC_4 
*.PININFO  TSMC_1:B TSMC_2:B TSMC_3:B TSMC_4:B 
MP0 TSMC_5 TSMC_5 TSMC_1 TSMC_1 pch_lvt_mac l=20n nfin=3 m=1 
MP2 TSMC_6 TSMC_7 TSMC_1 TSMC_1 pch_lvt_mac l=20n nfin=3 m=6 
MP7 TSMC_5 TSMC_7 TSMC_1 TSMC_1 pch_lvt_mac l=20n nfin=3 m=1 
MN3 TSMC_4 TSMC_5 TSMC_7 TSMC_4 nch_lvt_mac l=20n nfin=3 m=1 
MN1 TSMC_4 TSMC_5 TSMC_8 TSMC_4 nch_lvt_mac l=20n nfin=3 m=5 
MN0 TSMC_4 TSMC_7 TSMC_7 TSMC_4 nch_lvt_mac l=20n nfin=3 m=1 
XI18 TSMC_4 TSMC_4 TSMC_6 TSMC_3 TSMC_1 TSMC_1 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=8 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XI393 TSMC_4 TSMC_4 TSMC_8 TSMC_2 TSMC_1 TSMC_1 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=4 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    CNT_M4_SB_NBL
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_CNT_M4_SB_NBL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 VDDM VDDMHD TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 
*.PININFO  TSMC_1:I TSMC_7:I TSMC_8:I TSMC_9:I TSMC_10:I 
*.PININFO  TSMC_11:I TSMC_13:I TSMC_15:I TSMC_2:O TSMC_3:O 
*.PININFO  TSMC_4:O TSMC_5:O TSMC_6:O VDDM:B VDDMHD:B 
*.PININFO  TSMC_12:B TSMC_14:B 
XWASDEC TSMC_16 VDDMHD VDDM TSMC_17 TSMC_12 TSMC_13 
+ S1CSLVTSW400W90_DECB1_WAS 
MM9 TSMC_18 TSMC_19 TSMC_20 TSMC_12 nch_lvt_mac l=20n nfin=8 m=3 
MM1 TSMC_20 TSMC_19 TSMC_12 TSMC_12 nch_lvt_mac l=20n nfin=8 m=6 
MM5 TSMC_14 TSMC_19 TSMC_18 TSMC_12 nch_lvt_mac l=20n nfin=4 m=2 
MP0 TSMC_14 TSMC_19 VDDM VDDM pch_lvt_mac l=20n nfin=7 m=2 
XI750q TSMC_21 TSMC_22 TSMC_17 TSMC_12 TSMC_12 VDDM VDDM TSMC_23 
+ S1CSLVTSW400W90_nand3_lvt_mac_pcell_2 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI763 TSMC_12 TSMC_12 TSMC_14 TSMC_24 VDDMHD VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
XI753 TSMC_12 TSMC_12 TSMC_25 TSMC_19 VDDMHD VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=4 n_nfin=4 n_l=20n p_totalM=4 
+ p_nfin=4 p_l=20n 
XI3 TSMC_12 TSMC_12 TSMC_23 TSMC_26 VDDMHD VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=2 n_nfin=2 n_l=20n p_totalM=2 
+ p_nfin=2 p_l=20n 
XI764 TSMC_12 TSMC_12 TSMC_24 TSMC_27 VDDM VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=8 n_l=20n p_totalM=1 
+ p_nfin=8 p_l=20n 
XI765 TSMC_12 TSMC_12 TSMC_14 TSMC_28 VDDMHD VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
XI766 TSMC_12 TSMC_12 TSMC_28 TSMC_29 VDDM VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=8 n_l=20n p_totalM=1 
+ p_nfin=8 p_l=20n 
XI773 TSMC_12 TSMC_12 TSMC_30 TSMC_2 VDDM VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=6 n_nfin=8 n_l=20n p_totalM=6 
+ p_nfin=8 p_l=20n 
XI774 TSMC_12 TSMC_12 TSMC_29 TSMC_31 VDDMHD VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=6 n_nfin=4 n_l=20n p_totalM=6 
+ p_nfin=4 p_l=20n 
XI777 TSMC_12 TSMC_12 TSMC_27 TSMC_30 VDDMHD VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=6 n_nfin=4 n_l=20n p_totalM=6 
+ p_nfin=4 p_l=20n 
XI779 TSMC_12 TSMC_12 TSMC_31 TSMC_3 VDDM VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=6 n_nfin=8 n_l=20n p_totalM=6 
+ p_nfin=8 p_l=20n 
XI806 TSMC_12 TSMC_12 TSMC_32 TSMC_16 VDDMHD VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=2 n_nfin=2 n_l=20n p_totalM=2 
+ p_nfin=2 p_l=20n 
XI4 TSMC_12 TSMC_12 TSMC_26 TSMC_25 VDDM VDDM 
+ S1CSLVTSW400W90_inv_lvt_mac_pcell_0 n_totalM=2 n_nfin=2 n_l=20n p_totalM=2 
+ p_nfin=2 p_l=20n 
XI805 TSMC_1 TSMC_15 TSMC_12 TSMC_12 VDDM VDDM TSMC_32 
+ S1CSLVTSW400W90_nand2_lvt_mac_pcell_1 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XTSEL_WRITE TSMC_17 VDDMHD VDDM TSMC_10 TSMC_11 TSMC_12 TSMC_22 TSMC_21 
+ S1CSLVTSW400W90_RESETD_TSEL_NBL 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    XDRV_STRAP_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_XDRV_STRAP_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 
*.PININFO  TSMC_1:B TSMC_2:B TSMC_3:B TSMC_4:B 
MM10 TSMC_2 TSMC_1 TSMC_4 TSMC_4 nch_lvt_mac l=20n nfin=6 m=20 
MM1 TSMC_2 TSMC_1 TSMC_3 TSMC_3 pch_lvt_mac l=20n nfin=3 m=10 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    MCB_D0734_ONCELL
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_MCB_D0734_ONCELL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
*.PININFO  TSMC_1:B TSMC_2:B TSMC_3:B TSMC_4:B TSMC_5:B TSMC_6:B TSMC_7:B 
*.PININFO  TSMC_8:B 
Mpd11 TSMC_9 TSMC_5 TSMC_6 TSMC_6 nchpd_hdsr_mac l=20n nfin=1 m=1 
Mpd21 TSMC_10 TSMC_9 TSMC_6 TSMC_6 nchpd_hdsr_mac l=20n nfin=1 m=1 
Mpg21 TSMC_11 TSMC_7 TSMC_10 TSMC_6 nchpg_hdsr_mac l=20n nfin=1 m=1 
Mpd20 TSMC_12 TSMC_13 TSMC_6 TSMC_6 nchpd_hdsr_mac l=20n nfin=1 m=1 
Mpg11 TSMC_1 TSMC_2 TSMC_9 TSMC_6 nchpg_hdsr_mac l=20n nfin=1 m=1 
Mpg10 TSMC_1 TSMC_3 TSMC_13 TSMC_6 nchpg_hdsr_mac l=20n nfin=1 m=1 
Mpd10 TSMC_13 TSMC_5 TSMC_6 TSMC_6 nchpd_hdsr_mac l=20n nfin=1 m=1 
Mpg20 TSMC_11 TSMC_8 TSMC_12 TSMC_6 nchpg_hdsr_mac l=20n nfin=1 m=1 
Mpu11 TSMC_9 TSMC_5 TSMC_5 TSMC_4 pchpu_hdsr_mac l=20n nfin=1 m=1 
Mpu10 TSMC_13 TSMC_5 TSMC_5 TSMC_4 pchpu_hdsr_mac l=20n nfin=1 m=1 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    MCB_D0734_ONCELL_ISO
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_MCB_D0734_ONCELL_ISO TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 
*.PININFO  TSMC_1:B TSMC_2:B TSMC_3:B TSMC_4:B TSMC_5:B TSMC_6:B TSMC_7:B 
*.PININFO  TSMC_8:B 
*.PININFO  TSMC_9:B 
Mpg11 TSMC_1 TSMC_2 TSMC_10 TSMC_6 nchpg_hdsr_mac l=20n nfin=1 m=1 
Mpd11 TSMC_10 TSMC_5 TSMC_6 TSMC_6 nchpd_hdsr_mac l=20n nfin=1 m=1 
Mpd21 TSMC_11 TSMC_10 TSMC_6 TSMC_6 nchpd_hdsr_mac l=20n nfin=1 m=1 
Mpg21 TSMC_12 TSMC_8 TSMC_11 TSMC_6 nchpg_hdsr_mac l=20n nfin=1 m=1 
Mpd10 TSMC_13 TSMC_5 TSMC_6 TSMC_6 nchpd_hdsr_mac l=20n nfin=1 m=1 
Mpd20 TSMC_14 TSMC_13 TSMC_6 TSMC_6 nchpd_hdsr_mac l=20n nfin=1 m=1 
Mpg10 TSMC_1 TSMC_3 TSMC_13 TSMC_6 nchpg_hdsr_mac l=20n nfin=1 m=1 
Mpg20 TSMC_12 TSMC_7 TSMC_14 TSMC_6 nchpg_hdsr_mac l=20n nfin=1 m=1 
Mpu11 TSMC_10 TSMC_5 TSMC_5 TSMC_4 pchpu_hdsr_mac l=20n nfin=1 m=1 
Mpu10 TSMC_13 TSMC_5 TSMC_5 TSMC_4 pchpu_hdsr_mac l=20n nfin=1 m=1 
Mpu20 TSMC_15 TSMC_13 TSMC_9 TSMC_4 pchpu_hdsr_mac l=20n nfin=1 m=1 
.ENDS

************************************************************************
* Library Name: N16_HDSPSB_LEAFCELL
* Cell Name:    MCB_D0734_OFFCELL
* View Name:    schematic
************************************************************************

.SUBCKT S1CSLVTSW400W90_MCB_D0734_OFFCELL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
*.PININFO  TSMC_1:B TSMC_2:B TSMC_3:B TSMC_4:B TSMC_5:B TSMC_6:B TSMC_7:B 
*.PININFO  TSMC_8:B 
Mpu11 TSMC_9 TSMC_10 TSMC_3 TSMC_2 pchpu_hdsr_mac l=20n nfin=1 m=1 
Mpu21 TSMC_10 TSMC_9 TSMC_8 TSMC_2 pchpu_hdsr_mac l=20n nfin=1 m=1 
Mpu10 TSMC_11 TSMC_12 TSMC_3 TSMC_2 pchpu_hdsr_mac l=20n nfin=1 m=1 
Mpu20 TSMC_12 TSMC_11 TSMC_7 TSMC_2 pchpu_hdsr_mac l=20n nfin=1 m=1 
Mpg21 TSMC_13 TSMC_5 TSMC_10 TSMC_4 nchpg_hdsr_mac l=20n nfin=1 m=1 
Mpd11 TSMC_9 TSMC_10 TSMC_14 TSMC_4 nchpd_hdsr_mac l=20n nfin=1 m=1 
Mpd21 TSMC_10 TSMC_9 TSMC_4 TSMC_4 nchpd_hdsr_mac l=20n nfin=1 m=1 
Mpd20 TSMC_12 TSMC_11 TSMC_4 TSMC_4 nchpd_hdsr_mac l=20n nfin=1 m=1 
Mpg11 TSMC_1 TSMC_4 TSMC_9 TSMC_4 nchpg_hdsr_mac l=20n nfin=1 m=1 
Mpg20 TSMC_13 TSMC_6 TSMC_12 TSMC_4 nchpg_hdsr_mac l=20n nfin=1 m=1 
Mpg10 TSMC_1 TSMC_4 TSMC_11 TSMC_4 nchpg_hdsr_mac l=20n nfin=1 m=1 
Mpd10 TSMC_11 TSMC_12 TSMC_14 TSMC_4 nchpd_hdsr_mac l=20n nfin=1 m=1 
.ENDS




**** End of leaf cells

.SUBCKT S1CSLVTSW400W90_MCB_ARR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDDAI TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 
+ TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 
+ TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 
+ TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 
+ TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 
XMCB_0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_11 TSMC_12 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_13 TSMC_14 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_15 TSMC_16 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_3 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_17 TSMC_18 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_19 TSMC_20 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_5 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_21 TSMC_22 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_6 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_23 TSMC_24 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_7 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_25 TSMC_26 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_27 TSMC_28 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_9 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_29 TSMC_30 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_10 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_31 TSMC_32 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_11 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_33 TSMC_34 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_12 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_35 TSMC_36 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_13 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_37 TSMC_38 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_14 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_39 TSMC_40 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_15 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_41 TSMC_42 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_16 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_43 TSMC_44 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_17 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_45 TSMC_46 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_18 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_47 TSMC_48 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_19 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_49 TSMC_50 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_20 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_51 TSMC_52 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_21 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_53 TSMC_54 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_22 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_55 TSMC_56 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_23 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_57 TSMC_58 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_24 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_59 TSMC_60 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_25 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_61 TSMC_62 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_26 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_63 TSMC_64 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_27 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_65 TSMC_66 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_28 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_67 TSMC_68 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_29 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_69 TSMC_70 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_30 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_71 TSMC_72 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_31 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_73 TSMC_74 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_32 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_75 TSMC_76 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_33 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_77 TSMC_78 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_34 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_79 TSMC_80 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_35 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_81 TSMC_82 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_36 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_83 TSMC_84 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_37 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_85 TSMC_86 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_38 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_87 TSMC_88 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_39 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_89 TSMC_90 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_40 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_91 TSMC_92 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_41 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_93 TSMC_94 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_42 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_95 TSMC_96 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_43 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_97 TSMC_98 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_44 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_99 TSMC_100 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_45 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_101 TSMC_102 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_46 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_103 TSMC_104 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_47 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_105 TSMC_106 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_48 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_107 TSMC_108 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_49 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_109 TSMC_110 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_50 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_111 TSMC_112 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_51 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_113 TSMC_114 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_52 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_115 TSMC_116 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_53 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_117 TSMC_118 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_54 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_119 TSMC_120 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_55 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_121 TSMC_122 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_56 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_123 TSMC_124 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_57 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_125 TSMC_126 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_58 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_127 TSMC_128 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_59 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_129 TSMC_130 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_60 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_131 TSMC_132 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_61 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_133 TSMC_134 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_62 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_135 TSMC_136 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_63 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_137 TSMC_138 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_64 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_139 TSMC_140 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_65 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_141 TSMC_142 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_66 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_143 TSMC_144 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_67 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_145 TSMC_146 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_68 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_147 TSMC_148 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_69 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_149 TSMC_150 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_70 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_151 TSMC_152 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_71 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_153 TSMC_154 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_72 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_155 TSMC_156 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_73 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_157 TSMC_158 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_74 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_159 TSMC_160 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_75 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_161 TSMC_162 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_76 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_163 TSMC_164 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_77 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_165 TSMC_166 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_78 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_167 TSMC_168 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_79 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_169 TSMC_170 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_80 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_171 TSMC_172 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_81 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_173 TSMC_174 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_82 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_175 TSMC_176 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_83 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_177 TSMC_178 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_84 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_179 TSMC_180 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_85 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_181 TSMC_182 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_86 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_183 TSMC_184 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_87 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_185 TSMC_186 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_88 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_187 TSMC_188 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_89 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_189 TSMC_190 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_90 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_191 TSMC_192 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_91 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_193 TSMC_194 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_92 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_195 TSMC_196 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_93 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_197 TSMC_198 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_94 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_199 TSMC_200 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_95 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_201 TSMC_202 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_96 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_203 TSMC_204 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_97 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_205 TSMC_206 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_98 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_207 TSMC_208 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_99 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_209 TSMC_210 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_100 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_211 TSMC_212 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_101 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_213 TSMC_214 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_102 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_215 TSMC_216 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_103 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_217 TSMC_218 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_104 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_219 TSMC_220 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_105 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_221 TSMC_222 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_106 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_223 TSMC_224 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_107 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_225 TSMC_226 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_108 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_227 TSMC_228 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_109 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_229 TSMC_230 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_110 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_231 TSMC_232 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_111 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_233 TSMC_234 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_112 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_235 TSMC_236 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_113 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_237 TSMC_238 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_114 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_239 TSMC_240 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_115 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_241 TSMC_242 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_116 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_243 TSMC_244 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_117 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_245 TSMC_246 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_118 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_247 TSMC_248 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_119 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_249 TSMC_250 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_120 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_251 TSMC_252 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_121 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_253 TSMC_254 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_122 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_255 TSMC_256 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_123 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_257 TSMC_258 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_124 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_259 TSMC_260 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_125 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_261 TSMC_262 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_126 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_263 TSMC_264 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
XMCB_127 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDAI 
+ VDDAI VDDAI TSMC_9 TSMC_10 TSMC_265 TSMC_266 
+ S1CSLVTSW400W90_MCB_2X4_SD_HD 
.ENDS

.SUBCKT S1CSLVTSW400W90_TRACKING_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 
+ TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 
+ TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 
+ TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_281 
+ TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 
+ TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_297 
+ TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 TSMC_305 
+ TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 TSMC_313 
+ TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 TSMC_320 TSMC_321 
+ TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_326 TSMC_327 TSMC_328 TSMC_329 
+ TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_337 
+ TSMC_338 TSMC_339 TSMC_340 TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_345 
+ TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_353 
+ TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_361 
+ TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 TSMC_368 TSMC_369 
+ TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 TSMC_376 TSMC_377 
+ TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 TSMC_383 TSMC_384 TSMC_385 
+ TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 TSMC_391 TSMC_392 TSMC_393 
+ TSMC_394 TSMC_395 TSMC_396 TSMC_397 TSMC_398 TSMC_399 TSMC_400 TSMC_401 
+ TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 
+ TSMC_410 TSMC_411 TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 
+ TSMC_418 TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 TSMC_433 
+ TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 TSMC_441 
+ TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 TSMC_448 TSMC_449 
+ TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 TSMC_455 TSMC_456 TSMC_457 
+ TSMC_458 TSMC_459 TSMC_460 TSMC_461 TSMC_462 TSMC_463 TSMC_464 TSMC_465 
+ TSMC_466 TSMC_467 TSMC_468 TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 
+ TSMC_474 TSMC_475 TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 
+ TSMC_482 TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 TSMC_497 
+ TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 TSMC_504 TSMC_505 
+ TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 TSMC_511 TSMC_512 TSMC_513 
+ TSMC_514 TSMC_515 TSMC_516 TSMC_517 TSMC_518 TSMC_519 TSMC_520 TSMC_521 
+ TSMC_522 TSMC_523 TSMC_524 TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 
+ TSMC_530 TSMC_531 TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 
+ TSMC_538 TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 
XTKBL_ON_CELL_0 TSMC_289 TSMC_549 TSMC_549 TSMC_291 TSMC_290 TSMC_292 TSMC_547 
+ TSMC_548 S1CSLVTSW400W90_MCB_D0734_ONCELL 
XTKBL_ON_CELL_1 TSMC_289 TSMC_549 TSMC_549 TSMC_291 TSMC_290 TSMC_292 TSMC_545 
+ TSMC_546 S1CSLVTSW400W90_MCB_D0734_ONCELL 
XTKBL_ON_CELL_2 TSMC_289 TSMC_549 TSMC_549 TSMC_291 TSMC_290 TSMC_292 TSMC_543 
+ TSMC_544 S1CSLVTSW400W90_MCB_D0734_ONCELL 
XTKBL_ON_CELL_ISO TSMC_289 TSMC_549 TSMC_549 TSMC_291 TSMC_290 TSMC_292 
+ TSMC_541 TSMC_542 TSMC_550 
+ S1CSLVTSW400W90_MCB_D0734_ONCELL_ISO 
XTKBL_OFF_CELL_4 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_539 TSMC_540 TSMC_550 
+ TSMC_551 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_5 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_537 TSMC_538 TSMC_551 
+ TSMC_552 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_6 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_535 TSMC_536 TSMC_552 
+ TSMC_553 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_7 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_533 TSMC_534 TSMC_553 
+ TSMC_554 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_8 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_531 TSMC_532 TSMC_554 
+ TSMC_555 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_9 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_529 TSMC_530 TSMC_555 
+ TSMC_556 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_10 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_527 TSMC_528 
+ TSMC_556 TSMC_557 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_11 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_525 TSMC_526 
+ TSMC_557 TSMC_558 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_12 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_523 TSMC_524 
+ TSMC_558 TSMC_559 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_13 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_521 TSMC_522 
+ TSMC_559 TSMC_560 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_14 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_519 TSMC_520 
+ TSMC_560 TSMC_561 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_15 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_517 TSMC_518 
+ TSMC_561 TSMC_562 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_16 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_515 TSMC_516 
+ TSMC_562 TSMC_563 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_17 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_513 TSMC_514 
+ TSMC_563 TSMC_564 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_18 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_511 TSMC_512 
+ TSMC_564 TSMC_565 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_19 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_509 TSMC_510 
+ TSMC_565 TSMC_566 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_20 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_507 TSMC_508 
+ TSMC_566 TSMC_567 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_21 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_505 TSMC_506 
+ TSMC_567 TSMC_568 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_22 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_503 TSMC_504 
+ TSMC_568 TSMC_569 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_23 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_501 TSMC_502 
+ TSMC_569 TSMC_570 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_24 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_499 TSMC_500 
+ TSMC_570 TSMC_571 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_25 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_497 TSMC_498 
+ TSMC_571 TSMC_572 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_26 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_495 TSMC_496 
+ TSMC_572 TSMC_573 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_27 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_493 TSMC_494 
+ TSMC_573 TSMC_574 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_28 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_491 TSMC_492 
+ TSMC_574 TSMC_575 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_29 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_489 TSMC_490 
+ TSMC_575 TSMC_576 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_30 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_487 TSMC_488 
+ TSMC_576 TSMC_577 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_31 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_485 TSMC_486 
+ TSMC_577 TSMC_578 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_32 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_483 TSMC_484 
+ TSMC_578 TSMC_579 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_33 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_481 TSMC_482 
+ TSMC_579 TSMC_580 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_34 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_479 TSMC_480 
+ TSMC_580 TSMC_581 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_35 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_477 TSMC_478 
+ TSMC_581 TSMC_582 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_36 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_475 TSMC_476 
+ TSMC_582 TSMC_583 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_37 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_473 TSMC_474 
+ TSMC_583 TSMC_584 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_38 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_471 TSMC_472 
+ TSMC_584 TSMC_585 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_39 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_469 TSMC_470 
+ TSMC_585 TSMC_586 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_40 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_467 TSMC_468 
+ TSMC_586 TSMC_587 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_41 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_465 TSMC_466 
+ TSMC_587 TSMC_588 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_42 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_463 TSMC_464 
+ TSMC_588 TSMC_589 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_43 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_461 TSMC_462 
+ TSMC_589 TSMC_590 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_44 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_459 TSMC_460 
+ TSMC_590 TSMC_591 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_45 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_457 TSMC_458 
+ TSMC_591 TSMC_592 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_46 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_455 TSMC_456 
+ TSMC_592 TSMC_593 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_47 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_453 TSMC_454 
+ TSMC_593 TSMC_594 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_48 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_451 TSMC_452 
+ TSMC_594 TSMC_595 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_49 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_449 TSMC_450 
+ TSMC_595 TSMC_596 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_50 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_447 TSMC_448 
+ TSMC_596 TSMC_597 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_51 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_445 TSMC_446 
+ TSMC_597 TSMC_598 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_52 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_443 TSMC_444 
+ TSMC_598 TSMC_599 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_53 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_441 TSMC_442 
+ TSMC_599 TSMC_600 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_54 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_439 TSMC_440 
+ TSMC_600 TSMC_601 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_55 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_437 TSMC_438 
+ TSMC_601 TSMC_602 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_56 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_435 TSMC_436 
+ TSMC_602 TSMC_603 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_57 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_433 TSMC_434 
+ TSMC_603 TSMC_604 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_58 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_431 TSMC_432 
+ TSMC_604 TSMC_605 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_59 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_429 TSMC_430 
+ TSMC_605 TSMC_606 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_60 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_427 TSMC_428 
+ TSMC_606 TSMC_607 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_61 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_425 TSMC_426 
+ TSMC_607 TSMC_608 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_62 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_423 TSMC_424 
+ TSMC_608 TSMC_609 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_63 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_421 TSMC_422 
+ TSMC_609 TSMC_610 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_64 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_419 TSMC_420 
+ TSMC_610 TSMC_611 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_65 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_417 TSMC_418 
+ TSMC_611 TSMC_612 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_66 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_415 TSMC_416 
+ TSMC_612 TSMC_613 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_67 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_413 TSMC_414 
+ TSMC_613 TSMC_614 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_68 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_411 TSMC_412 
+ TSMC_614 TSMC_615 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_69 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_409 TSMC_410 
+ TSMC_615 TSMC_616 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_70 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_407 TSMC_408 
+ TSMC_616 TSMC_617 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_71 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_405 TSMC_406 
+ TSMC_617 TSMC_618 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_72 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_403 TSMC_404 
+ TSMC_618 TSMC_619 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_73 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_401 TSMC_402 
+ TSMC_619 TSMC_620 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_74 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_399 TSMC_400 
+ TSMC_620 TSMC_621 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_75 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_397 TSMC_398 
+ TSMC_621 TSMC_622 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_76 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_395 TSMC_396 
+ TSMC_622 TSMC_623 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_77 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_393 TSMC_394 
+ TSMC_623 TSMC_624 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_78 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_391 TSMC_392 
+ TSMC_624 TSMC_625 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_79 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_389 TSMC_390 
+ TSMC_625 TSMC_626 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_80 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_387 TSMC_388 
+ TSMC_626 TSMC_627 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_81 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_385 TSMC_386 
+ TSMC_627 TSMC_628 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_82 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_383 TSMC_384 
+ TSMC_628 TSMC_629 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_83 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_381 TSMC_382 
+ TSMC_629 TSMC_630 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_84 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_379 TSMC_380 
+ TSMC_630 TSMC_631 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_85 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_377 TSMC_378 
+ TSMC_631 TSMC_632 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_86 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_375 TSMC_376 
+ TSMC_632 TSMC_633 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_87 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_373 TSMC_374 
+ TSMC_633 TSMC_634 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_88 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_371 TSMC_372 
+ TSMC_634 TSMC_635 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_89 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_369 TSMC_370 
+ TSMC_635 TSMC_636 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_90 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_367 TSMC_368 
+ TSMC_636 TSMC_637 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_91 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_365 TSMC_366 
+ TSMC_637 TSMC_638 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_92 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_363 TSMC_364 
+ TSMC_638 TSMC_639 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_93 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_361 TSMC_362 
+ TSMC_639 TSMC_640 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_94 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_359 TSMC_360 
+ TSMC_640 TSMC_641 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_95 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_357 TSMC_358 
+ TSMC_641 TSMC_642 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_96 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_355 TSMC_356 
+ TSMC_642 TSMC_643 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_97 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_353 TSMC_354 
+ TSMC_643 TSMC_644 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_98 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_351 TSMC_352 
+ TSMC_644 TSMC_645 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_99 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_349 TSMC_350 
+ TSMC_645 TSMC_646 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_100 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_347 TSMC_348 
+ TSMC_646 TSMC_647 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_101 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_345 TSMC_346 
+ TSMC_647 TSMC_648 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_102 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_343 TSMC_344 
+ TSMC_648 TSMC_649 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_103 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_341 TSMC_342 
+ TSMC_649 TSMC_650 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_104 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_339 TSMC_340 
+ TSMC_650 TSMC_651 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_105 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_337 TSMC_338 
+ TSMC_651 TSMC_652 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_106 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_335 TSMC_336 
+ TSMC_652 TSMC_653 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_107 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_333 TSMC_334 
+ TSMC_653 TSMC_654 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_108 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_331 TSMC_332 
+ TSMC_654 TSMC_655 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_109 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_329 TSMC_330 
+ TSMC_655 TSMC_656 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_110 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_327 TSMC_328 
+ TSMC_656 TSMC_657 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_111 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_325 TSMC_326 
+ TSMC_657 TSMC_658 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_112 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_323 TSMC_324 
+ TSMC_658 TSMC_659 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_113 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_321 TSMC_322 
+ TSMC_659 TSMC_660 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_114 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_319 TSMC_320 
+ TSMC_660 TSMC_661 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_115 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_317 TSMC_318 
+ TSMC_661 TSMC_662 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_116 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_315 TSMC_316 
+ TSMC_662 TSMC_663 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_117 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_313 TSMC_314 
+ TSMC_663 TSMC_664 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_118 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_311 TSMC_312 
+ TSMC_664 TSMC_665 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_119 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_309 TSMC_310 
+ TSMC_665 TSMC_666 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_120 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_307 TSMC_308 
+ TSMC_666 TSMC_667 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_121 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_305 TSMC_306 
+ TSMC_667 TSMC_668 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_122 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_303 TSMC_304 
+ TSMC_668 TSMC_669 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_123 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_301 TSMC_302 
+ TSMC_669 TSMC_670 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_124 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_299 TSMC_300 
+ TSMC_670 TSMC_671 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_125 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_297 TSMC_298 
+ TSMC_671 TSMC_672 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_126 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_295 TSMC_296 
+ TSMC_672 TSMC_673 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTKBL_OFF_CELL_127 TSMC_289 TSMC_291 TSMC_290 TSMC_292 TSMC_293 TSMC_294 
+ TSMC_673 TSMC_674 S1CSLVTSW400W90_MCB_D0734_OFFCELL 
XTRKWL_CELL_0 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_1 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_2 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_3 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_4 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_5 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_6 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_7 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_8 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_9 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_10 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_11 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_12 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_13 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_14 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_15 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_16 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_17 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_18 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_19 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_20 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_21 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_22 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_23 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_24 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_25 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_26 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_27 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_28 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_29 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_30 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_31 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_32 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_33 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_34 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
XTRKWL_CELL_35 TSMC_292 TSMC_549 TSMC_549 
+ S1CSLVTSW400W90_LOGIC_D0734_TRKWL 
.ENDS

.SUBCKT S1CSLVTSW400W90_MIO_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 
+ TSMC_18 VDD TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 TSMC_26 
+ TSMC_27 
XMIO_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 
+ TSMC_28 TSMC_11 TSMC_29 TSMC_30 TSMC_17 TSMC_18 VDD TSMC_19 TSMC_20 
+ TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 
+ S1CSLVTSW400W90_MIO_M4_SB_BASE 
XMIO_MX_SB_NBL TSMC_31 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_30 VDD VDD 
+ TSMC_19 S1CSLVTSW400W90_MIO_M4_SB_NBL_S 
XMIO_MX_SB_BUF TSMC_10 TSMC_28 TSMC_12 TSMC_29 VDD TSMC_19 
+ S1CSLVTSW400W90_MIO_M4_SB_BUF 
.ENDS

.SUBCKT S1CSLVTSW400W90_CNT_M4_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 VDD TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 
XCNT_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_73 TSMC_5 TSMC_6 TSMC_74 TSMC_7 
+ TSMC_75 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 VDD TSMC_55 TSMC_76 
+ TSMC_77 TSMC_58 TSMC_59 TSMC_60 TSMC_78 TSMC_79 TSMC_80 TSMC_81 
+ TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 TSMC_89 
+ S1CSLVTSW400W90_CNT_M4_SB_BASE 
XCNT_MX_SB_NBL TSMC_74 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 
+ TSMC_46 TSMC_47 TSMC_48 TSMC_49 VDD VDD TSMC_55 TSMC_56 TSMC_90 TSMC_77 
+ S1CSLVTSW400W90_CNT_M4_SB_NBL 
XCNT_MX_SB_BUF TSMC_4 TSMC_73 TSMC_7 TSMC_75 VDD TSMC_55 TSMC_57 TSMC_76 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 
+ TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_69 
+ TSMC_70 TSMC_71 TSMC_72 TSMC_86 TSMC_87 TSMC_88 TSMC_89 
+ S1CSLVTSW400W90_CNT_M4_SB_BUF 
.ENDS

.SUBCKT TS1N16FFCLLSBLVTC1024X144M4SW D[0] D[1] D[2] D[3] D[4] D[5] D[6] D[7] 
+ D[8] D[9] D[10] D[11] D[12] D[13] D[14] D[15] D[16] D[17] D[18] D[19] D[20] 
+ D[21] D[22] D[23] D[24] D[25] D[26] D[27] D[28] D[29] D[30] D[31] D[32] D[33] 
+ D[34] D[35] D[36] D[37] D[38] D[39] D[40] D[41] D[42] D[43] D[44] D[45] D[46] 
+ D[47] D[48] D[49] D[50] D[51] D[52] D[53] D[54] D[55] D[56] D[57] D[58] D[59] 
+ D[60] D[61] D[62] D[63] D[64] D[65] D[66] D[67] D[68] D[69] D[70] D[71] D[72] 
+ D[73] D[74] D[75] D[76] D[77] D[78] D[79] D[80] D[81] D[82] D[83] D[84] D[85] 
+ D[86] D[87] D[88] D[89] D[90] D[91] D[92] D[93] D[94] D[95] D[96] D[97] D[98] 
+ D[99] D[100] D[101] D[102] D[103] D[104] D[105] D[106] D[107] D[108] D[109] 
+ D[110] D[111] D[112] D[113] D[114] D[115] D[116] D[117] D[118] D[119] D[120] 
+ D[121] D[122] D[123] D[124] D[125] D[126] D[127] D[128] D[129] D[130] D[131] 
+ D[132] D[133] D[134] D[135] D[136] D[137] D[138] D[139] D[140] D[141] D[142] 
+ D[143] BWEB[0] BWEB[1] BWEB[2] BWEB[3] BWEB[4] BWEB[5] BWEB[6] BWEB[7] 
+ BWEB[8] BWEB[9] BWEB[10] BWEB[11] BWEB[12] BWEB[13] BWEB[14] BWEB[15] 
+ BWEB[16] BWEB[17] BWEB[18] BWEB[19] BWEB[20] BWEB[21] BWEB[22] BWEB[23] 
+ BWEB[24] BWEB[25] BWEB[26] BWEB[27] BWEB[28] BWEB[29] BWEB[30] BWEB[31] 
+ BWEB[32] BWEB[33] BWEB[34] BWEB[35] BWEB[36] BWEB[37] BWEB[38] BWEB[39] 
+ BWEB[40] BWEB[41] BWEB[42] BWEB[43] BWEB[44] BWEB[45] BWEB[46] BWEB[47] 
+ BWEB[48] BWEB[49] BWEB[50] BWEB[51] BWEB[52] BWEB[53] BWEB[54] BWEB[55] 
+ BWEB[56] BWEB[57] BWEB[58] BWEB[59] BWEB[60] BWEB[61] BWEB[62] BWEB[63] 
+ BWEB[64] BWEB[65] BWEB[66] BWEB[67] BWEB[68] BWEB[69] BWEB[70] BWEB[71] 
+ BWEB[72] BWEB[73] BWEB[74] BWEB[75] BWEB[76] BWEB[77] BWEB[78] BWEB[79] 
+ BWEB[80] BWEB[81] BWEB[82] BWEB[83] BWEB[84] BWEB[85] BWEB[86] BWEB[87] 
+ BWEB[88] BWEB[89] BWEB[90] BWEB[91] BWEB[92] BWEB[93] BWEB[94] BWEB[95] 
+ BWEB[96] BWEB[97] BWEB[98] BWEB[99] BWEB[100] BWEB[101] BWEB[102] BWEB[103] 
+ BWEB[104] BWEB[105] BWEB[106] BWEB[107] BWEB[108] BWEB[109] BWEB[110] 
+ BWEB[111] BWEB[112] BWEB[113] BWEB[114] BWEB[115] BWEB[116] BWEB[117] 
+ BWEB[118] BWEB[119] BWEB[120] BWEB[121] BWEB[122] BWEB[123] BWEB[124] 
+ BWEB[125] BWEB[126] BWEB[127] BWEB[128] BWEB[129] BWEB[130] BWEB[131] 
+ BWEB[132] BWEB[133] BWEB[134] BWEB[135] BWEB[136] BWEB[137] BWEB[138] 
+ BWEB[139] BWEB[140] BWEB[141] BWEB[142] BWEB[143] A[0] A[1] A[2] A[3] A[4] 
+ A[5] A[6] A[7] A[8] A[9] Q[0] Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] 
+ Q[10] Q[11] Q[12] Q[13] Q[14] Q[15] Q[16] Q[17] Q[18] Q[19] Q[20] Q[21] Q[22] 
+ Q[23] Q[24] Q[25] Q[26] Q[27] Q[28] Q[29] Q[30] Q[31] Q[32] Q[33] Q[34] Q[35] 
+ Q[36] Q[37] Q[38] Q[39] Q[40] Q[41] Q[42] Q[43] Q[44] Q[45] Q[46] Q[47] Q[48] 
+ Q[49] Q[50] Q[51] Q[52] Q[53] Q[54] Q[55] Q[56] Q[57] Q[58] Q[59] Q[60] Q[61] 
+ Q[62] Q[63] Q[64] Q[65] Q[66] Q[67] Q[68] Q[69] Q[70] Q[71] Q[72] Q[73] Q[74] 
+ Q[75] Q[76] Q[77] Q[78] Q[79] Q[80] Q[81] Q[82] Q[83] Q[84] Q[85] Q[86] Q[87] 
+ Q[88] Q[89] Q[90] Q[91] Q[92] Q[93] Q[94] Q[95] Q[96] Q[97] Q[98] Q[99] 
+ Q[100] Q[101] Q[102] Q[103] Q[104] Q[105] Q[106] Q[107] Q[108] Q[109] Q[110] 
+ Q[111] Q[112] Q[113] Q[114] Q[115] Q[116] Q[117] Q[118] Q[119] Q[120] Q[121] 
+ Q[122] Q[123] Q[124] Q[125] Q[126] Q[127] Q[128] Q[129] Q[130] Q[131] Q[132] 
+ Q[133] Q[134] Q[135] Q[136] Q[137] Q[138] Q[139] Q[140] Q[141] Q[142] Q[143] 
+ CEB CLK WEB RTSEL[1] RTSEL[0] WTSEL[1] WTSEL[0] VDD VSS 
XMCB256X4_L_0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDD VDD 
+ VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 
+ TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 
+ TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 
+ TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 
+ TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 
+ TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 
+ TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 
+ TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 
+ TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 
+ TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 
+ TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 TSMC_131 TSMC_132 
+ TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_139 
+ TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 
+ TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 
+ TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 
+ TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 
+ TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 
+ TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 TSMC_187 TSMC_188 
+ TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 TSMC_194 TSMC_195 
+ TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 
+ TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 
+ TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 
+ TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 
+ TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 TSMC_236 TSMC_237 
+ TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 TSMC_243 TSMC_244 
+ TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 TSMC_250 TSMC_251 
+ TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 TSMC_258 
+ TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_1 TSMC_265 TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 
+ TSMC_272 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_2 TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 
+ TSMC_280 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_3 TSMC_281 TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 
+ TSMC_288 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_4 TSMC_289 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 
+ TSMC_296 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_5 TSMC_297 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 
+ TSMC_304 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_6 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 
+ TSMC_312 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_7 TSMC_313 TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 
+ TSMC_320 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_8 TSMC_321 TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_326 TSMC_327 
+ TSMC_328 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_9 TSMC_329 TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 TSMC_335 
+ TSMC_336 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_10 TSMC_337 TSMC_338 TSMC_339 TSMC_340 TSMC_341 TSMC_342 TSMC_343 
+ TSMC_344 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_11 TSMC_345 TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 
+ TSMC_352 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_12 TSMC_353 TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 
+ TSMC_360 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_13 TSMC_361 TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 
+ TSMC_368 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_14 TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 
+ TSMC_376 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_15 TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 TSMC_383 
+ TSMC_384 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_16 TSMC_385 TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 TSMC_391 
+ TSMC_392 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_17 TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 TSMC_398 TSMC_399 
+ TSMC_400 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_18 TSMC_401 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_407 
+ TSMC_408 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_19 TSMC_409 TSMC_410 TSMC_411 TSMC_412 TSMC_413 TSMC_414 TSMC_415 
+ TSMC_416 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_20 TSMC_417 TSMC_418 TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 
+ TSMC_424 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_21 TSMC_425 TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 
+ TSMC_432 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_22 TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 
+ TSMC_440 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_23 TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_24 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 TSMC_455 
+ TSMC_456 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_25 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 TSMC_462 
+ TSMC_463 TSMC_464 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_26 TSMC_465 TSMC_466 TSMC_467 TSMC_468 TSMC_469 TSMC_470 
+ TSMC_471 TSMC_472 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_27 TSMC_473 TSMC_474 TSMC_475 TSMC_476 TSMC_477 TSMC_478 
+ TSMC_479 TSMC_480 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_28 TSMC_481 TSMC_482 TSMC_483 TSMC_484 TSMC_485 TSMC_486 
+ TSMC_487 TSMC_488 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_29 TSMC_489 TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 
+ TSMC_495 TSMC_496 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_30 TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 
+ TSMC_503 TSMC_504 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_31 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_32 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 TSMC_518 
+ TSMC_519 TSMC_520 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_33 TSMC_521 TSMC_522 TSMC_523 TSMC_524 TSMC_525 TSMC_526 
+ TSMC_527 TSMC_528 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_34 TSMC_529 TSMC_530 TSMC_531 TSMC_532 TSMC_533 TSMC_534 
+ TSMC_535 TSMC_536 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_35 TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 TSMC_542 
+ TSMC_543 TSMC_544 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_36 TSMC_545 TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 
+ TSMC_551 TSMC_552 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_37 TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 
+ TSMC_559 TSMC_560 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_38 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_39 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 TSMC_574 
+ TSMC_575 TSMC_576 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_40 TSMC_577 TSMC_578 TSMC_579 TSMC_580 TSMC_581 TSMC_582 
+ TSMC_583 TSMC_584 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_41 TSMC_585 TSMC_586 TSMC_587 TSMC_588 TSMC_589 TSMC_590 
+ TSMC_591 TSMC_592 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_42 TSMC_593 TSMC_594 TSMC_595 TSMC_596 TSMC_597 TSMC_598 
+ TSMC_599 TSMC_600 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_43 TSMC_601 TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 
+ TSMC_607 TSMC_608 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_44 TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 
+ TSMC_615 TSMC_616 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_45 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_46 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 TSMC_630 
+ TSMC_631 TSMC_632 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_47 TSMC_633 TSMC_634 TSMC_635 TSMC_636 TSMC_637 TSMC_638 
+ TSMC_639 TSMC_640 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_48 TSMC_641 TSMC_642 TSMC_643 TSMC_644 TSMC_645 TSMC_646 
+ TSMC_647 TSMC_648 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_49 TSMC_649 TSMC_650 TSMC_651 TSMC_652 TSMC_653 TSMC_654 
+ TSMC_655 TSMC_656 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_50 TSMC_657 TSMC_658 TSMC_659 TSMC_660 TSMC_661 TSMC_662 
+ TSMC_663 TSMC_664 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_51 TSMC_665 TSMC_666 TSMC_667 TSMC_668 TSMC_669 TSMC_670 
+ TSMC_671 TSMC_672 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_52 TSMC_673 TSMC_674 TSMC_675 TSMC_676 TSMC_677 TSMC_678 
+ TSMC_679 TSMC_680 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_53 TSMC_681 TSMC_682 TSMC_683 TSMC_684 TSMC_685 TSMC_686 
+ TSMC_687 TSMC_688 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_54 TSMC_689 TSMC_690 TSMC_691 TSMC_692 TSMC_693 TSMC_694 
+ TSMC_695 TSMC_696 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_55 TSMC_697 TSMC_698 TSMC_699 TSMC_700 TSMC_701 TSMC_702 
+ TSMC_703 TSMC_704 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_56 TSMC_705 TSMC_706 TSMC_707 TSMC_708 TSMC_709 TSMC_710 
+ TSMC_711 TSMC_712 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_57 TSMC_713 TSMC_714 TSMC_715 TSMC_716 TSMC_717 TSMC_718 
+ TSMC_719 TSMC_720 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_58 TSMC_721 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_727 TSMC_728 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_59 TSMC_729 TSMC_730 TSMC_731 TSMC_732 TSMC_733 TSMC_734 
+ TSMC_735 TSMC_736 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_60 TSMC_737 TSMC_738 TSMC_739 TSMC_740 TSMC_741 TSMC_742 
+ TSMC_743 TSMC_744 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_61 TSMC_745 TSMC_746 TSMC_747 TSMC_748 TSMC_749 TSMC_750 
+ TSMC_751 TSMC_752 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_62 TSMC_753 TSMC_754 TSMC_755 TSMC_756 TSMC_757 TSMC_758 
+ TSMC_759 TSMC_760 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_63 TSMC_761 TSMC_762 TSMC_763 TSMC_764 TSMC_765 TSMC_766 
+ TSMC_767 TSMC_768 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_64 TSMC_769 TSMC_770 TSMC_771 TSMC_772 TSMC_773 TSMC_774 
+ TSMC_775 TSMC_776 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_65 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 TSMC_782 
+ TSMC_783 TSMC_784 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_66 TSMC_785 TSMC_786 TSMC_787 TSMC_788 TSMC_789 TSMC_790 
+ TSMC_791 TSMC_792 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_67 TSMC_793 TSMC_794 TSMC_795 TSMC_796 TSMC_797 TSMC_798 
+ TSMC_799 TSMC_800 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_68 TSMC_801 TSMC_802 TSMC_803 TSMC_804 TSMC_805 TSMC_806 
+ TSMC_807 TSMC_808 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_69 TSMC_809 TSMC_810 TSMC_811 TSMC_812 TSMC_813 TSMC_814 
+ TSMC_815 TSMC_816 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_70 TSMC_817 TSMC_818 TSMC_819 TSMC_820 TSMC_821 TSMC_822 
+ TSMC_823 TSMC_824 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_L_71 TSMC_825 TSMC_826 TSMC_827 TSMC_828 TSMC_829 TSMC_830 
+ TSMC_831 TSMC_832 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_72 TSMC_833 TSMC_834 TSMC_835 TSMC_836 TSMC_837 TSMC_838 
+ TSMC_839 TSMC_840 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 TSMC_845 
+ TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 TSMC_852 
+ TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 TSMC_859 
+ TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 TSMC_866 
+ TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 TSMC_873 
+ TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 TSMC_880 
+ TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 TSMC_895 
+ TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 TSMC_902 
+ TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 TSMC_909 
+ TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 TSMC_916 
+ TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 TSMC_923 
+ TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 TSMC_930 
+ TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 TSMC_937 
+ TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 TSMC_944 
+ TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 TSMC_951 
+ TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 TSMC_958 
+ TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 TSMC_965 
+ TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 TSMC_972 
+ TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 TSMC_979 
+ TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 TSMC_986 
+ TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 TSMC_993 
+ TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 TSMC_1000 
+ TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 TSMC_1013 
+ TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 TSMC_1019 
+ TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 TSMC_1025 
+ TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 TSMC_1031 
+ TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 TSMC_1037 
+ TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 TSMC_1043 
+ TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 TSMC_1049 
+ TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 TSMC_1062 
+ TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 TSMC_1068 
+ TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 TSMC_1074 
+ TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 TSMC_1080 
+ TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 TSMC_1086 
+ TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 TSMC_1092 
+ TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_73 TSMC_1097 TSMC_1098 TSMC_1099 TSMC_1100 TSMC_1101 TSMC_1102 
+ TSMC_1103 TSMC_1104 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_74 TSMC_1105 TSMC_1106 TSMC_1107 TSMC_1108 TSMC_1109 TSMC_1110 
+ TSMC_1111 TSMC_1112 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_75 TSMC_1113 TSMC_1114 TSMC_1115 TSMC_1116 TSMC_1117 TSMC_1118 
+ TSMC_1119 TSMC_1120 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_76 TSMC_1121 TSMC_1122 TSMC_1123 TSMC_1124 TSMC_1125 TSMC_1126 
+ TSMC_1127 TSMC_1128 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_77 TSMC_1129 TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 
+ TSMC_1135 TSMC_1136 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_78 TSMC_1137 TSMC_1138 TSMC_1139 TSMC_1140 TSMC_1141 TSMC_1142 
+ TSMC_1143 TSMC_1144 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_79 TSMC_1145 TSMC_1146 TSMC_1147 TSMC_1148 TSMC_1149 TSMC_1150 
+ TSMC_1151 TSMC_1152 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_80 TSMC_1153 TSMC_1154 TSMC_1155 TSMC_1156 TSMC_1157 TSMC_1158 
+ TSMC_1159 TSMC_1160 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_81 TSMC_1161 TSMC_1162 TSMC_1163 TSMC_1164 TSMC_1165 TSMC_1166 
+ TSMC_1167 TSMC_1168 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_82 TSMC_1169 TSMC_1170 TSMC_1171 TSMC_1172 TSMC_1173 TSMC_1174 
+ TSMC_1175 TSMC_1176 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_83 TSMC_1177 TSMC_1178 TSMC_1179 TSMC_1180 TSMC_1181 TSMC_1182 
+ TSMC_1183 TSMC_1184 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_84 TSMC_1185 TSMC_1186 TSMC_1187 TSMC_1188 TSMC_1189 TSMC_1190 
+ TSMC_1191 TSMC_1192 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_85 TSMC_1193 TSMC_1194 TSMC_1195 TSMC_1196 TSMC_1197 TSMC_1198 
+ TSMC_1199 TSMC_1200 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_86 TSMC_1201 TSMC_1202 TSMC_1203 TSMC_1204 TSMC_1205 TSMC_1206 
+ TSMC_1207 TSMC_1208 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_87 TSMC_1209 TSMC_1210 TSMC_1211 TSMC_1212 TSMC_1213 TSMC_1214 
+ TSMC_1215 TSMC_1216 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_88 TSMC_1217 TSMC_1218 TSMC_1219 TSMC_1220 TSMC_1221 TSMC_1222 
+ TSMC_1223 TSMC_1224 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_89 TSMC_1225 TSMC_1226 TSMC_1227 TSMC_1228 TSMC_1229 TSMC_1230 
+ TSMC_1231 TSMC_1232 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_90 TSMC_1233 TSMC_1234 TSMC_1235 TSMC_1236 TSMC_1237 TSMC_1238 
+ TSMC_1239 TSMC_1240 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_91 TSMC_1241 TSMC_1242 TSMC_1243 TSMC_1244 TSMC_1245 TSMC_1246 
+ TSMC_1247 TSMC_1248 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_92 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_93 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 TSMC_1261 TSMC_1262 
+ TSMC_1263 TSMC_1264 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_94 TSMC_1265 TSMC_1266 TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 
+ TSMC_1271 TSMC_1272 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_95 TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_96 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_97 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 TSMC_1294 
+ TSMC_1295 TSMC_1296 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_98 TSMC_1297 TSMC_1298 TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 
+ TSMC_1303 TSMC_1304 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_99 TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_100 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_101 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 TSMC_1326 
+ TSMC_1327 TSMC_1328 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_102 TSMC_1329 TSMC_1330 TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 
+ TSMC_1335 TSMC_1336 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_103 TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 
+ TSMC_1343 TSMC_1344 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_104 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_105 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 TSMC_1358 
+ TSMC_1359 TSMC_1360 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_106 TSMC_1361 TSMC_1362 TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 
+ TSMC_1367 TSMC_1368 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_107 TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_108 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 
+ TSMC_1383 TSMC_1384 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_109 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 TSMC_1389 TSMC_1390 
+ TSMC_1391 TSMC_1392 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_110 TSMC_1393 TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 
+ TSMC_1399 TSMC_1400 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_111 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_112 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 TSMC_1414 
+ TSMC_1415 TSMC_1416 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_113 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 
+ TSMC_1423 TSMC_1424 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_114 TSMC_1425 TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 
+ TSMC_1431 TSMC_1432 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_115 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_116 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 TSMC_1446 
+ TSMC_1447 TSMC_1448 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_117 TSMC_1449 TSMC_1450 TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 
+ TSMC_1455 TSMC_1456 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_118 TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_119 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_120 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 TSMC_1477 TSMC_1478 
+ TSMC_1479 TSMC_1480 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_121 TSMC_1481 TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 
+ TSMC_1487 TSMC_1488 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_122 TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_123 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 TSMC_1502 
+ TSMC_1503 TSMC_1504 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_124 TSMC_1505 TSMC_1506 TSMC_1507 TSMC_1508 TSMC_1509 TSMC_1510 
+ TSMC_1511 TSMC_1512 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_125 TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 
+ TSMC_1519 TSMC_1520 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_126 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_127 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 TSMC_1534 
+ TSMC_1535 TSMC_1536 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_128 TSMC_1537 TSMC_1538 TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 
+ TSMC_1543 TSMC_1544 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_129 TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_130 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_131 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 TSMC_1565 TSMC_1566 
+ TSMC_1567 TSMC_1568 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_132 TSMC_1569 TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 
+ TSMC_1575 TSMC_1576 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_133 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_134 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 TSMC_1590 
+ TSMC_1591 TSMC_1592 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_135 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 
+ TSMC_1599 TSMC_1600 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_136 TSMC_1601 TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 
+ TSMC_1607 TSMC_1608 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_137 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 
+ TSMC_1615 TSMC_1616 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_138 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 TSMC_1622 
+ TSMC_1623 TSMC_1624 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_139 TSMC_1625 TSMC_1626 TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 
+ TSMC_1631 TSMC_1632 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_140 TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_141 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_142 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 TSMC_1653 TSMC_1654 
+ TSMC_1655 TSMC_1656 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XMCB256X4_R_143 TSMC_1657 TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 
+ TSMC_1663 TSMC_1664 VDD VDD VSS TSMC_841 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 
+ TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 
+ TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 
+ TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_985 
+ TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 
+ TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 
+ TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 
+ TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 
+ TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ S1CSLVTSW400W90_MCB_ARR 
XXDRV_STRAP_BT_SB_0 TSMC_1665 TSMC_1666 VDD VSS 
+ S1CSLVTSW400W90_XDRV_STRAP_BT_SB 
XXDRV_LA512_SB_0 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 
+ TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_841 
+ TSMC_842 TSMC_843 TSMC_844 TSMC_1665 TSMC_1666 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_1 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1675 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 VDD VSS TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_845 
+ TSMC_846 TSMC_847 TSMC_848 TSMC_1665 TSMC_1666 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_2 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1704 
+ TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 TSMC_1710 
+ TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 TSMC_1716 
+ TSMC_1717 TSMC_1718 VDD VSS TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_849 
+ TSMC_850 TSMC_851 TSMC_852 TSMC_1665 TSMC_1666 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_3 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1719 
+ TSMC_1720 TSMC_1721 TSMC_1722 TSMC_1708 TSMC_1723 TSMC_1724 
+ TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 TSMC_1729 TSMC_1730 
+ TSMC_1731 TSMC_1732 VDD VSS TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_853 
+ TSMC_854 TSMC_855 TSMC_856 TSMC_1665 TSMC_1666 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_4 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 
+ TSMC_1746 TSMC_1747 VDD VSS TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_857 
+ TSMC_858 TSMC_859 TSMC_860 TSMC_1665 TSMC_1666 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_5 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1748 
+ TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1737 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 VDD VSS TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_861 
+ TSMC_862 TSMC_863 TSMC_864 TSMC_1665 TSMC_1666 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_6 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1762 
+ TSMC_1763 TSMC_1764 TSMC_1765 TSMC_1766 TSMC_1767 TSMC_1768 
+ TSMC_1769 TSMC_1770 TSMC_1771 TSMC_1772 TSMC_1773 TSMC_1774 
+ TSMC_1775 TSMC_1776 VDD VSS TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_1665 TSMC_1666 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_7 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1777 
+ TSMC_1778 TSMC_1779 TSMC_1780 TSMC_1766 TSMC_1781 TSMC_1782 
+ TSMC_1783 TSMC_1784 TSMC_1785 TSMC_1786 TSMC_1787 TSMC_1788 
+ TSMC_1789 TSMC_1790 VDD VSS TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_869 
+ TSMC_870 TSMC_871 TSMC_872 TSMC_1665 TSMC_1666 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_8 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1791 
+ TSMC_1792 TSMC_1793 TSMC_1794 TSMC_1795 TSMC_1796 TSMC_1797 
+ TSMC_1798 TSMC_1799 TSMC_1800 TSMC_1801 TSMC_1802 TSMC_1803 
+ TSMC_1804 TSMC_1805 VDD VSS TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_873 
+ TSMC_874 TSMC_875 TSMC_876 TSMC_1665 TSMC_1666 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_9 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1806 
+ TSMC_1807 TSMC_1808 TSMC_1809 TSMC_1795 TSMC_1810 TSMC_1811 
+ TSMC_1812 TSMC_1813 TSMC_1814 TSMC_1815 TSMC_1816 TSMC_1817 
+ TSMC_1818 TSMC_1819 VDD VSS TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_877 
+ TSMC_878 TSMC_879 TSMC_880 TSMC_1665 TSMC_1666 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_10 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1820 
+ TSMC_1821 TSMC_1822 TSMC_1823 TSMC_1824 TSMC_1825 TSMC_1826 
+ TSMC_1827 TSMC_1828 TSMC_1829 TSMC_1830 TSMC_1831 TSMC_1832 
+ TSMC_1833 TSMC_1834 VDD VSS TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_1665 TSMC_1666 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_11 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1835 
+ TSMC_1836 TSMC_1837 TSMC_1838 TSMC_1824 TSMC_1839 TSMC_1840 
+ TSMC_1841 TSMC_1842 TSMC_1843 TSMC_1844 TSMC_1845 TSMC_1846 
+ TSMC_1847 TSMC_1848 VDD VSS TSMC_53 TSMC_54 TSMC_55 TSMC_56 
+ TSMC_885 TSMC_886 TSMC_887 TSMC_888 TSMC_1665 TSMC_1666 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_12 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1849 
+ TSMC_1850 TSMC_1851 TSMC_1852 TSMC_1853 TSMC_1854 TSMC_1855 
+ TSMC_1856 TSMC_1857 TSMC_1858 TSMC_1859 TSMC_1860 TSMC_1861 
+ TSMC_1862 TSMC_1863 VDD VSS TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_1665 TSMC_1666 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_13 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1864 
+ TSMC_1865 TSMC_1866 TSMC_1867 TSMC_1853 TSMC_1868 TSMC_1869 
+ TSMC_1870 TSMC_1871 TSMC_1872 TSMC_1873 TSMC_1874 TSMC_1875 
+ TSMC_1876 TSMC_1877 VDD VSS TSMC_61 TSMC_62 TSMC_63 TSMC_64 
+ TSMC_893 TSMC_894 TSMC_895 TSMC_896 TSMC_1665 TSMC_1666 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_14 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1878 
+ TSMC_1879 TSMC_1880 TSMC_1881 TSMC_1882 TSMC_1883 TSMC_1884 
+ TSMC_1885 TSMC_1886 TSMC_1887 TSMC_1888 TSMC_1889 TSMC_1890 
+ TSMC_1891 TSMC_1892 VDD VSS TSMC_65 TSMC_66 TSMC_67 TSMC_68 
+ TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_1665 TSMC_1666 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_15 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1893 
+ TSMC_1894 TSMC_1895 TSMC_1896 TSMC_1882 TSMC_1897 TSMC_1898 
+ TSMC_1899 TSMC_1900 TSMC_1901 TSMC_1902 TSMC_1903 TSMC_1904 
+ TSMC_1905 TSMC_1906 VDD VSS TSMC_69 TSMC_70 TSMC_71 TSMC_72 
+ TSMC_901 TSMC_902 TSMC_903 TSMC_904 TSMC_1665 TSMC_1666 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_STRAP_SB_16 TSMC_1907 TSMC_1908 VDD VSS 
+ S1CSLVTSW400W90_XDRV_STRAP_SB 
XXDRV_LA512_SB_16 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1909 
+ TSMC_1910 TSMC_1911 TSMC_1912 TSMC_1675 TSMC_1913 TSMC_1914 
+ TSMC_1915 TSMC_1916 TSMC_1917 TSMC_1918 TSMC_1919 TSMC_1920 
+ TSMC_1921 TSMC_1922 VDD VSS TSMC_73 TSMC_74 TSMC_75 TSMC_76 
+ TSMC_905 TSMC_906 TSMC_907 TSMC_908 TSMC_1907 TSMC_1908 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_17 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1923 
+ TSMC_1924 TSMC_1925 TSMC_1926 TSMC_1675 TSMC_1927 TSMC_1928 
+ TSMC_1929 TSMC_1930 TSMC_1931 TSMC_1932 TSMC_1933 TSMC_1934 
+ TSMC_1935 TSMC_1936 VDD VSS TSMC_77 TSMC_78 TSMC_79 TSMC_80 
+ TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_1907 TSMC_1908 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_18 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1937 
+ TSMC_1938 TSMC_1939 TSMC_1940 TSMC_1708 TSMC_1941 TSMC_1942 
+ TSMC_1943 TSMC_1944 TSMC_1945 TSMC_1946 TSMC_1947 TSMC_1948 
+ TSMC_1949 TSMC_1950 VDD VSS TSMC_81 TSMC_82 TSMC_83 TSMC_84 
+ TSMC_913 TSMC_914 TSMC_915 TSMC_916 TSMC_1907 TSMC_1908 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_19 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1951 
+ TSMC_1952 TSMC_1953 TSMC_1954 TSMC_1708 TSMC_1955 TSMC_1956 
+ TSMC_1957 TSMC_1958 TSMC_1959 TSMC_1960 TSMC_1961 TSMC_1962 
+ TSMC_1963 TSMC_1964 VDD VSS TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_1907 TSMC_1908 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_20 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1965 
+ TSMC_1966 TSMC_1967 TSMC_1968 TSMC_1737 TSMC_1969 TSMC_1970 
+ TSMC_1971 TSMC_1972 TSMC_1973 TSMC_1974 TSMC_1975 TSMC_1976 
+ TSMC_1977 TSMC_1978 VDD VSS TSMC_89 TSMC_90 TSMC_91 TSMC_92 
+ TSMC_921 TSMC_922 TSMC_923 TSMC_924 TSMC_1907 TSMC_1908 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_21 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1979 
+ TSMC_1980 TSMC_1981 TSMC_1982 TSMC_1737 TSMC_1983 TSMC_1984 
+ TSMC_1985 TSMC_1986 TSMC_1987 TSMC_1988 TSMC_1989 TSMC_1990 
+ TSMC_1991 TSMC_1992 VDD VSS TSMC_93 TSMC_94 TSMC_95 TSMC_96 
+ TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_1907 TSMC_1908 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_22 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1993 
+ TSMC_1994 TSMC_1995 TSMC_1996 TSMC_1766 TSMC_1997 TSMC_1998 
+ TSMC_1999 TSMC_2000 TSMC_2001 TSMC_2002 TSMC_2003 TSMC_2004 
+ TSMC_2005 TSMC_2006 VDD VSS TSMC_97 TSMC_98 TSMC_99 TSMC_100 
+ TSMC_929 TSMC_930 TSMC_931 TSMC_932 TSMC_1907 TSMC_1908 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_23 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2007 
+ TSMC_2008 TSMC_2009 TSMC_2010 TSMC_1766 TSMC_2011 TSMC_2012 
+ TSMC_2013 TSMC_2014 TSMC_2015 TSMC_2016 TSMC_2017 TSMC_2018 
+ TSMC_2019 TSMC_2020 VDD VSS TSMC_101 TSMC_102 TSMC_103 TSMC_104 
+ TSMC_933 TSMC_934 TSMC_935 TSMC_936 TSMC_1907 TSMC_1908 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_24 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2021 
+ TSMC_2022 TSMC_2023 TSMC_2024 TSMC_1795 TSMC_2025 TSMC_2026 
+ TSMC_2027 TSMC_2028 TSMC_2029 TSMC_2030 TSMC_2031 TSMC_2032 
+ TSMC_2033 TSMC_2034 VDD VSS TSMC_105 TSMC_106 TSMC_107 TSMC_108 
+ TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_1907 TSMC_1908 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_25 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2035 
+ TSMC_2036 TSMC_2037 TSMC_2038 TSMC_1795 TSMC_2039 TSMC_2040 
+ TSMC_2041 TSMC_2042 TSMC_2043 TSMC_2044 TSMC_2045 TSMC_2046 
+ TSMC_2047 TSMC_2048 VDD VSS TSMC_109 TSMC_110 TSMC_111 TSMC_112 
+ TSMC_941 TSMC_942 TSMC_943 TSMC_944 TSMC_1907 TSMC_1908 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_26 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2049 
+ TSMC_2050 TSMC_2051 TSMC_2052 TSMC_1824 TSMC_2053 TSMC_2054 
+ TSMC_2055 TSMC_2056 TSMC_2057 TSMC_2058 TSMC_2059 TSMC_2060 
+ TSMC_2061 TSMC_2062 VDD VSS TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_1907 TSMC_1908 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_27 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2063 
+ TSMC_2064 TSMC_2065 TSMC_2066 TSMC_1824 TSMC_2067 TSMC_2068 
+ TSMC_2069 TSMC_2070 TSMC_2071 TSMC_2072 TSMC_2073 TSMC_2074 
+ TSMC_2075 TSMC_2076 VDD VSS TSMC_117 TSMC_118 TSMC_119 TSMC_120 
+ TSMC_949 TSMC_950 TSMC_951 TSMC_952 TSMC_1907 TSMC_1908 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_28 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2077 
+ TSMC_2078 TSMC_2079 TSMC_2080 TSMC_1853 TSMC_2081 TSMC_2082 
+ TSMC_2083 TSMC_2084 TSMC_2085 TSMC_2086 TSMC_2087 TSMC_2088 
+ TSMC_2089 TSMC_2090 VDD VSS TSMC_121 TSMC_122 TSMC_123 TSMC_124 
+ TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_1907 TSMC_1908 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_29 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2091 
+ TSMC_2092 TSMC_2093 TSMC_2094 TSMC_1853 TSMC_2095 TSMC_2096 
+ TSMC_2097 TSMC_2098 TSMC_2099 TSMC_2100 TSMC_2101 TSMC_2102 
+ TSMC_2103 TSMC_2104 VDD VSS TSMC_125 TSMC_126 TSMC_127 TSMC_128 
+ TSMC_957 TSMC_958 TSMC_959 TSMC_960 TSMC_1907 TSMC_1908 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_30 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2105 
+ TSMC_2106 TSMC_2107 TSMC_2108 TSMC_1882 TSMC_2109 TSMC_2110 
+ TSMC_2111 TSMC_2112 TSMC_2113 TSMC_2114 TSMC_2115 TSMC_2116 
+ TSMC_2117 TSMC_2118 VDD VSS TSMC_129 TSMC_130 TSMC_131 TSMC_132 
+ TSMC_961 TSMC_962 TSMC_963 TSMC_964 TSMC_1907 TSMC_1908 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_31 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2119 
+ TSMC_2120 TSMC_2121 TSMC_2122 TSMC_1882 TSMC_2123 TSMC_2124 
+ TSMC_2125 TSMC_2126 TSMC_2127 TSMC_2128 TSMC_2129 TSMC_2130 
+ TSMC_2131 TSMC_2132 VDD VSS TSMC_133 TSMC_134 TSMC_135 TSMC_136 
+ TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_1907 TSMC_1908 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_STRAP_SB_32 TSMC_2133 TSMC_2134 VDD VSS 
+ S1CSLVTSW400W90_XDRV_STRAP_SB 
XXDRV_LA512_SB_32 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2135 
+ TSMC_2136 TSMC_2137 TSMC_2138 TSMC_1675 TSMC_2139 TSMC_2140 
+ TSMC_2141 TSMC_2142 TSMC_2143 TSMC_2144 TSMC_2145 TSMC_2146 
+ TSMC_2147 TSMC_2148 VDD VSS TSMC_137 TSMC_138 TSMC_139 TSMC_140 
+ TSMC_969 TSMC_970 TSMC_971 TSMC_972 TSMC_2133 TSMC_2134 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_33 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2149 
+ TSMC_2150 TSMC_2151 TSMC_2152 TSMC_1675 TSMC_2153 TSMC_2154 
+ TSMC_2155 TSMC_2156 TSMC_2157 TSMC_2158 TSMC_2159 TSMC_2160 
+ TSMC_2161 TSMC_2162 VDD VSS TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_2133 TSMC_2134 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_34 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2163 
+ TSMC_2164 TSMC_2165 TSMC_2166 TSMC_1708 TSMC_2167 TSMC_2168 
+ TSMC_2169 TSMC_2170 TSMC_2171 TSMC_2172 TSMC_2173 TSMC_2174 
+ TSMC_2175 TSMC_2176 VDD VSS TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ TSMC_977 TSMC_978 TSMC_979 TSMC_980 TSMC_2133 TSMC_2134 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_35 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2177 
+ TSMC_2178 TSMC_2179 TSMC_2180 TSMC_1708 TSMC_2181 TSMC_2182 
+ TSMC_2183 TSMC_2184 TSMC_2185 TSMC_2186 TSMC_2187 TSMC_2188 
+ TSMC_2189 TSMC_2190 VDD VSS TSMC_149 TSMC_150 TSMC_151 TSMC_152 
+ TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_2133 TSMC_2134 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_36 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2191 
+ TSMC_2192 TSMC_2193 TSMC_2194 TSMC_1737 TSMC_2195 TSMC_2196 
+ TSMC_2197 TSMC_2198 TSMC_2199 TSMC_2200 TSMC_2201 TSMC_2202 
+ TSMC_2203 TSMC_2204 VDD VSS TSMC_153 TSMC_154 TSMC_155 TSMC_156 
+ TSMC_985 TSMC_986 TSMC_987 TSMC_988 TSMC_2133 TSMC_2134 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_37 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2205 
+ TSMC_2206 TSMC_2207 TSMC_2208 TSMC_1737 TSMC_2209 TSMC_2210 
+ TSMC_2211 TSMC_2212 TSMC_2213 TSMC_2214 TSMC_2215 TSMC_2216 
+ TSMC_2217 TSMC_2218 VDD VSS TSMC_157 TSMC_158 TSMC_159 TSMC_160 
+ TSMC_989 TSMC_990 TSMC_991 TSMC_992 TSMC_2133 TSMC_2134 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_38 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2219 
+ TSMC_2220 TSMC_2221 TSMC_2222 TSMC_1766 TSMC_2223 TSMC_2224 
+ TSMC_2225 TSMC_2226 TSMC_2227 TSMC_2228 TSMC_2229 TSMC_2230 
+ TSMC_2231 TSMC_2232 VDD VSS TSMC_161 TSMC_162 TSMC_163 TSMC_164 
+ TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_2133 TSMC_2134 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_39 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2233 
+ TSMC_2234 TSMC_2235 TSMC_2236 TSMC_1766 TSMC_2237 TSMC_2238 
+ TSMC_2239 TSMC_2240 TSMC_2241 TSMC_2242 TSMC_2243 TSMC_2244 
+ TSMC_2245 TSMC_2246 VDD VSS TSMC_165 TSMC_166 TSMC_167 TSMC_168 
+ TSMC_997 TSMC_998 TSMC_999 TSMC_1000 TSMC_2133 TSMC_2134 
+ S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_40 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2247 
+ TSMC_2248 TSMC_2249 TSMC_2250 TSMC_1795 TSMC_2251 TSMC_2252 
+ TSMC_2253 TSMC_2254 TSMC_2255 TSMC_2256 TSMC_2257 TSMC_2258 
+ TSMC_2259 TSMC_2260 VDD VSS TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_2133 
+ TSMC_2134 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_41 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2261 
+ TSMC_2262 TSMC_2263 TSMC_2264 TSMC_1795 TSMC_2265 TSMC_2266 
+ TSMC_2267 TSMC_2268 TSMC_2269 TSMC_2270 TSMC_2271 TSMC_2272 
+ TSMC_2273 TSMC_2274 VDD VSS TSMC_173 TSMC_174 TSMC_175 TSMC_176 
+ TSMC_1005 TSMC_1006 TSMC_1007 TSMC_1008 TSMC_2133 
+ TSMC_2134 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_42 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2275 
+ TSMC_2276 TSMC_2277 TSMC_2278 TSMC_1824 TSMC_2279 TSMC_2280 
+ TSMC_2281 TSMC_2282 TSMC_2283 TSMC_2284 TSMC_2285 TSMC_2286 
+ TSMC_2287 TSMC_2288 VDD VSS TSMC_177 TSMC_178 TSMC_179 TSMC_180 
+ TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 TSMC_2133 
+ TSMC_2134 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_43 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2289 
+ TSMC_2290 TSMC_2291 TSMC_2292 TSMC_1824 TSMC_2293 TSMC_2294 
+ TSMC_2295 TSMC_2296 TSMC_2297 TSMC_2298 TSMC_2299 TSMC_2300 
+ TSMC_2301 TSMC_2302 VDD VSS TSMC_181 TSMC_182 TSMC_183 TSMC_184 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_2133 
+ TSMC_2134 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_44 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2303 
+ TSMC_2304 TSMC_2305 TSMC_2306 TSMC_1853 TSMC_2307 TSMC_2308 
+ TSMC_2309 TSMC_2310 TSMC_2311 TSMC_2312 TSMC_2313 TSMC_2314 
+ TSMC_2315 TSMC_2316 VDD VSS TSMC_185 TSMC_186 TSMC_187 TSMC_188 
+ TSMC_1017 TSMC_1018 TSMC_1019 TSMC_1020 TSMC_2133 
+ TSMC_2134 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_45 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2317 
+ TSMC_2318 TSMC_2319 TSMC_2320 TSMC_1853 TSMC_2321 TSMC_2322 
+ TSMC_2323 TSMC_2324 TSMC_2325 TSMC_2326 TSMC_2327 TSMC_2328 
+ TSMC_2329 TSMC_2330 VDD VSS TSMC_189 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 TSMC_2133 
+ TSMC_2134 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_46 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2331 
+ TSMC_2332 TSMC_2333 TSMC_2334 TSMC_1882 TSMC_2335 TSMC_2336 
+ TSMC_2337 TSMC_2338 TSMC_2339 TSMC_2340 TSMC_2341 TSMC_2342 
+ TSMC_2343 TSMC_2344 VDD VSS TSMC_193 TSMC_194 TSMC_195 TSMC_196 
+ TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_2133 
+ TSMC_2134 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_47 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2345 
+ TSMC_2346 TSMC_2347 TSMC_2348 TSMC_1882 TSMC_2349 TSMC_2350 
+ TSMC_2351 TSMC_2352 TSMC_2353 TSMC_2354 TSMC_2355 TSMC_2356 
+ TSMC_2357 TSMC_2358 VDD VSS TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_1029 TSMC_1030 TSMC_1031 TSMC_1032 TSMC_2133 
+ TSMC_2134 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_STRAP_SB_48 TSMC_2359 TSMC_2360 VDD VSS 
+ S1CSLVTSW400W90_XDRV_STRAP_SB 
XXDRV_LA512_SB_48 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2361 
+ TSMC_2362 TSMC_2363 TSMC_2364 TSMC_1675 TSMC_2365 TSMC_2366 
+ TSMC_2367 TSMC_2368 TSMC_2369 TSMC_2370 TSMC_2371 TSMC_2372 
+ TSMC_2373 TSMC_2374 VDD VSS TSMC_201 TSMC_202 TSMC_203 TSMC_204 
+ TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 TSMC_2359 
+ TSMC_2360 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_49 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2375 
+ TSMC_2376 TSMC_2377 TSMC_2378 TSMC_1675 TSMC_2379 TSMC_2380 
+ TSMC_2381 TSMC_2382 TSMC_2383 TSMC_2384 TSMC_2385 TSMC_2386 
+ TSMC_2387 TSMC_2388 VDD VSS TSMC_205 TSMC_206 TSMC_207 TSMC_208 
+ TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_2359 
+ TSMC_2360 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_50 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2389 
+ TSMC_2390 TSMC_2391 TSMC_2392 TSMC_1708 TSMC_2393 TSMC_2394 
+ TSMC_2395 TSMC_2396 TSMC_2397 TSMC_2398 TSMC_2399 TSMC_2400 
+ TSMC_2401 TSMC_2402 VDD VSS TSMC_209 TSMC_210 TSMC_211 TSMC_212 
+ TSMC_1041 TSMC_1042 TSMC_1043 TSMC_1044 TSMC_2359 
+ TSMC_2360 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_51 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2403 
+ TSMC_2404 TSMC_2405 TSMC_2406 TSMC_1708 TSMC_2407 TSMC_2408 
+ TSMC_2409 TSMC_2410 TSMC_2411 TSMC_2412 TSMC_2413 TSMC_2414 
+ TSMC_2415 TSMC_2416 VDD VSS TSMC_213 TSMC_214 TSMC_215 TSMC_216 
+ TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 TSMC_2359 
+ TSMC_2360 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_52 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2417 
+ TSMC_2418 TSMC_2419 TSMC_2420 TSMC_1737 TSMC_2421 TSMC_2422 
+ TSMC_2423 TSMC_2424 TSMC_2425 TSMC_2426 TSMC_2427 TSMC_2428 
+ TSMC_2429 TSMC_2430 VDD VSS TSMC_217 TSMC_218 TSMC_219 TSMC_220 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_2359 
+ TSMC_2360 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_53 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2431 
+ TSMC_2432 TSMC_2433 TSMC_2434 TSMC_1737 TSMC_2435 TSMC_2436 
+ TSMC_2437 TSMC_2438 TSMC_2439 TSMC_2440 TSMC_2441 TSMC_2442 
+ TSMC_2443 TSMC_2444 VDD VSS TSMC_221 TSMC_222 TSMC_223 TSMC_224 
+ TSMC_1053 TSMC_1054 TSMC_1055 TSMC_1056 TSMC_2359 
+ TSMC_2360 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_54 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2445 
+ TSMC_2446 TSMC_2447 TSMC_2448 TSMC_1766 TSMC_2449 TSMC_2450 
+ TSMC_2451 TSMC_2452 TSMC_2453 TSMC_2454 TSMC_2455 TSMC_2456 
+ TSMC_2457 TSMC_2458 VDD VSS TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_2359 
+ TSMC_2360 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_55 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2459 
+ TSMC_2460 TSMC_2461 TSMC_2462 TSMC_1766 TSMC_2463 TSMC_2464 
+ TSMC_2465 TSMC_2466 TSMC_2467 TSMC_2468 TSMC_2469 TSMC_2470 
+ TSMC_2471 TSMC_2472 VDD VSS TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_1061 TSMC_1062 TSMC_1063 TSMC_1064 TSMC_2359 
+ TSMC_2360 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_56 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2473 
+ TSMC_2474 TSMC_2475 TSMC_2476 TSMC_1795 TSMC_2477 TSMC_2478 
+ TSMC_2479 TSMC_2480 TSMC_2481 TSMC_2482 TSMC_2483 TSMC_2484 
+ TSMC_2485 TSMC_2486 VDD VSS TSMC_233 TSMC_234 TSMC_235 TSMC_236 
+ TSMC_1065 TSMC_1066 TSMC_1067 TSMC_1068 TSMC_2359 
+ TSMC_2360 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_57 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2487 
+ TSMC_2488 TSMC_2489 TSMC_2490 TSMC_1795 TSMC_2491 TSMC_2492 
+ TSMC_2493 TSMC_2494 TSMC_2495 TSMC_2496 TSMC_2497 TSMC_2498 
+ TSMC_2499 TSMC_2500 VDD VSS TSMC_237 TSMC_238 TSMC_239 TSMC_240 
+ TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_2359 
+ TSMC_2360 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_58 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2501 
+ TSMC_2502 TSMC_2503 TSMC_2504 TSMC_1824 TSMC_2505 TSMC_2506 
+ TSMC_2507 TSMC_2508 TSMC_2509 TSMC_2510 TSMC_2511 TSMC_2512 
+ TSMC_2513 TSMC_2514 VDD VSS TSMC_241 TSMC_242 TSMC_243 TSMC_244 
+ TSMC_1073 TSMC_1074 TSMC_1075 TSMC_1076 TSMC_2359 
+ TSMC_2360 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_59 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2515 
+ TSMC_2516 TSMC_2517 TSMC_2518 TSMC_1824 TSMC_2519 TSMC_2520 
+ TSMC_2521 TSMC_2522 TSMC_2523 TSMC_2524 TSMC_2525 TSMC_2526 
+ TSMC_2527 TSMC_2528 VDD VSS TSMC_245 TSMC_246 TSMC_247 TSMC_248 
+ TSMC_1077 TSMC_1078 TSMC_1079 TSMC_1080 TSMC_2359 
+ TSMC_2360 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_60 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2529 
+ TSMC_2530 TSMC_2531 TSMC_2532 TSMC_1853 TSMC_2533 TSMC_2534 
+ TSMC_2535 TSMC_2536 TSMC_2537 TSMC_2538 TSMC_2539 TSMC_2540 
+ TSMC_2541 TSMC_2542 VDD VSS TSMC_249 TSMC_250 TSMC_251 TSMC_252 
+ TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_2359 
+ TSMC_2360 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_61 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2543 
+ TSMC_2544 TSMC_2545 TSMC_2546 TSMC_1853 TSMC_2547 TSMC_2548 
+ TSMC_2549 TSMC_2550 TSMC_2551 TSMC_2552 TSMC_2553 TSMC_2554 
+ TSMC_2555 TSMC_2556 VDD VSS TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_1085 TSMC_1086 TSMC_1087 TSMC_1088 TSMC_2359 
+ TSMC_2360 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_62 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_2557 
+ TSMC_2558 TSMC_2559 TSMC_2560 TSMC_1882 TSMC_2561 TSMC_2562 
+ TSMC_2563 TSMC_2564 TSMC_2565 TSMC_2566 TSMC_2567 TSMC_2568 
+ TSMC_2569 TSMC_2570 VDD VSS TSMC_257 TSMC_258 TSMC_259 TSMC_260 
+ TSMC_1089 TSMC_1090 TSMC_1091 TSMC_1092 TSMC_2359 
+ TSMC_2360 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XXDRV_LA512_SB_63 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_2571 
+ TSMC_2572 TSMC_2573 TSMC_2574 TSMC_1882 TSMC_2575 TSMC_2576 
+ TSMC_2577 TSMC_2578 TSMC_2579 TSMC_2580 TSMC_2581 TSMC_2582 
+ TSMC_2583 TSMC_2584 VDD VSS TSMC_261 TSMC_262 TSMC_263 TSMC_264 
+ TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 TSMC_2359 
+ TSMC_2360 S1CSLVTSW400W90_XDRV_LA512_884_SB 
XTRACKING_XB256X4 TSMC_833 TSMC_834 TSMC_835 TSMC_836 TSMC_1097 TSMC_1098 
+ TSMC_1099 TSMC_1100 TSMC_1105 TSMC_1106 TSMC_1107 TSMC_1108 
+ TSMC_1113 TSMC_1114 TSMC_1115 TSMC_1116 TSMC_1121 TSMC_1122 
+ TSMC_1123 TSMC_1124 TSMC_1129 TSMC_1130 TSMC_1131 TSMC_1132 
+ TSMC_1137 TSMC_1138 TSMC_1139 TSMC_1140 TSMC_1145 TSMC_1146 
+ TSMC_1147 TSMC_1148 TSMC_1153 TSMC_1154 TSMC_1155 TSMC_1156 TSMC_1161 
+ TSMC_1162 TSMC_1163 TSMC_1164 TSMC_1169 TSMC_1170 TSMC_1171 
+ TSMC_1172 TSMC_1177 TSMC_1178 TSMC_1179 TSMC_1180 TSMC_1185 
+ TSMC_1186 TSMC_1187 TSMC_1188 TSMC_1193 TSMC_1194 TSMC_1195 
+ TSMC_1196 TSMC_1201 TSMC_1202 TSMC_1203 TSMC_1204 TSMC_1209 TSMC_1210 
+ TSMC_1211 TSMC_1212 TSMC_1217 TSMC_1218 TSMC_1219 TSMC_1220 
+ TSMC_1225 TSMC_1226 TSMC_1227 TSMC_1228 TSMC_1233 TSMC_1234 
+ TSMC_1235 TSMC_1236 TSMC_1241 TSMC_1242 TSMC_1243 TSMC_1244 
+ TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1257 TSMC_1258 
+ TSMC_1259 TSMC_1260 TSMC_1265 TSMC_1266 TSMC_1267 TSMC_1268 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1281 TSMC_1282 TSMC_1283 
+ TSMC_1284 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1297 
+ TSMC_1298 TSMC_1299 TSMC_1300 TSMC_1305 TSMC_1306 TSMC_1307 
+ TSMC_1308 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1321 TSMC_1322 
+ TSMC_1323 TSMC_1324 TSMC_1329 TSMC_1330 TSMC_1331 TSMC_1332 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1345 TSMC_1346 
+ TSMC_1347 TSMC_1348 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1361 TSMC_1362 TSMC_1363 TSMC_1364 TSMC_1369 TSMC_1370 
+ TSMC_1371 TSMC_1372 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1385 
+ TSMC_1386 TSMC_1387 TSMC_1388 TSMC_1393 TSMC_1394 TSMC_1395 
+ TSMC_1396 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1409 
+ TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1425 TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1433 TSMC_1434 
+ TSMC_1435 TSMC_1436 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1449 TSMC_1450 TSMC_1451 TSMC_1452 TSMC_1457 TSMC_1458 
+ TSMC_1459 TSMC_1460 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 
+ TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1497 
+ TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1505 TSMC_1506 TSMC_1507 
+ TSMC_1508 TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1521 
+ TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1537 TSMC_1538 TSMC_1539 TSMC_1540 TSMC_1545 TSMC_1546 
+ TSMC_1547 TSMC_1548 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 
+ TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 
+ TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1601 TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1609 
+ TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1617 TSMC_1618 TSMC_1619 
+ TSMC_1620 TSMC_1625 TSMC_1626 TSMC_1627 TSMC_1628 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1641 TSMC_1642 TSMC_1643 
+ TSMC_1644 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 TSMC_1657 TSMC_1658 
+ TSMC_1659 TSMC_1660 TSMC_2585 VDD VDD VSS TSMC_841 TSMC_842 
+ TSMC_843 TSMC_844 TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 
+ TSMC_850 TSMC_851 TSMC_852 TSMC_853 TSMC_854 TSMC_855 TSMC_856 
+ TSMC_857 TSMC_858 TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 
+ TSMC_864 TSMC_865 TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 
+ TSMC_871 TSMC_872 TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 
+ TSMC_879 TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 
+ TSMC_886 TSMC_887 TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 
+ TSMC_893 TSMC_894 TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 
+ TSMC_900 TSMC_901 TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 
+ TSMC_907 TSMC_908 TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 
+ TSMC_914 TSMC_915 TSMC_916 TSMC_917 TSMC_918 TSMC_919 TSMC_920 
+ TSMC_921 TSMC_922 TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 
+ TSMC_928 TSMC_929 TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 
+ TSMC_935 TSMC_936 TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 
+ TSMC_943 TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 
+ TSMC_950 TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 
+ TSMC_957 TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 
+ TSMC_964 TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 
+ TSMC_971 TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 
+ TSMC_978 TSMC_979 TSMC_980 TSMC_981 TSMC_982 TSMC_983 TSMC_984 
+ TSMC_985 TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 
+ TSMC_992 TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 
+ TSMC_999 TSMC_1000 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 
+ TSMC_1006 TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 
+ TSMC_1012 TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 
+ TSMC_1018 TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 
+ TSMC_1024 TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 
+ TSMC_1030 TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 TSMC_1035 
+ TSMC_1036 TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 
+ TSMC_1042 TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 TSMC_1047 
+ TSMC_1048 TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 
+ TSMC_1055 TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 
+ TSMC_1061 TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 
+ TSMC_1067 TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 
+ TSMC_1073 TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 
+ TSMC_1079 TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 TSMC_1084 
+ TSMC_1085 TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 
+ TSMC_1091 TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 TSMC_1096 
+ TSMC_2586 S1CSLVTSW400W90_TRACKING_SB 
XMIOM4_L_0 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_2587 
+ BWEB[0] TSMC_2588 D[0] TSMC_2589 TSMC_2590 TSMC_2591 TSMC_2592 Q[0] 
+ TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 
+ TSMC_2599 TSMC_2600 TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_1 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_265 TSMC_266 TSMC_267 
+ TSMC_268 TSMC_2587 BWEB[1] TSMC_2588 D[1] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[1] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 TSMC_2596 
+ TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_2 TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_273 TSMC_274 TSMC_275 
+ TSMC_276 TSMC_2587 BWEB[2] TSMC_2588 D[2] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[2] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 TSMC_2596 
+ TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_3 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_281 TSMC_282 TSMC_283 
+ TSMC_284 TSMC_2587 BWEB[3] TSMC_2588 D[3] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[3] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 TSMC_2596 
+ TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_4 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_289 TSMC_290 TSMC_291 
+ TSMC_292 TSMC_2587 BWEB[4] TSMC_2588 D[4] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[4] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 TSMC_2596 
+ TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_5 TSMC_301 TSMC_302 TSMC_303 TSMC_304 TSMC_297 TSMC_298 TSMC_299 
+ TSMC_300 TSMC_2587 BWEB[5] TSMC_2588 D[5] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[5] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 TSMC_2596 
+ TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_6 TSMC_309 TSMC_310 TSMC_311 TSMC_312 TSMC_305 TSMC_306 TSMC_307 
+ TSMC_308 TSMC_2587 BWEB[6] TSMC_2588 D[6] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[6] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 TSMC_2596 
+ TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_7 TSMC_317 TSMC_318 TSMC_319 TSMC_320 TSMC_313 TSMC_314 TSMC_315 
+ TSMC_316 TSMC_2587 BWEB[7] TSMC_2588 D[7] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[7] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 TSMC_2596 
+ TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_8 TSMC_325 TSMC_326 TSMC_327 TSMC_328 TSMC_321 TSMC_322 TSMC_323 
+ TSMC_324 TSMC_2587 BWEB[8] TSMC_2588 D[8] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[8] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 TSMC_2596 
+ TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_9 TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_329 TSMC_330 TSMC_331 
+ TSMC_332 TSMC_2587 BWEB[9] TSMC_2588 D[9] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[9] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 TSMC_2596 
+ TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_10 TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_337 TSMC_338 TSMC_339 
+ TSMC_340 TSMC_2587 BWEB[10] TSMC_2588 D[10] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[10] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_11 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_345 TSMC_346 TSMC_347 
+ TSMC_348 TSMC_2587 BWEB[11] TSMC_2588 D[11] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[11] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_12 TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_353 TSMC_354 TSMC_355 
+ TSMC_356 TSMC_2587 BWEB[12] TSMC_2588 D[12] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[12] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_13 TSMC_365 TSMC_366 TSMC_367 TSMC_368 TSMC_361 TSMC_362 TSMC_363 
+ TSMC_364 TSMC_2587 BWEB[13] TSMC_2588 D[13] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[13] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_14 TSMC_373 TSMC_374 TSMC_375 TSMC_376 TSMC_369 TSMC_370 TSMC_371 
+ TSMC_372 TSMC_2587 BWEB[14] TSMC_2588 D[14] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[14] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_15 TSMC_381 TSMC_382 TSMC_383 TSMC_384 TSMC_377 TSMC_378 TSMC_379 
+ TSMC_380 TSMC_2587 BWEB[15] TSMC_2588 D[15] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[15] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_16 TSMC_389 TSMC_390 TSMC_391 TSMC_392 TSMC_385 TSMC_386 TSMC_387 
+ TSMC_388 TSMC_2587 BWEB[16] TSMC_2588 D[16] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[16] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_17 TSMC_397 TSMC_398 TSMC_399 TSMC_400 TSMC_393 TSMC_394 TSMC_395 
+ TSMC_396 TSMC_2587 BWEB[17] TSMC_2588 D[17] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[17] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_18 TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_401 TSMC_402 TSMC_403 
+ TSMC_404 TSMC_2587 BWEB[18] TSMC_2588 D[18] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[18] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_19 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_2587 BWEB[19] TSMC_2588 D[19] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[19] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_20 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_417 TSMC_418 TSMC_419 
+ TSMC_420 TSMC_2587 BWEB[20] TSMC_2588 D[20] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[20] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_21 TSMC_429 TSMC_430 TSMC_431 TSMC_432 TSMC_425 TSMC_426 TSMC_427 
+ TSMC_428 TSMC_2587 BWEB[21] TSMC_2588 D[21] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[21] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_22 TSMC_437 TSMC_438 TSMC_439 TSMC_440 TSMC_433 TSMC_434 TSMC_435 
+ TSMC_436 TSMC_2587 BWEB[22] TSMC_2588 D[22] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[22] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_23 TSMC_445 TSMC_446 TSMC_447 TSMC_448 TSMC_441 TSMC_442 TSMC_443 
+ TSMC_444 TSMC_2587 BWEB[23] TSMC_2588 D[23] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[23] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_24 TSMC_453 TSMC_454 TSMC_455 TSMC_456 TSMC_449 TSMC_450 TSMC_451 
+ TSMC_452 TSMC_2587 BWEB[24] TSMC_2588 D[24] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[24] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_25 TSMC_461 TSMC_462 TSMC_463 TSMC_464 TSMC_457 TSMC_458 TSMC_459 
+ TSMC_460 TSMC_2587 BWEB[25] TSMC_2588 D[25] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[25] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_26 TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_465 TSMC_466 TSMC_467 
+ TSMC_468 TSMC_2587 BWEB[26] TSMC_2588 D[26] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[26] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_27 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_2587 BWEB[27] TSMC_2588 D[27] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[27] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_28 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_481 TSMC_482 TSMC_483 
+ TSMC_484 TSMC_2587 BWEB[28] TSMC_2588 D[28] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[28] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_29 TSMC_493 TSMC_494 TSMC_495 TSMC_496 TSMC_489 TSMC_490 TSMC_491 
+ TSMC_492 TSMC_2587 BWEB[29] TSMC_2588 D[29] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[29] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_30 TSMC_501 TSMC_502 TSMC_503 TSMC_504 TSMC_497 TSMC_498 TSMC_499 
+ TSMC_500 TSMC_2587 BWEB[30] TSMC_2588 D[30] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[30] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_31 TSMC_509 TSMC_510 TSMC_511 TSMC_512 TSMC_505 TSMC_506 TSMC_507 
+ TSMC_508 TSMC_2587 BWEB[31] TSMC_2588 D[31] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[31] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_32 TSMC_517 TSMC_518 TSMC_519 TSMC_520 TSMC_513 TSMC_514 TSMC_515 
+ TSMC_516 TSMC_2587 BWEB[32] TSMC_2588 D[32] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[32] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_33 TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_521 TSMC_522 TSMC_523 
+ TSMC_524 TSMC_2587 BWEB[33] TSMC_2588 D[33] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[33] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_34 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_2587 BWEB[34] TSMC_2588 D[34] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[34] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_35 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_537 TSMC_538 TSMC_539 
+ TSMC_540 TSMC_2587 BWEB[35] TSMC_2588 D[35] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[35] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_36 TSMC_549 TSMC_550 TSMC_551 TSMC_552 TSMC_545 TSMC_546 TSMC_547 
+ TSMC_548 TSMC_2587 BWEB[36] TSMC_2588 D[36] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[36] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_37 TSMC_557 TSMC_558 TSMC_559 TSMC_560 TSMC_553 TSMC_554 TSMC_555 
+ TSMC_556 TSMC_2587 BWEB[37] TSMC_2588 D[37] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[37] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_38 TSMC_565 TSMC_566 TSMC_567 TSMC_568 TSMC_561 TSMC_562 TSMC_563 
+ TSMC_564 TSMC_2587 BWEB[38] TSMC_2588 D[38] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[38] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_39 TSMC_573 TSMC_574 TSMC_575 TSMC_576 TSMC_569 TSMC_570 TSMC_571 
+ TSMC_572 TSMC_2587 BWEB[39] TSMC_2588 D[39] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[39] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_40 TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_577 TSMC_578 TSMC_579 
+ TSMC_580 TSMC_2587 BWEB[40] TSMC_2588 D[40] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[40] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_41 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_2587 BWEB[41] TSMC_2588 D[41] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[41] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_42 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_593 TSMC_594 TSMC_595 
+ TSMC_596 TSMC_2587 BWEB[42] TSMC_2588 D[42] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[42] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_43 TSMC_605 TSMC_606 TSMC_607 TSMC_608 TSMC_601 TSMC_602 TSMC_603 
+ TSMC_604 TSMC_2587 BWEB[43] TSMC_2588 D[43] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[43] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_44 TSMC_613 TSMC_614 TSMC_615 TSMC_616 TSMC_609 TSMC_610 TSMC_611 
+ TSMC_612 TSMC_2587 BWEB[44] TSMC_2588 D[44] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[44] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_45 TSMC_621 TSMC_622 TSMC_623 TSMC_624 TSMC_617 TSMC_618 TSMC_619 
+ TSMC_620 TSMC_2587 BWEB[45] TSMC_2588 D[45] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[45] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_46 TSMC_629 TSMC_630 TSMC_631 TSMC_632 TSMC_625 TSMC_626 TSMC_627 
+ TSMC_628 TSMC_2587 BWEB[46] TSMC_2588 D[46] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[46] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_47 TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_633 TSMC_634 TSMC_635 
+ TSMC_636 TSMC_2587 BWEB[47] TSMC_2588 D[47] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[47] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_48 TSMC_645 TSMC_646 TSMC_647 TSMC_648 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_2587 BWEB[48] TSMC_2588 D[48] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[48] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_49 TSMC_653 TSMC_654 TSMC_655 TSMC_656 TSMC_649 TSMC_650 TSMC_651 
+ TSMC_652 TSMC_2587 BWEB[49] TSMC_2588 D[49] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[49] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_50 TSMC_661 TSMC_662 TSMC_663 TSMC_664 TSMC_657 TSMC_658 TSMC_659 
+ TSMC_660 TSMC_2587 BWEB[50] TSMC_2588 D[50] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[50] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_51 TSMC_669 TSMC_670 TSMC_671 TSMC_672 TSMC_665 TSMC_666 TSMC_667 
+ TSMC_668 TSMC_2587 BWEB[51] TSMC_2588 D[51] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[51] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_52 TSMC_677 TSMC_678 TSMC_679 TSMC_680 TSMC_673 TSMC_674 TSMC_675 
+ TSMC_676 TSMC_2587 BWEB[52] TSMC_2588 D[52] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[52] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_53 TSMC_685 TSMC_686 TSMC_687 TSMC_688 TSMC_681 TSMC_682 TSMC_683 
+ TSMC_684 TSMC_2587 BWEB[53] TSMC_2588 D[53] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[53] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_54 TSMC_693 TSMC_694 TSMC_695 TSMC_696 TSMC_689 TSMC_690 TSMC_691 
+ TSMC_692 TSMC_2587 BWEB[54] TSMC_2588 D[54] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[54] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_55 TSMC_701 TSMC_702 TSMC_703 TSMC_704 TSMC_697 TSMC_698 TSMC_699 
+ TSMC_700 TSMC_2587 BWEB[55] TSMC_2588 D[55] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[55] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_56 TSMC_709 TSMC_710 TSMC_711 TSMC_712 TSMC_705 TSMC_706 TSMC_707 
+ TSMC_708 TSMC_2587 BWEB[56] TSMC_2588 D[56] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[56] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_57 TSMC_717 TSMC_718 TSMC_719 TSMC_720 TSMC_713 TSMC_714 TSMC_715 
+ TSMC_716 TSMC_2587 BWEB[57] TSMC_2588 D[57] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[57] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_58 TSMC_725 TSMC_726 TSMC_727 TSMC_728 TSMC_721 TSMC_722 TSMC_723 
+ TSMC_724 TSMC_2587 BWEB[58] TSMC_2588 D[58] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[58] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_59 TSMC_733 TSMC_734 TSMC_735 TSMC_736 TSMC_729 TSMC_730 TSMC_731 
+ TSMC_732 TSMC_2587 BWEB[59] TSMC_2588 D[59] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[59] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_60 TSMC_741 TSMC_742 TSMC_743 TSMC_744 TSMC_737 TSMC_738 TSMC_739 
+ TSMC_740 TSMC_2587 BWEB[60] TSMC_2588 D[60] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[60] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_61 TSMC_749 TSMC_750 TSMC_751 TSMC_752 TSMC_745 TSMC_746 TSMC_747 
+ TSMC_748 TSMC_2587 BWEB[61] TSMC_2588 D[61] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[61] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_62 TSMC_757 TSMC_758 TSMC_759 TSMC_760 TSMC_753 TSMC_754 TSMC_755 
+ TSMC_756 TSMC_2587 BWEB[62] TSMC_2588 D[62] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[62] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_63 TSMC_765 TSMC_766 TSMC_767 TSMC_768 TSMC_761 TSMC_762 TSMC_763 
+ TSMC_764 TSMC_2587 BWEB[63] TSMC_2588 D[63] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[63] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_64 TSMC_773 TSMC_774 TSMC_775 TSMC_776 TSMC_769 TSMC_770 TSMC_771 
+ TSMC_772 TSMC_2587 BWEB[64] TSMC_2588 D[64] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[64] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_65 TSMC_781 TSMC_782 TSMC_783 TSMC_784 TSMC_777 TSMC_778 TSMC_779 
+ TSMC_780 TSMC_2587 BWEB[65] TSMC_2588 D[65] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[65] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_66 TSMC_789 TSMC_790 TSMC_791 TSMC_792 TSMC_785 TSMC_786 TSMC_787 
+ TSMC_788 TSMC_2587 BWEB[66] TSMC_2588 D[66] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[66] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_67 TSMC_797 TSMC_798 TSMC_799 TSMC_800 TSMC_793 TSMC_794 TSMC_795 
+ TSMC_796 TSMC_2587 BWEB[67] TSMC_2588 D[67] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[67] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_68 TSMC_805 TSMC_806 TSMC_807 TSMC_808 TSMC_801 TSMC_802 TSMC_803 
+ TSMC_804 TSMC_2587 BWEB[68] TSMC_2588 D[68] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[68] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_69 TSMC_813 TSMC_814 TSMC_815 TSMC_816 TSMC_809 TSMC_810 TSMC_811 
+ TSMC_812 TSMC_2587 BWEB[69] TSMC_2588 D[69] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[69] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_70 TSMC_821 TSMC_822 TSMC_823 TSMC_824 TSMC_817 TSMC_818 TSMC_819 
+ TSMC_820 TSMC_2587 BWEB[70] TSMC_2588 D[70] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[70] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_L_71 TSMC_829 TSMC_830 TSMC_831 TSMC_832 TSMC_825 TSMC_826 TSMC_827 
+ TSMC_828 TSMC_2587 BWEB[71] TSMC_2588 D[71] TSMC_2589 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[71] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_72 TSMC_837 TSMC_838 TSMC_839 TSMC_840 TSMC_833 TSMC_834 TSMC_835 
+ TSMC_836 TSMC_2602 BWEB[72] TSMC_2603 D[72] TSMC_2604 TSMC_2590 
+ TSMC_2591 TSMC_2592 Q[72] TSMC_2593 VDD VSS TSMC_2594 TSMC_2595 
+ TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 TSMC_2601 
+ S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_73 TSMC_1101 TSMC_1102 TSMC_1103 TSMC_1104 TSMC_1097 TSMC_1098 
+ TSMC_1099 TSMC_1100 TSMC_2602 BWEB[73] TSMC_2603 D[73] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[73] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_74 TSMC_1109 TSMC_1110 TSMC_1111 TSMC_1112 TSMC_1105 TSMC_1106 
+ TSMC_1107 TSMC_1108 TSMC_2602 BWEB[74] TSMC_2603 D[74] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[74] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_75 TSMC_1117 TSMC_1118 TSMC_1119 TSMC_1120 TSMC_1113 TSMC_1114 
+ TSMC_1115 TSMC_1116 TSMC_2602 BWEB[75] TSMC_2603 D[75] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[75] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_76 TSMC_1125 TSMC_1126 TSMC_1127 TSMC_1128 TSMC_1121 TSMC_1122 
+ TSMC_1123 TSMC_1124 TSMC_2602 BWEB[76] TSMC_2603 D[76] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[76] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_77 TSMC_1133 TSMC_1134 TSMC_1135 TSMC_1136 TSMC_1129 TSMC_1130 
+ TSMC_1131 TSMC_1132 TSMC_2602 BWEB[77] TSMC_2603 D[77] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[77] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_78 TSMC_1141 TSMC_1142 TSMC_1143 TSMC_1144 TSMC_1137 TSMC_1138 
+ TSMC_1139 TSMC_1140 TSMC_2602 BWEB[78] TSMC_2603 D[78] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[78] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_79 TSMC_1149 TSMC_1150 TSMC_1151 TSMC_1152 TSMC_1145 TSMC_1146 
+ TSMC_1147 TSMC_1148 TSMC_2602 BWEB[79] TSMC_2603 D[79] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[79] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_80 TSMC_1157 TSMC_1158 TSMC_1159 TSMC_1160 TSMC_1153 TSMC_1154 
+ TSMC_1155 TSMC_1156 TSMC_2602 BWEB[80] TSMC_2603 D[80] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[80] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_81 TSMC_1165 TSMC_1166 TSMC_1167 TSMC_1168 TSMC_1161 TSMC_1162 
+ TSMC_1163 TSMC_1164 TSMC_2602 BWEB[81] TSMC_2603 D[81] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[81] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_82 TSMC_1173 TSMC_1174 TSMC_1175 TSMC_1176 TSMC_1169 TSMC_1170 
+ TSMC_1171 TSMC_1172 TSMC_2602 BWEB[82] TSMC_2603 D[82] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[82] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_83 TSMC_1181 TSMC_1182 TSMC_1183 TSMC_1184 TSMC_1177 TSMC_1178 
+ TSMC_1179 TSMC_1180 TSMC_2602 BWEB[83] TSMC_2603 D[83] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[83] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_84 TSMC_1189 TSMC_1190 TSMC_1191 TSMC_1192 TSMC_1185 TSMC_1186 
+ TSMC_1187 TSMC_1188 TSMC_2602 BWEB[84] TSMC_2603 D[84] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[84] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_85 TSMC_1197 TSMC_1198 TSMC_1199 TSMC_1200 TSMC_1193 TSMC_1194 
+ TSMC_1195 TSMC_1196 TSMC_2602 BWEB[85] TSMC_2603 D[85] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[85] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_86 TSMC_1205 TSMC_1206 TSMC_1207 TSMC_1208 TSMC_1201 TSMC_1202 
+ TSMC_1203 TSMC_1204 TSMC_2602 BWEB[86] TSMC_2603 D[86] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[86] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_87 TSMC_1213 TSMC_1214 TSMC_1215 TSMC_1216 TSMC_1209 TSMC_1210 
+ TSMC_1211 TSMC_1212 TSMC_2602 BWEB[87] TSMC_2603 D[87] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[87] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_88 TSMC_1221 TSMC_1222 TSMC_1223 TSMC_1224 TSMC_1217 TSMC_1218 
+ TSMC_1219 TSMC_1220 TSMC_2602 BWEB[88] TSMC_2603 D[88] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[88] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_89 TSMC_1229 TSMC_1230 TSMC_1231 TSMC_1232 TSMC_1225 TSMC_1226 
+ TSMC_1227 TSMC_1228 TSMC_2602 BWEB[89] TSMC_2603 D[89] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[89] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_90 TSMC_1237 TSMC_1238 TSMC_1239 TSMC_1240 TSMC_1233 TSMC_1234 
+ TSMC_1235 TSMC_1236 TSMC_2602 BWEB[90] TSMC_2603 D[90] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[90] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_91 TSMC_1245 TSMC_1246 TSMC_1247 TSMC_1248 TSMC_1241 TSMC_1242 
+ TSMC_1243 TSMC_1244 TSMC_2602 BWEB[91] TSMC_2603 D[91] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[91] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_92 TSMC_1253 TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1249 TSMC_1250 
+ TSMC_1251 TSMC_1252 TSMC_2602 BWEB[92] TSMC_2603 D[92] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[92] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_93 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1257 TSMC_1258 
+ TSMC_1259 TSMC_1260 TSMC_2602 BWEB[93] TSMC_2603 D[93] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[93] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_94 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_2602 BWEB[94] TSMC_2603 D[94] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[94] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_95 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1273 TSMC_1274 
+ TSMC_1275 TSMC_1276 TSMC_2602 BWEB[95] TSMC_2603 D[95] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[95] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_96 TSMC_1285 TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1281 TSMC_1282 
+ TSMC_1283 TSMC_1284 TSMC_2602 BWEB[96] TSMC_2603 D[96] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[96] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_97 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1289 TSMC_1290 
+ TSMC_1291 TSMC_1292 TSMC_2602 BWEB[97] TSMC_2603 D[97] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[97] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_98 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_2602 BWEB[98] TSMC_2603 D[98] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[98] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_99 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 TSMC_1305 TSMC_1306 
+ TSMC_1307 TSMC_1308 TSMC_2602 BWEB[99] TSMC_2603 D[99] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[99] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_100 TSMC_1317 TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1313 TSMC_1314 
+ TSMC_1315 TSMC_1316 TSMC_2602 BWEB[100] TSMC_2603 D[100] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[100] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_101 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1321 TSMC_1322 
+ TSMC_1323 TSMC_1324 TSMC_2602 BWEB[101] TSMC_2603 D[101] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[101] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_102 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_2602 BWEB[102] TSMC_2603 D[102] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[102] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_103 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 TSMC_1337 TSMC_1338 
+ TSMC_1339 TSMC_1340 TSMC_2602 BWEB[103] TSMC_2603 D[103] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[103] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_104 TSMC_1349 TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1345 TSMC_1346 
+ TSMC_1347 TSMC_1348 TSMC_2602 BWEB[104] TSMC_2603 D[104] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[104] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_105 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1353 TSMC_1354 
+ TSMC_1355 TSMC_1356 TSMC_2602 BWEB[105] TSMC_2603 D[105] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[105] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_106 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_2602 BWEB[106] TSMC_2603 D[106] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[106] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_107 TSMC_1373 TSMC_1374 TSMC_1375 TSMC_1376 TSMC_1369 TSMC_1370 
+ TSMC_1371 TSMC_1372 TSMC_2602 BWEB[107] TSMC_2603 D[107] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[107] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_108 TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1377 TSMC_1378 
+ TSMC_1379 TSMC_1380 TSMC_2602 BWEB[108] TSMC_2603 D[108] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[108] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_109 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1385 TSMC_1386 
+ TSMC_1387 TSMC_1388 TSMC_2602 BWEB[109] TSMC_2603 D[109] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[109] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_110 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_2602 BWEB[110] TSMC_2603 D[110] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[110] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_111 TSMC_1405 TSMC_1406 TSMC_1407 TSMC_1408 TSMC_1401 TSMC_1402 
+ TSMC_1403 TSMC_1404 TSMC_2602 BWEB[111] TSMC_2603 D[111] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[111] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_112 TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1409 TSMC_1410 
+ TSMC_1411 TSMC_1412 TSMC_2602 BWEB[112] TSMC_2603 D[112] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[112] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_113 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_2602 BWEB[113] TSMC_2603 D[113] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[113] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_114 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_2602 BWEB[114] TSMC_2603 D[114] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[114] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_115 TSMC_1437 TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1433 TSMC_1434 
+ TSMC_1435 TSMC_1436 TSMC_2602 BWEB[115] TSMC_2603 D[115] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[115] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_116 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1441 TSMC_1442 
+ TSMC_1443 TSMC_1444 TSMC_2602 BWEB[116] TSMC_2603 D[116] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[116] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_117 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_2602 BWEB[117] TSMC_2603 D[117] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[117] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_118 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 TSMC_1457 TSMC_1458 
+ TSMC_1459 TSMC_1460 TSMC_2602 BWEB[118] TSMC_2603 D[118] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[118] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_119 TSMC_1469 TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1465 TSMC_1466 
+ TSMC_1467 TSMC_1468 TSMC_2602 BWEB[119] TSMC_2603 D[119] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[119] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_120 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1473 TSMC_1474 
+ TSMC_1475 TSMC_1476 TSMC_2602 BWEB[120] TSMC_2603 D[120] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[120] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_121 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_2602 BWEB[121] TSMC_2603 D[121] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[121] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_122 TSMC_1493 TSMC_1494 TSMC_1495 TSMC_1496 TSMC_1489 TSMC_1490 
+ TSMC_1491 TSMC_1492 TSMC_2602 BWEB[122] TSMC_2603 D[122] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[122] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_123 TSMC_1501 TSMC_1502 TSMC_1503 TSMC_1504 TSMC_1497 TSMC_1498 
+ TSMC_1499 TSMC_1500 TSMC_2602 BWEB[123] TSMC_2603 D[123] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[123] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_124 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1505 TSMC_1506 
+ TSMC_1507 TSMC_1508 TSMC_2602 BWEB[124] TSMC_2603 D[124] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[124] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_125 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_2602 BWEB[125] TSMC_2603 D[125] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[125] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_126 TSMC_1525 TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1521 TSMC_1522 
+ TSMC_1523 TSMC_1524 TSMC_2602 BWEB[126] TSMC_2603 D[126] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[126] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_127 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1529 TSMC_1530 
+ TSMC_1531 TSMC_1532 TSMC_2602 BWEB[127] TSMC_2603 D[127] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[127] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_128 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_2602 BWEB[128] TSMC_2603 D[128] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[128] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_129 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 TSMC_1545 TSMC_1546 
+ TSMC_1547 TSMC_1548 TSMC_2602 BWEB[129] TSMC_2603 D[129] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[129] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_130 TSMC_1557 TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1553 TSMC_1554 
+ TSMC_1555 TSMC_1556 TSMC_2602 BWEB[130] TSMC_2603 D[130] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[130] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_131 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1561 TSMC_1562 
+ TSMC_1563 TSMC_1564 TSMC_2602 BWEB[131] TSMC_2603 D[131] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[131] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_132 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_2602 BWEB[132] TSMC_2603 D[132] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[132] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_133 TSMC_1581 TSMC_1582 TSMC_1583 TSMC_1584 TSMC_1577 TSMC_1578 
+ TSMC_1579 TSMC_1580 TSMC_2602 BWEB[133] TSMC_2603 D[133] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[133] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_134 TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1585 TSMC_1586 
+ TSMC_1587 TSMC_1588 TSMC_2602 BWEB[134] TSMC_2603 D[134] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[134] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_135 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_2602 BWEB[135] TSMC_2603 D[135] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[135] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_136 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_2602 BWEB[136] TSMC_2603 D[136] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[136] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_137 TSMC_1613 TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1609 TSMC_1610 
+ TSMC_1611 TSMC_1612 TSMC_2602 BWEB[137] TSMC_2603 D[137] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[137] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_138 TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1617 TSMC_1618 
+ TSMC_1619 TSMC_1620 TSMC_2602 BWEB[138] TSMC_2603 D[138] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[138] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_139 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_2602 BWEB[139] TSMC_2603 D[139] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[139] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_140 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 TSMC_1633 TSMC_1634 
+ TSMC_1635 TSMC_1636 TSMC_2602 BWEB[140] TSMC_2603 D[140] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[140] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_141 TSMC_1645 TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1641 TSMC_1642 
+ TSMC_1643 TSMC_1644 TSMC_2602 BWEB[141] TSMC_2603 D[141] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[141] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_142 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1649 TSMC_1650 
+ TSMC_1651 TSMC_1652 TSMC_2602 BWEB[142] TSMC_2603 D[142] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[142] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIOM4_R_143 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1657 TSMC_1658 
+ TSMC_1659 TSMC_1660 TSMC_2602 BWEB[143] TSMC_2603 D[143] TSMC_2604 
+ TSMC_2590 TSMC_2591 TSMC_2592 Q[143] TSMC_2593 VDD VSS TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 S1CSLVTSW400W90_MIO_SB 
XMIO_SB_EDGE_L VDD TSMC_2605 TSMC_2606 VSS 
+ S1CSLVTSW400W90_MIO_SB_EDGE 
XMIO_SB_EDGE_R VDD TSMC_2605 TSMC_2606 VSS 
+ S1CSLVTSW400W90_MIO_SB_EDGE 
XCNT_M4_SB TSMC_2587 TSMC_2602 TSMC_2586 CEB TSMC_2588 TSMC_2603 CLK TSMC_1667 
+ TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1686 TSMC_1687 TSMC_1688 
+ TSMC_1689 TSMC_1675 TSMC_1708 TSMC_1737 TSMC_1766 TSMC_1795 
+ TSMC_1824 TSMC_1853 TSMC_1882 TSMC_1665 TSMC_1907 TSMC_2133 
+ TSMC_2359 TSMC_2607 TSMC_2608 TSMC_2609 TSMC_2610 TSMC_2594 
+ TSMC_2595 TSMC_2596 TSMC_2597 TSMC_2598 TSMC_2599 TSMC_2600 
+ TSMC_2601 TSMC_2589 TSMC_2604 TSMC_2590 TSMC_2591 TSMC_2592 
+ TSMC_2606 TSMC_2606 TSMC_2606 TSMC_2606 TSMC_2606 RTSEL[0] RTSEL[1] TSMC_2593 
+ TSMC_2606 TSMC_2585 VDD VSS TSMC_2605 WEB WTSEL[0] WTSEL[1] 
+ TSMC_2606 A[2] A[3] A[4] A[5] A[6] A[7] A[8] A[9] A[0] A[1] TSMC_2606 
+ TSMC_2606 S1CSLVTSW400W90_CNT_M4_SB 
XD_WEB WEB TSMC_2606 VSS S1CSLVTSW400W90_DIODE 
XD_CEB CEB TSMC_2606 VSS S1CSLVTSW400W90_DIODE 
XD_CLK CLK TSMC_2606 VSS S1CSLVTSW400W90_DIODE 
XD_A0 A[0] TSMC_2606 VSS S1CSLVTSW400W90_DIODE 
XD_A1 A[1] TSMC_2606 VSS S1CSLVTSW400W90_DIODE 
XD_A2 A[2] TSMC_2606 VSS S1CSLVTSW400W90_DIODE 
XD_A3 A[3] TSMC_2606 VSS S1CSLVTSW400W90_DIODE 
XD_A4 A[4] TSMC_2606 VSS S1CSLVTSW400W90_DIODE 
XD_A5 A[5] TSMC_2606 VSS S1CSLVTSW400W90_DIODE 
XD_A6 A[6] TSMC_2606 VSS S1CSLVTSW400W90_DIODE 
XD_A7 A[7] TSMC_2606 VSS S1CSLVTSW400W90_DIODE 
XD_A8 A[8] TSMC_2606 VSS S1CSLVTSW400W90_DIODE 
XD_A9 A[9] TSMC_2606 VSS S1CSLVTSW400W90_DIODE 
XD_D0 D[0] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D1 D[1] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D2 D[2] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D3 D[3] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D4 D[4] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D5 D[5] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D6 D[6] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D7 D[7] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D8 D[8] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D9 D[9] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D10 D[10] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D11 D[11] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D12 D[12] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D13 D[13] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D14 D[14] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D15 D[15] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D16 D[16] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D17 D[17] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D18 D[18] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D19 D[19] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D20 D[20] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D21 D[21] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D22 D[22] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D23 D[23] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D24 D[24] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D25 D[25] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D26 D[26] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D27 D[27] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D28 D[28] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D29 D[29] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D30 D[30] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D31 D[31] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D32 D[32] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D33 D[33] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D34 D[34] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D35 D[35] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D36 D[36] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D37 D[37] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D38 D[38] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D39 D[39] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D40 D[40] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D41 D[41] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D42 D[42] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D43 D[43] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D44 D[44] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D45 D[45] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D46 D[46] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D47 D[47] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D48 D[48] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D49 D[49] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D50 D[50] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D51 D[51] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D52 D[52] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D53 D[53] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D54 D[54] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D55 D[55] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D56 D[56] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D57 D[57] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D58 D[58] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D59 D[59] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D60 D[60] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D61 D[61] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D62 D[62] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D63 D[63] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D64 D[64] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D65 D[65] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D66 D[66] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D67 D[67] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D68 D[68] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D69 D[69] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D70 D[70] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D71 D[71] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D72 D[72] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D73 D[73] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D74 D[74] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D75 D[75] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D76 D[76] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D77 D[77] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D78 D[78] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D79 D[79] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D80 D[80] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D81 D[81] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D82 D[82] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D83 D[83] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D84 D[84] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D85 D[85] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D86 D[86] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D87 D[87] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D88 D[88] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D89 D[89] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D90 D[90] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D91 D[91] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D92 D[92] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D93 D[93] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D94 D[94] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D95 D[95] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D96 D[96] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D97 D[97] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D98 D[98] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D99 D[99] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D100 D[100] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D101 D[101] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D102 D[102] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D103 D[103] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D104 D[104] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D105 D[105] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D106 D[106] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D107 D[107] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D108 D[108] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D109 D[109] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D110 D[110] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D111 D[111] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D112 D[112] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D113 D[113] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D114 D[114] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D115 D[115] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D116 D[116] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D117 D[117] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D118 D[118] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D119 D[119] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D120 D[120] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D121 D[121] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D122 D[122] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D123 D[123] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D124 D[124] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D125 D[125] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D126 D[126] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D127 D[127] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D128 D[128] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D129 D[129] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D130 D[130] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D131 D[131] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D132 D[132] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D133 D[133] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D134 D[134] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D135 D[135] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D136 D[136] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D137 D[137] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D138 D[138] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D139 D[139] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D140 D[140] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D141 D[141] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D142 D[142] VSS S1CSLVTSW400W90_DIO_TALL 
XD_D143 D[143] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB0 BWEB[0] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB1 BWEB[1] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB2 BWEB[2] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB3 BWEB[3] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB4 BWEB[4] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB5 BWEB[5] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB6 BWEB[6] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB7 BWEB[7] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB8 BWEB[8] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB9 BWEB[9] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB10 BWEB[10] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB11 BWEB[11] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB12 BWEB[12] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB13 BWEB[13] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB14 BWEB[14] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB15 BWEB[15] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB16 BWEB[16] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB17 BWEB[17] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB18 BWEB[18] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB19 BWEB[19] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB20 BWEB[20] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB21 BWEB[21] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB22 BWEB[22] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB23 BWEB[23] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB24 BWEB[24] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB25 BWEB[25] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB26 BWEB[26] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB27 BWEB[27] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB28 BWEB[28] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB29 BWEB[29] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB30 BWEB[30] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB31 BWEB[31] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB32 BWEB[32] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB33 BWEB[33] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB34 BWEB[34] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB35 BWEB[35] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB36 BWEB[36] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB37 BWEB[37] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB38 BWEB[38] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB39 BWEB[39] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB40 BWEB[40] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB41 BWEB[41] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB42 BWEB[42] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB43 BWEB[43] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB44 BWEB[44] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB45 BWEB[45] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB46 BWEB[46] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB47 BWEB[47] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB48 BWEB[48] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB49 BWEB[49] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB50 BWEB[50] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB51 BWEB[51] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB52 BWEB[52] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB53 BWEB[53] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB54 BWEB[54] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB55 BWEB[55] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB56 BWEB[56] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB57 BWEB[57] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB58 BWEB[58] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB59 BWEB[59] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB60 BWEB[60] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB61 BWEB[61] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB62 BWEB[62] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB63 BWEB[63] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB64 BWEB[64] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB65 BWEB[65] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB66 BWEB[66] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB67 BWEB[67] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB68 BWEB[68] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB69 BWEB[69] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB70 BWEB[70] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB71 BWEB[71] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB72 BWEB[72] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB73 BWEB[73] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB74 BWEB[74] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB75 BWEB[75] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB76 BWEB[76] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB77 BWEB[77] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB78 BWEB[78] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB79 BWEB[79] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB80 BWEB[80] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB81 BWEB[81] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB82 BWEB[82] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB83 BWEB[83] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB84 BWEB[84] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB85 BWEB[85] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB86 BWEB[86] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB87 BWEB[87] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB88 BWEB[88] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB89 BWEB[89] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB90 BWEB[90] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB91 BWEB[91] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB92 BWEB[92] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB93 BWEB[93] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB94 BWEB[94] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB95 BWEB[95] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB96 BWEB[96] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB97 BWEB[97] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB98 BWEB[98] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB99 BWEB[99] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB100 BWEB[100] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB101 BWEB[101] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB102 BWEB[102] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB103 BWEB[103] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB104 BWEB[104] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB105 BWEB[105] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB106 BWEB[106] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB107 BWEB[107] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB108 BWEB[108] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB109 BWEB[109] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB110 BWEB[110] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB111 BWEB[111] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB112 BWEB[112] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB113 BWEB[113] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB114 BWEB[114] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB115 BWEB[115] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB116 BWEB[116] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB117 BWEB[117] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB118 BWEB[118] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB119 BWEB[119] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB120 BWEB[120] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB121 BWEB[121] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB122 BWEB[122] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB123 BWEB[123] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB124 BWEB[124] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB125 BWEB[125] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB126 BWEB[126] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB127 BWEB[127] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB128 BWEB[128] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB129 BWEB[129] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB130 BWEB[130] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB131 BWEB[131] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB132 BWEB[132] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB133 BWEB[133] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB134 BWEB[134] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB135 BWEB[135] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB136 BWEB[136] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB137 BWEB[137] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB138 BWEB[138] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB139 BWEB[139] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB140 BWEB[140] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB141 BWEB[141] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB142 BWEB[142] VSS S1CSLVTSW400W90_DIO_TALL 
XD_BWEB143 BWEB[143] VSS S1CSLVTSW400W90_DIO_TALL 
XD_WTESL_1 WTSEL[1] TSMC_2606 VSS S1CSLVTSW400W90_DIODE 
XD_WTESL_0 WTSEL[0] TSMC_2606 VSS S1CSLVTSW400W90_DIODE 
XD_RTESL_1 RTSEL[1] TSMC_2606 VSS S1CSLVTSW400W90_DIODE 
XD_RTESL_0 RTSEL[0] TSMC_2606 VSS S1CSLVTSW400W90_DIODE 
.ENDS


