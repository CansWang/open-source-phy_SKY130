magic
tech sky130A
magscale 1 2
timestamp 1619862920
<< checkpaint >>
rect -1717 -1250 3163 3819
<< nwell >>
rect 0 1318 1889 2559
<< pwell >>
rect 11 982 1893 1172
rect -269 520 1893 982
rect -269 330 1049 520
rect 11 120 1049 330
rect 12 96 1049 120
rect 1323 120 1893 520
rect 1323 96 1888 120
rect 12 10 1888 96
<< mvnmos >>
rect -190 356 -90 956
rect 90 146 190 1146
rect 246 146 346 1146
rect 402 146 502 1146
rect 558 146 658 1146
rect 714 146 814 1146
rect 870 146 970 1146
rect 1136 546 1236 1146
rect 1402 146 1502 1146
rect 1558 146 1658 1146
rect 1714 146 1814 1146
<< mvpmos >>
rect 248 1552 348 2152
rect 404 1552 504 2152
rect 780 1384 880 2384
rect 1046 1384 1146 2384
rect 1202 1384 1302 2384
rect 1358 1384 1458 2384
rect 1514 1384 1614 2384
rect 1670 1384 1770 2384
<< mvndiff >>
rect 37 1076 90 1146
rect 37 1042 45 1076
rect 79 1042 90 1076
rect 37 1008 90 1042
rect 37 974 45 1008
rect 79 974 90 1008
rect -243 878 -190 956
rect -243 844 -235 878
rect -201 844 -190 878
rect -243 810 -190 844
rect -243 776 -235 810
rect -201 776 -190 810
rect -243 742 -190 776
rect -243 708 -235 742
rect -201 708 -190 742
rect -243 674 -190 708
rect -243 640 -235 674
rect -201 640 -190 674
rect -243 606 -190 640
rect -243 572 -235 606
rect -201 572 -190 606
rect -243 538 -190 572
rect -243 504 -235 538
rect -201 504 -190 538
rect -243 470 -190 504
rect -243 436 -235 470
rect -201 436 -190 470
rect -243 402 -190 436
rect -243 368 -235 402
rect -201 368 -190 402
rect -243 356 -190 368
rect -90 878 -37 956
rect -90 844 -79 878
rect -45 844 -37 878
rect -90 810 -37 844
rect -90 776 -79 810
rect -45 776 -37 810
rect -90 742 -37 776
rect -90 708 -79 742
rect -45 708 -37 742
rect -90 674 -37 708
rect -90 640 -79 674
rect -45 640 -37 674
rect -90 606 -37 640
rect -90 572 -79 606
rect -45 572 -37 606
rect -90 538 -37 572
rect -90 504 -79 538
rect -45 504 -37 538
rect -90 470 -37 504
rect -90 436 -79 470
rect -45 436 -37 470
rect -90 402 -37 436
rect -90 368 -79 402
rect -45 368 -37 402
rect -90 356 -37 368
rect 37 940 90 974
rect 37 906 45 940
rect 79 906 90 940
rect 37 872 90 906
rect 37 838 45 872
rect 79 838 90 872
rect 37 804 90 838
rect 37 770 45 804
rect 79 770 90 804
rect 37 736 90 770
rect 37 702 45 736
rect 79 702 90 736
rect 37 668 90 702
rect 37 634 45 668
rect 79 634 90 668
rect 37 600 90 634
rect 37 566 45 600
rect 79 566 90 600
rect 37 532 90 566
rect 37 498 45 532
rect 79 498 90 532
rect 37 464 90 498
rect 37 430 45 464
rect 79 430 90 464
rect 37 396 90 430
rect 37 362 45 396
rect 79 362 90 396
rect 37 328 90 362
rect 37 294 45 328
rect 79 294 90 328
rect 37 260 90 294
rect 37 226 45 260
rect 79 226 90 260
rect 37 192 90 226
rect 37 158 45 192
rect 79 158 90 192
rect 37 146 90 158
rect 190 1076 246 1146
rect 190 1042 201 1076
rect 235 1042 246 1076
rect 190 1008 246 1042
rect 190 974 201 1008
rect 235 974 246 1008
rect 190 940 246 974
rect 190 906 201 940
rect 235 906 246 940
rect 190 872 246 906
rect 190 838 201 872
rect 235 838 246 872
rect 190 804 246 838
rect 190 770 201 804
rect 235 770 246 804
rect 190 736 246 770
rect 190 702 201 736
rect 235 702 246 736
rect 190 668 246 702
rect 190 634 201 668
rect 235 634 246 668
rect 190 600 246 634
rect 190 566 201 600
rect 235 566 246 600
rect 190 532 246 566
rect 190 498 201 532
rect 235 498 246 532
rect 190 464 246 498
rect 190 430 201 464
rect 235 430 246 464
rect 190 396 246 430
rect 190 362 201 396
rect 235 362 246 396
rect 190 328 246 362
rect 190 294 201 328
rect 235 294 246 328
rect 190 260 246 294
rect 190 226 201 260
rect 235 226 246 260
rect 190 192 246 226
rect 190 158 201 192
rect 235 158 246 192
rect 190 146 246 158
rect 346 1076 402 1146
rect 346 1042 357 1076
rect 391 1042 402 1076
rect 346 1008 402 1042
rect 346 974 357 1008
rect 391 974 402 1008
rect 346 940 402 974
rect 346 906 357 940
rect 391 906 402 940
rect 346 872 402 906
rect 346 838 357 872
rect 391 838 402 872
rect 346 804 402 838
rect 346 770 357 804
rect 391 770 402 804
rect 346 736 402 770
rect 346 702 357 736
rect 391 702 402 736
rect 346 668 402 702
rect 346 634 357 668
rect 391 634 402 668
rect 346 600 402 634
rect 346 566 357 600
rect 391 566 402 600
rect 346 532 402 566
rect 346 498 357 532
rect 391 498 402 532
rect 346 464 402 498
rect 346 430 357 464
rect 391 430 402 464
rect 346 396 402 430
rect 346 362 357 396
rect 391 362 402 396
rect 346 328 402 362
rect 346 294 357 328
rect 391 294 402 328
rect 346 260 402 294
rect 346 226 357 260
rect 391 226 402 260
rect 346 192 402 226
rect 346 158 357 192
rect 391 158 402 192
rect 346 146 402 158
rect 502 1076 558 1146
rect 502 1042 513 1076
rect 547 1042 558 1076
rect 502 1008 558 1042
rect 502 974 513 1008
rect 547 974 558 1008
rect 502 940 558 974
rect 502 906 513 940
rect 547 906 558 940
rect 502 872 558 906
rect 502 838 513 872
rect 547 838 558 872
rect 502 804 558 838
rect 502 770 513 804
rect 547 770 558 804
rect 502 736 558 770
rect 502 702 513 736
rect 547 702 558 736
rect 502 668 558 702
rect 502 634 513 668
rect 547 634 558 668
rect 502 600 558 634
rect 502 566 513 600
rect 547 566 558 600
rect 502 532 558 566
rect 502 498 513 532
rect 547 498 558 532
rect 502 464 558 498
rect 502 430 513 464
rect 547 430 558 464
rect 502 396 558 430
rect 502 362 513 396
rect 547 362 558 396
rect 502 328 558 362
rect 502 294 513 328
rect 547 294 558 328
rect 502 260 558 294
rect 502 226 513 260
rect 547 226 558 260
rect 502 192 558 226
rect 502 158 513 192
rect 547 158 558 192
rect 502 146 558 158
rect 658 1076 714 1146
rect 658 1042 669 1076
rect 703 1042 714 1076
rect 658 1008 714 1042
rect 658 974 669 1008
rect 703 974 714 1008
rect 658 940 714 974
rect 658 906 669 940
rect 703 906 714 940
rect 658 872 714 906
rect 658 838 669 872
rect 703 838 714 872
rect 658 804 714 838
rect 658 770 669 804
rect 703 770 714 804
rect 658 736 714 770
rect 658 702 669 736
rect 703 702 714 736
rect 658 668 714 702
rect 658 634 669 668
rect 703 634 714 668
rect 658 600 714 634
rect 658 566 669 600
rect 703 566 714 600
rect 658 532 714 566
rect 658 498 669 532
rect 703 498 714 532
rect 658 464 714 498
rect 658 430 669 464
rect 703 430 714 464
rect 658 396 714 430
rect 658 362 669 396
rect 703 362 714 396
rect 658 328 714 362
rect 658 294 669 328
rect 703 294 714 328
rect 658 260 714 294
rect 658 226 669 260
rect 703 226 714 260
rect 658 192 714 226
rect 658 158 669 192
rect 703 158 714 192
rect 658 146 714 158
rect 814 1076 870 1146
rect 814 1042 825 1076
rect 859 1042 870 1076
rect 814 1008 870 1042
rect 814 974 825 1008
rect 859 974 870 1008
rect 814 940 870 974
rect 814 906 825 940
rect 859 906 870 940
rect 814 872 870 906
rect 814 838 825 872
rect 859 838 870 872
rect 814 804 870 838
rect 814 770 825 804
rect 859 770 870 804
rect 814 736 870 770
rect 814 702 825 736
rect 859 702 870 736
rect 814 668 870 702
rect 814 634 825 668
rect 859 634 870 668
rect 814 600 870 634
rect 814 566 825 600
rect 859 566 870 600
rect 814 532 870 566
rect 814 498 825 532
rect 859 498 870 532
rect 814 464 870 498
rect 814 430 825 464
rect 859 430 870 464
rect 814 396 870 430
rect 814 362 825 396
rect 859 362 870 396
rect 814 328 870 362
rect 814 294 825 328
rect 859 294 870 328
rect 814 260 870 294
rect 814 226 825 260
rect 859 226 870 260
rect 814 192 870 226
rect 814 158 825 192
rect 859 158 870 192
rect 814 146 870 158
rect 970 1076 1023 1146
rect 970 1042 981 1076
rect 1015 1042 1023 1076
rect 970 1008 1023 1042
rect 970 974 981 1008
rect 1015 974 1023 1008
rect 970 940 1023 974
rect 970 906 981 940
rect 1015 906 1023 940
rect 970 872 1023 906
rect 970 838 981 872
rect 1015 838 1023 872
rect 970 804 1023 838
rect 970 770 981 804
rect 1015 770 1023 804
rect 970 736 1023 770
rect 970 702 981 736
rect 1015 702 1023 736
rect 970 668 1023 702
rect 970 634 981 668
rect 1015 634 1023 668
rect 970 600 1023 634
rect 970 566 981 600
rect 1015 566 1023 600
rect 970 532 1023 566
rect 1083 1068 1136 1146
rect 1083 1034 1091 1068
rect 1125 1034 1136 1068
rect 1083 1000 1136 1034
rect 1083 966 1091 1000
rect 1125 966 1136 1000
rect 1083 932 1136 966
rect 1083 898 1091 932
rect 1125 898 1136 932
rect 1083 864 1136 898
rect 1083 830 1091 864
rect 1125 830 1136 864
rect 1083 796 1136 830
rect 1083 762 1091 796
rect 1125 762 1136 796
rect 1083 728 1136 762
rect 1083 694 1091 728
rect 1125 694 1136 728
rect 1083 660 1136 694
rect 1083 626 1091 660
rect 1125 626 1136 660
rect 1083 592 1136 626
rect 1083 558 1091 592
rect 1125 558 1136 592
rect 1083 546 1136 558
rect 1236 1068 1289 1146
rect 1236 1034 1247 1068
rect 1281 1034 1289 1068
rect 1236 1000 1289 1034
rect 1236 966 1247 1000
rect 1281 966 1289 1000
rect 1236 932 1289 966
rect 1236 898 1247 932
rect 1281 898 1289 932
rect 1236 864 1289 898
rect 1236 830 1247 864
rect 1281 830 1289 864
rect 1236 796 1289 830
rect 1236 762 1247 796
rect 1281 762 1289 796
rect 1236 728 1289 762
rect 1236 694 1247 728
rect 1281 694 1289 728
rect 1236 660 1289 694
rect 1236 626 1247 660
rect 1281 626 1289 660
rect 1236 592 1289 626
rect 1236 558 1247 592
rect 1281 558 1289 592
rect 1236 546 1289 558
rect 1349 1076 1402 1146
rect 1349 1042 1357 1076
rect 1391 1042 1402 1076
rect 1349 1008 1402 1042
rect 1349 974 1357 1008
rect 1391 974 1402 1008
rect 1349 940 1402 974
rect 1349 906 1357 940
rect 1391 906 1402 940
rect 1349 872 1402 906
rect 1349 838 1357 872
rect 1391 838 1402 872
rect 1349 804 1402 838
rect 1349 770 1357 804
rect 1391 770 1402 804
rect 1349 736 1402 770
rect 1349 702 1357 736
rect 1391 702 1402 736
rect 1349 668 1402 702
rect 1349 634 1357 668
rect 1391 634 1402 668
rect 1349 600 1402 634
rect 1349 566 1357 600
rect 1391 566 1402 600
rect 970 498 981 532
rect 1015 498 1023 532
rect 1349 532 1402 566
rect 970 464 1023 498
rect 970 430 981 464
rect 1015 430 1023 464
rect 970 396 1023 430
rect 970 362 981 396
rect 1015 362 1023 396
rect 970 328 1023 362
rect 970 294 981 328
rect 1015 294 1023 328
rect 970 260 1023 294
rect 970 226 981 260
rect 1015 226 1023 260
rect 970 192 1023 226
rect 970 158 981 192
rect 1015 158 1023 192
rect 970 146 1023 158
rect 1349 498 1357 532
rect 1391 498 1402 532
rect 1349 464 1402 498
rect 1349 430 1357 464
rect 1391 430 1402 464
rect 1349 396 1402 430
rect 1349 362 1357 396
rect 1391 362 1402 396
rect 1349 328 1402 362
rect 1349 294 1357 328
rect 1391 294 1402 328
rect 1349 260 1402 294
rect 1349 226 1357 260
rect 1391 226 1402 260
rect 1349 192 1402 226
rect 1349 158 1357 192
rect 1391 158 1402 192
rect 1349 146 1402 158
rect 1502 1076 1558 1146
rect 1502 1042 1513 1076
rect 1547 1042 1558 1076
rect 1502 1008 1558 1042
rect 1502 974 1513 1008
rect 1547 974 1558 1008
rect 1502 940 1558 974
rect 1502 906 1513 940
rect 1547 906 1558 940
rect 1502 872 1558 906
rect 1502 838 1513 872
rect 1547 838 1558 872
rect 1502 804 1558 838
rect 1502 770 1513 804
rect 1547 770 1558 804
rect 1502 736 1558 770
rect 1502 702 1513 736
rect 1547 702 1558 736
rect 1502 668 1558 702
rect 1502 634 1513 668
rect 1547 634 1558 668
rect 1502 600 1558 634
rect 1502 566 1513 600
rect 1547 566 1558 600
rect 1502 532 1558 566
rect 1502 498 1513 532
rect 1547 498 1558 532
rect 1502 464 1558 498
rect 1502 430 1513 464
rect 1547 430 1558 464
rect 1502 396 1558 430
rect 1502 362 1513 396
rect 1547 362 1558 396
rect 1502 328 1558 362
rect 1502 294 1513 328
rect 1547 294 1558 328
rect 1502 260 1558 294
rect 1502 226 1513 260
rect 1547 226 1558 260
rect 1502 192 1558 226
rect 1502 158 1513 192
rect 1547 158 1558 192
rect 1502 146 1558 158
rect 1658 1076 1714 1146
rect 1658 1042 1669 1076
rect 1703 1042 1714 1076
rect 1658 1008 1714 1042
rect 1658 974 1669 1008
rect 1703 974 1714 1008
rect 1658 940 1714 974
rect 1658 906 1669 940
rect 1703 906 1714 940
rect 1658 872 1714 906
rect 1658 838 1669 872
rect 1703 838 1714 872
rect 1658 804 1714 838
rect 1658 770 1669 804
rect 1703 770 1714 804
rect 1658 736 1714 770
rect 1658 702 1669 736
rect 1703 702 1714 736
rect 1658 668 1714 702
rect 1658 634 1669 668
rect 1703 634 1714 668
rect 1658 600 1714 634
rect 1658 566 1669 600
rect 1703 566 1714 600
rect 1658 532 1714 566
rect 1658 498 1669 532
rect 1703 498 1714 532
rect 1658 464 1714 498
rect 1658 430 1669 464
rect 1703 430 1714 464
rect 1658 396 1714 430
rect 1658 362 1669 396
rect 1703 362 1714 396
rect 1658 328 1714 362
rect 1658 294 1669 328
rect 1703 294 1714 328
rect 1658 260 1714 294
rect 1658 226 1669 260
rect 1703 226 1714 260
rect 1658 192 1714 226
rect 1658 158 1669 192
rect 1703 158 1714 192
rect 1658 146 1714 158
rect 1814 1076 1867 1146
rect 1814 1042 1825 1076
rect 1859 1042 1867 1076
rect 1814 1008 1867 1042
rect 1814 974 1825 1008
rect 1859 974 1867 1008
rect 1814 940 1867 974
rect 1814 906 1825 940
rect 1859 906 1867 940
rect 1814 872 1867 906
rect 1814 838 1825 872
rect 1859 838 1867 872
rect 1814 804 1867 838
rect 1814 770 1825 804
rect 1859 770 1867 804
rect 1814 736 1867 770
rect 1814 702 1825 736
rect 1859 702 1867 736
rect 1814 668 1867 702
rect 1814 634 1825 668
rect 1859 634 1867 668
rect 1814 600 1867 634
rect 1814 566 1825 600
rect 1859 566 1867 600
rect 1814 532 1867 566
rect 1814 498 1825 532
rect 1859 498 1867 532
rect 1814 464 1867 498
rect 1814 430 1825 464
rect 1859 430 1867 464
rect 1814 396 1867 430
rect 1814 362 1825 396
rect 1859 362 1867 396
rect 1814 328 1867 362
rect 1814 294 1825 328
rect 1859 294 1867 328
rect 1814 260 1867 294
rect 1814 226 1825 260
rect 1859 226 1867 260
rect 1814 192 1867 226
rect 1814 158 1825 192
rect 1859 158 1867 192
rect 1814 146 1867 158
<< mvpdiff >>
rect 727 2314 780 2384
rect 727 2280 735 2314
rect 769 2280 780 2314
rect 727 2246 780 2280
rect 727 2212 735 2246
rect 769 2212 780 2246
rect 727 2178 780 2212
rect 195 2074 248 2152
rect 195 2040 203 2074
rect 237 2040 248 2074
rect 195 2006 248 2040
rect 195 1972 203 2006
rect 237 1972 248 2006
rect 195 1938 248 1972
rect 195 1904 203 1938
rect 237 1904 248 1938
rect 195 1870 248 1904
rect 195 1836 203 1870
rect 237 1836 248 1870
rect 195 1802 248 1836
rect 195 1768 203 1802
rect 237 1768 248 1802
rect 195 1734 248 1768
rect 195 1700 203 1734
rect 237 1700 248 1734
rect 195 1666 248 1700
rect 195 1632 203 1666
rect 237 1632 248 1666
rect 195 1598 248 1632
rect 195 1564 203 1598
rect 237 1564 248 1598
rect 195 1552 248 1564
rect 348 2074 404 2152
rect 348 2040 359 2074
rect 393 2040 404 2074
rect 348 2006 404 2040
rect 348 1972 359 2006
rect 393 1972 404 2006
rect 348 1938 404 1972
rect 348 1904 359 1938
rect 393 1904 404 1938
rect 348 1870 404 1904
rect 348 1836 359 1870
rect 393 1836 404 1870
rect 348 1802 404 1836
rect 348 1768 359 1802
rect 393 1768 404 1802
rect 348 1734 404 1768
rect 348 1700 359 1734
rect 393 1700 404 1734
rect 348 1666 404 1700
rect 348 1632 359 1666
rect 393 1632 404 1666
rect 348 1598 404 1632
rect 348 1564 359 1598
rect 393 1564 404 1598
rect 348 1552 404 1564
rect 504 2074 557 2152
rect 504 2040 515 2074
rect 549 2040 557 2074
rect 504 2006 557 2040
rect 504 1972 515 2006
rect 549 1972 557 2006
rect 504 1938 557 1972
rect 504 1904 515 1938
rect 549 1904 557 1938
rect 504 1870 557 1904
rect 504 1836 515 1870
rect 549 1836 557 1870
rect 504 1802 557 1836
rect 504 1768 515 1802
rect 549 1768 557 1802
rect 504 1734 557 1768
rect 504 1700 515 1734
rect 549 1700 557 1734
rect 504 1666 557 1700
rect 504 1632 515 1666
rect 549 1632 557 1666
rect 504 1598 557 1632
rect 504 1564 515 1598
rect 549 1564 557 1598
rect 504 1552 557 1564
rect 727 2144 735 2178
rect 769 2144 780 2178
rect 727 2110 780 2144
rect 727 2076 735 2110
rect 769 2076 780 2110
rect 727 2042 780 2076
rect 727 2008 735 2042
rect 769 2008 780 2042
rect 727 1974 780 2008
rect 727 1940 735 1974
rect 769 1940 780 1974
rect 727 1906 780 1940
rect 727 1872 735 1906
rect 769 1872 780 1906
rect 727 1838 780 1872
rect 727 1804 735 1838
rect 769 1804 780 1838
rect 727 1770 780 1804
rect 727 1736 735 1770
rect 769 1736 780 1770
rect 727 1702 780 1736
rect 727 1668 735 1702
rect 769 1668 780 1702
rect 727 1634 780 1668
rect 727 1600 735 1634
rect 769 1600 780 1634
rect 727 1566 780 1600
rect 727 1532 735 1566
rect 769 1532 780 1566
rect 727 1498 780 1532
rect 727 1464 735 1498
rect 769 1464 780 1498
rect 727 1430 780 1464
rect 727 1396 735 1430
rect 769 1396 780 1430
rect 727 1384 780 1396
rect 880 2314 933 2384
rect 880 2280 891 2314
rect 925 2280 933 2314
rect 880 2246 933 2280
rect 880 2212 891 2246
rect 925 2212 933 2246
rect 880 2178 933 2212
rect 880 2144 891 2178
rect 925 2144 933 2178
rect 880 2110 933 2144
rect 880 2076 891 2110
rect 925 2076 933 2110
rect 880 2042 933 2076
rect 880 2008 891 2042
rect 925 2008 933 2042
rect 880 1974 933 2008
rect 880 1940 891 1974
rect 925 1940 933 1974
rect 880 1906 933 1940
rect 880 1872 891 1906
rect 925 1872 933 1906
rect 880 1838 933 1872
rect 880 1804 891 1838
rect 925 1804 933 1838
rect 880 1770 933 1804
rect 880 1736 891 1770
rect 925 1736 933 1770
rect 880 1702 933 1736
rect 880 1668 891 1702
rect 925 1668 933 1702
rect 880 1634 933 1668
rect 880 1600 891 1634
rect 925 1600 933 1634
rect 880 1566 933 1600
rect 880 1532 891 1566
rect 925 1532 933 1566
rect 880 1498 933 1532
rect 880 1464 891 1498
rect 925 1464 933 1498
rect 880 1430 933 1464
rect 880 1396 891 1430
rect 925 1396 933 1430
rect 880 1384 933 1396
rect 993 2314 1046 2384
rect 993 2280 1001 2314
rect 1035 2280 1046 2314
rect 993 2246 1046 2280
rect 993 2212 1001 2246
rect 1035 2212 1046 2246
rect 993 2178 1046 2212
rect 993 2144 1001 2178
rect 1035 2144 1046 2178
rect 993 2110 1046 2144
rect 993 2076 1001 2110
rect 1035 2076 1046 2110
rect 993 2042 1046 2076
rect 993 2008 1001 2042
rect 1035 2008 1046 2042
rect 993 1974 1046 2008
rect 993 1940 1001 1974
rect 1035 1940 1046 1974
rect 993 1906 1046 1940
rect 993 1872 1001 1906
rect 1035 1872 1046 1906
rect 993 1838 1046 1872
rect 993 1804 1001 1838
rect 1035 1804 1046 1838
rect 993 1770 1046 1804
rect 993 1736 1001 1770
rect 1035 1736 1046 1770
rect 993 1702 1046 1736
rect 993 1668 1001 1702
rect 1035 1668 1046 1702
rect 993 1634 1046 1668
rect 993 1600 1001 1634
rect 1035 1600 1046 1634
rect 993 1566 1046 1600
rect 993 1532 1001 1566
rect 1035 1532 1046 1566
rect 993 1498 1046 1532
rect 993 1464 1001 1498
rect 1035 1464 1046 1498
rect 993 1430 1046 1464
rect 993 1396 1001 1430
rect 1035 1396 1046 1430
rect 993 1384 1046 1396
rect 1146 2314 1202 2384
rect 1146 2280 1157 2314
rect 1191 2280 1202 2314
rect 1146 2246 1202 2280
rect 1146 2212 1157 2246
rect 1191 2212 1202 2246
rect 1146 2178 1202 2212
rect 1146 2144 1157 2178
rect 1191 2144 1202 2178
rect 1146 2110 1202 2144
rect 1146 2076 1157 2110
rect 1191 2076 1202 2110
rect 1146 2042 1202 2076
rect 1146 2008 1157 2042
rect 1191 2008 1202 2042
rect 1146 1974 1202 2008
rect 1146 1940 1157 1974
rect 1191 1940 1202 1974
rect 1146 1906 1202 1940
rect 1146 1872 1157 1906
rect 1191 1872 1202 1906
rect 1146 1838 1202 1872
rect 1146 1804 1157 1838
rect 1191 1804 1202 1838
rect 1146 1770 1202 1804
rect 1146 1736 1157 1770
rect 1191 1736 1202 1770
rect 1146 1702 1202 1736
rect 1146 1668 1157 1702
rect 1191 1668 1202 1702
rect 1146 1634 1202 1668
rect 1146 1600 1157 1634
rect 1191 1600 1202 1634
rect 1146 1566 1202 1600
rect 1146 1532 1157 1566
rect 1191 1532 1202 1566
rect 1146 1498 1202 1532
rect 1146 1464 1157 1498
rect 1191 1464 1202 1498
rect 1146 1430 1202 1464
rect 1146 1396 1157 1430
rect 1191 1396 1202 1430
rect 1146 1384 1202 1396
rect 1302 2314 1358 2384
rect 1302 2280 1313 2314
rect 1347 2280 1358 2314
rect 1302 2246 1358 2280
rect 1302 2212 1313 2246
rect 1347 2212 1358 2246
rect 1302 2178 1358 2212
rect 1302 2144 1313 2178
rect 1347 2144 1358 2178
rect 1302 2110 1358 2144
rect 1302 2076 1313 2110
rect 1347 2076 1358 2110
rect 1302 2042 1358 2076
rect 1302 2008 1313 2042
rect 1347 2008 1358 2042
rect 1302 1974 1358 2008
rect 1302 1940 1313 1974
rect 1347 1940 1358 1974
rect 1302 1906 1358 1940
rect 1302 1872 1313 1906
rect 1347 1872 1358 1906
rect 1302 1838 1358 1872
rect 1302 1804 1313 1838
rect 1347 1804 1358 1838
rect 1302 1770 1358 1804
rect 1302 1736 1313 1770
rect 1347 1736 1358 1770
rect 1302 1702 1358 1736
rect 1302 1668 1313 1702
rect 1347 1668 1358 1702
rect 1302 1634 1358 1668
rect 1302 1600 1313 1634
rect 1347 1600 1358 1634
rect 1302 1566 1358 1600
rect 1302 1532 1313 1566
rect 1347 1532 1358 1566
rect 1302 1498 1358 1532
rect 1302 1464 1313 1498
rect 1347 1464 1358 1498
rect 1302 1430 1358 1464
rect 1302 1396 1313 1430
rect 1347 1396 1358 1430
rect 1302 1384 1358 1396
rect 1458 2314 1514 2384
rect 1458 2280 1469 2314
rect 1503 2280 1514 2314
rect 1458 2246 1514 2280
rect 1458 2212 1469 2246
rect 1503 2212 1514 2246
rect 1458 2178 1514 2212
rect 1458 2144 1469 2178
rect 1503 2144 1514 2178
rect 1458 2110 1514 2144
rect 1458 2076 1469 2110
rect 1503 2076 1514 2110
rect 1458 2042 1514 2076
rect 1458 2008 1469 2042
rect 1503 2008 1514 2042
rect 1458 1974 1514 2008
rect 1458 1940 1469 1974
rect 1503 1940 1514 1974
rect 1458 1906 1514 1940
rect 1458 1872 1469 1906
rect 1503 1872 1514 1906
rect 1458 1838 1514 1872
rect 1458 1804 1469 1838
rect 1503 1804 1514 1838
rect 1458 1770 1514 1804
rect 1458 1736 1469 1770
rect 1503 1736 1514 1770
rect 1458 1702 1514 1736
rect 1458 1668 1469 1702
rect 1503 1668 1514 1702
rect 1458 1634 1514 1668
rect 1458 1600 1469 1634
rect 1503 1600 1514 1634
rect 1458 1566 1514 1600
rect 1458 1532 1469 1566
rect 1503 1532 1514 1566
rect 1458 1498 1514 1532
rect 1458 1464 1469 1498
rect 1503 1464 1514 1498
rect 1458 1430 1514 1464
rect 1458 1396 1469 1430
rect 1503 1396 1514 1430
rect 1458 1384 1514 1396
rect 1614 2314 1670 2384
rect 1614 2280 1625 2314
rect 1659 2280 1670 2314
rect 1614 2246 1670 2280
rect 1614 2212 1625 2246
rect 1659 2212 1670 2246
rect 1614 2178 1670 2212
rect 1614 2144 1625 2178
rect 1659 2144 1670 2178
rect 1614 2110 1670 2144
rect 1614 2076 1625 2110
rect 1659 2076 1670 2110
rect 1614 2042 1670 2076
rect 1614 2008 1625 2042
rect 1659 2008 1670 2042
rect 1614 1974 1670 2008
rect 1614 1940 1625 1974
rect 1659 1940 1670 1974
rect 1614 1906 1670 1940
rect 1614 1872 1625 1906
rect 1659 1872 1670 1906
rect 1614 1838 1670 1872
rect 1614 1804 1625 1838
rect 1659 1804 1670 1838
rect 1614 1770 1670 1804
rect 1614 1736 1625 1770
rect 1659 1736 1670 1770
rect 1614 1702 1670 1736
rect 1614 1668 1625 1702
rect 1659 1668 1670 1702
rect 1614 1634 1670 1668
rect 1614 1600 1625 1634
rect 1659 1600 1670 1634
rect 1614 1566 1670 1600
rect 1614 1532 1625 1566
rect 1659 1532 1670 1566
rect 1614 1498 1670 1532
rect 1614 1464 1625 1498
rect 1659 1464 1670 1498
rect 1614 1430 1670 1464
rect 1614 1396 1625 1430
rect 1659 1396 1670 1430
rect 1614 1384 1670 1396
rect 1770 2314 1823 2384
rect 1770 2280 1781 2314
rect 1815 2280 1823 2314
rect 1770 2246 1823 2280
rect 1770 2212 1781 2246
rect 1815 2212 1823 2246
rect 1770 2178 1823 2212
rect 1770 2144 1781 2178
rect 1815 2144 1823 2178
rect 1770 2110 1823 2144
rect 1770 2076 1781 2110
rect 1815 2076 1823 2110
rect 1770 2042 1823 2076
rect 1770 2008 1781 2042
rect 1815 2008 1823 2042
rect 1770 1974 1823 2008
rect 1770 1940 1781 1974
rect 1815 1940 1823 1974
rect 1770 1906 1823 1940
rect 1770 1872 1781 1906
rect 1815 1872 1823 1906
rect 1770 1838 1823 1872
rect 1770 1804 1781 1838
rect 1815 1804 1823 1838
rect 1770 1770 1823 1804
rect 1770 1736 1781 1770
rect 1815 1736 1823 1770
rect 1770 1702 1823 1736
rect 1770 1668 1781 1702
rect 1815 1668 1823 1702
rect 1770 1634 1823 1668
rect 1770 1600 1781 1634
rect 1815 1600 1823 1634
rect 1770 1566 1823 1600
rect 1770 1532 1781 1566
rect 1815 1532 1823 1566
rect 1770 1498 1823 1532
rect 1770 1464 1781 1498
rect 1815 1464 1823 1498
rect 1770 1430 1823 1464
rect 1770 1396 1781 1430
rect 1815 1396 1823 1430
rect 1770 1384 1823 1396
<< mvndiffc >>
rect 45 1042 79 1076
rect 45 974 79 1008
rect -235 844 -201 878
rect -235 776 -201 810
rect -235 708 -201 742
rect -235 640 -201 674
rect -235 572 -201 606
rect -235 504 -201 538
rect -235 436 -201 470
rect -235 368 -201 402
rect -79 844 -45 878
rect -79 776 -45 810
rect -79 708 -45 742
rect -79 640 -45 674
rect -79 572 -45 606
rect -79 504 -45 538
rect -79 436 -45 470
rect -79 368 -45 402
rect 45 906 79 940
rect 45 838 79 872
rect 45 770 79 804
rect 45 702 79 736
rect 45 634 79 668
rect 45 566 79 600
rect 45 498 79 532
rect 45 430 79 464
rect 45 362 79 396
rect 45 294 79 328
rect 45 226 79 260
rect 45 158 79 192
rect 201 1042 235 1076
rect 201 974 235 1008
rect 201 906 235 940
rect 201 838 235 872
rect 201 770 235 804
rect 201 702 235 736
rect 201 634 235 668
rect 201 566 235 600
rect 201 498 235 532
rect 201 430 235 464
rect 201 362 235 396
rect 201 294 235 328
rect 201 226 235 260
rect 201 158 235 192
rect 357 1042 391 1076
rect 357 974 391 1008
rect 357 906 391 940
rect 357 838 391 872
rect 357 770 391 804
rect 357 702 391 736
rect 357 634 391 668
rect 357 566 391 600
rect 357 498 391 532
rect 357 430 391 464
rect 357 362 391 396
rect 357 294 391 328
rect 357 226 391 260
rect 357 158 391 192
rect 513 1042 547 1076
rect 513 974 547 1008
rect 513 906 547 940
rect 513 838 547 872
rect 513 770 547 804
rect 513 702 547 736
rect 513 634 547 668
rect 513 566 547 600
rect 513 498 547 532
rect 513 430 547 464
rect 513 362 547 396
rect 513 294 547 328
rect 513 226 547 260
rect 513 158 547 192
rect 669 1042 703 1076
rect 669 974 703 1008
rect 669 906 703 940
rect 669 838 703 872
rect 669 770 703 804
rect 669 702 703 736
rect 669 634 703 668
rect 669 566 703 600
rect 669 498 703 532
rect 669 430 703 464
rect 669 362 703 396
rect 669 294 703 328
rect 669 226 703 260
rect 669 158 703 192
rect 825 1042 859 1076
rect 825 974 859 1008
rect 825 906 859 940
rect 825 838 859 872
rect 825 770 859 804
rect 825 702 859 736
rect 825 634 859 668
rect 825 566 859 600
rect 825 498 859 532
rect 825 430 859 464
rect 825 362 859 396
rect 825 294 859 328
rect 825 226 859 260
rect 825 158 859 192
rect 981 1042 1015 1076
rect 981 974 1015 1008
rect 981 906 1015 940
rect 981 838 1015 872
rect 981 770 1015 804
rect 981 702 1015 736
rect 981 634 1015 668
rect 981 566 1015 600
rect 1091 1034 1125 1068
rect 1091 966 1125 1000
rect 1091 898 1125 932
rect 1091 830 1125 864
rect 1091 762 1125 796
rect 1091 694 1125 728
rect 1091 626 1125 660
rect 1091 558 1125 592
rect 1247 1034 1281 1068
rect 1247 966 1281 1000
rect 1247 898 1281 932
rect 1247 830 1281 864
rect 1247 762 1281 796
rect 1247 694 1281 728
rect 1247 626 1281 660
rect 1247 558 1281 592
rect 1357 1042 1391 1076
rect 1357 974 1391 1008
rect 1357 906 1391 940
rect 1357 838 1391 872
rect 1357 770 1391 804
rect 1357 702 1391 736
rect 1357 634 1391 668
rect 1357 566 1391 600
rect 981 498 1015 532
rect 981 430 1015 464
rect 981 362 1015 396
rect 981 294 1015 328
rect 981 226 1015 260
rect 981 158 1015 192
rect 1357 498 1391 532
rect 1357 430 1391 464
rect 1357 362 1391 396
rect 1357 294 1391 328
rect 1357 226 1391 260
rect 1357 158 1391 192
rect 1513 1042 1547 1076
rect 1513 974 1547 1008
rect 1513 906 1547 940
rect 1513 838 1547 872
rect 1513 770 1547 804
rect 1513 702 1547 736
rect 1513 634 1547 668
rect 1513 566 1547 600
rect 1513 498 1547 532
rect 1513 430 1547 464
rect 1513 362 1547 396
rect 1513 294 1547 328
rect 1513 226 1547 260
rect 1513 158 1547 192
rect 1669 1042 1703 1076
rect 1669 974 1703 1008
rect 1669 906 1703 940
rect 1669 838 1703 872
rect 1669 770 1703 804
rect 1669 702 1703 736
rect 1669 634 1703 668
rect 1669 566 1703 600
rect 1669 498 1703 532
rect 1669 430 1703 464
rect 1669 362 1703 396
rect 1669 294 1703 328
rect 1669 226 1703 260
rect 1669 158 1703 192
rect 1825 1042 1859 1076
rect 1825 974 1859 1008
rect 1825 906 1859 940
rect 1825 838 1859 872
rect 1825 770 1859 804
rect 1825 702 1859 736
rect 1825 634 1859 668
rect 1825 566 1859 600
rect 1825 498 1859 532
rect 1825 430 1859 464
rect 1825 362 1859 396
rect 1825 294 1859 328
rect 1825 226 1859 260
rect 1825 158 1859 192
<< mvpdiffc >>
rect 735 2280 769 2314
rect 735 2212 769 2246
rect 203 2040 237 2074
rect 203 1972 237 2006
rect 203 1904 237 1938
rect 203 1836 237 1870
rect 203 1768 237 1802
rect 203 1700 237 1734
rect 203 1632 237 1666
rect 203 1564 237 1598
rect 359 2040 393 2074
rect 359 1972 393 2006
rect 359 1904 393 1938
rect 359 1836 393 1870
rect 359 1768 393 1802
rect 359 1700 393 1734
rect 359 1632 393 1666
rect 359 1564 393 1598
rect 515 2040 549 2074
rect 515 1972 549 2006
rect 515 1904 549 1938
rect 515 1836 549 1870
rect 515 1768 549 1802
rect 515 1700 549 1734
rect 515 1632 549 1666
rect 515 1564 549 1598
rect 735 2144 769 2178
rect 735 2076 769 2110
rect 735 2008 769 2042
rect 735 1940 769 1974
rect 735 1872 769 1906
rect 735 1804 769 1838
rect 735 1736 769 1770
rect 735 1668 769 1702
rect 735 1600 769 1634
rect 735 1532 769 1566
rect 735 1464 769 1498
rect 735 1396 769 1430
rect 891 2280 925 2314
rect 891 2212 925 2246
rect 891 2144 925 2178
rect 891 2076 925 2110
rect 891 2008 925 2042
rect 891 1940 925 1974
rect 891 1872 925 1906
rect 891 1804 925 1838
rect 891 1736 925 1770
rect 891 1668 925 1702
rect 891 1600 925 1634
rect 891 1532 925 1566
rect 891 1464 925 1498
rect 891 1396 925 1430
rect 1001 2280 1035 2314
rect 1001 2212 1035 2246
rect 1001 2144 1035 2178
rect 1001 2076 1035 2110
rect 1001 2008 1035 2042
rect 1001 1940 1035 1974
rect 1001 1872 1035 1906
rect 1001 1804 1035 1838
rect 1001 1736 1035 1770
rect 1001 1668 1035 1702
rect 1001 1600 1035 1634
rect 1001 1532 1035 1566
rect 1001 1464 1035 1498
rect 1001 1396 1035 1430
rect 1157 2280 1191 2314
rect 1157 2212 1191 2246
rect 1157 2144 1191 2178
rect 1157 2076 1191 2110
rect 1157 2008 1191 2042
rect 1157 1940 1191 1974
rect 1157 1872 1191 1906
rect 1157 1804 1191 1838
rect 1157 1736 1191 1770
rect 1157 1668 1191 1702
rect 1157 1600 1191 1634
rect 1157 1532 1191 1566
rect 1157 1464 1191 1498
rect 1157 1396 1191 1430
rect 1313 2280 1347 2314
rect 1313 2212 1347 2246
rect 1313 2144 1347 2178
rect 1313 2076 1347 2110
rect 1313 2008 1347 2042
rect 1313 1940 1347 1974
rect 1313 1872 1347 1906
rect 1313 1804 1347 1838
rect 1313 1736 1347 1770
rect 1313 1668 1347 1702
rect 1313 1600 1347 1634
rect 1313 1532 1347 1566
rect 1313 1464 1347 1498
rect 1313 1396 1347 1430
rect 1469 2280 1503 2314
rect 1469 2212 1503 2246
rect 1469 2144 1503 2178
rect 1469 2076 1503 2110
rect 1469 2008 1503 2042
rect 1469 1940 1503 1974
rect 1469 1872 1503 1906
rect 1469 1804 1503 1838
rect 1469 1736 1503 1770
rect 1469 1668 1503 1702
rect 1469 1600 1503 1634
rect 1469 1532 1503 1566
rect 1469 1464 1503 1498
rect 1469 1396 1503 1430
rect 1625 2280 1659 2314
rect 1625 2212 1659 2246
rect 1625 2144 1659 2178
rect 1625 2076 1659 2110
rect 1625 2008 1659 2042
rect 1625 1940 1659 1974
rect 1625 1872 1659 1906
rect 1625 1804 1659 1838
rect 1625 1736 1659 1770
rect 1625 1668 1659 1702
rect 1625 1600 1659 1634
rect 1625 1532 1659 1566
rect 1625 1464 1659 1498
rect 1625 1396 1659 1430
rect 1781 2280 1815 2314
rect 1781 2212 1815 2246
rect 1781 2144 1815 2178
rect 1781 2076 1815 2110
rect 1781 2008 1815 2042
rect 1781 1940 1815 1974
rect 1781 1872 1815 1906
rect 1781 1804 1815 1838
rect 1781 1736 1815 1770
rect 1781 1668 1815 1702
rect 1781 1600 1815 1634
rect 1781 1532 1815 1566
rect 1781 1464 1815 1498
rect 1781 1396 1815 1430
<< mvpsubdiff >>
rect 38 36 62 70
rect 96 36 132 70
rect 166 36 202 70
rect 236 36 272 70
rect 306 36 342 70
rect 376 36 412 70
rect 446 36 482 70
rect 516 36 552 70
rect 586 36 622 70
rect 656 36 692 70
rect 726 36 762 70
rect 796 36 832 70
rect 866 36 902 70
rect 936 36 972 70
rect 1006 36 1042 70
rect 1076 36 1112 70
rect 1146 36 1182 70
rect 1216 36 1252 70
rect 1286 36 1321 70
rect 1355 36 1390 70
rect 1424 36 1459 70
rect 1493 36 1528 70
rect 1562 36 1597 70
rect 1631 36 1666 70
rect 1700 36 1735 70
rect 1769 36 1804 70
rect 1838 36 1862 70
<< mvnsubdiff >>
rect 67 2458 121 2492
rect 155 2458 189 2492
rect 223 2458 257 2492
rect 291 2458 325 2492
rect 359 2458 393 2492
rect 427 2458 461 2492
rect 495 2458 529 2492
rect 563 2458 597 2492
rect 631 2458 665 2492
rect 699 2458 733 2492
rect 767 2458 801 2492
rect 835 2458 869 2492
rect 903 2458 937 2492
rect 971 2458 1005 2492
rect 1039 2458 1073 2492
rect 1107 2458 1141 2492
rect 1175 2458 1209 2492
rect 1243 2458 1277 2492
rect 1311 2458 1345 2492
rect 1379 2458 1413 2492
rect 1447 2458 1481 2492
rect 1515 2458 1549 2492
rect 1583 2458 1617 2492
rect 1651 2458 1685 2492
rect 1719 2458 1753 2492
rect 1787 2458 1821 2492
<< mvpsubdiffcont >>
rect 62 36 96 70
rect 132 36 166 70
rect 202 36 236 70
rect 272 36 306 70
rect 342 36 376 70
rect 412 36 446 70
rect 482 36 516 70
rect 552 36 586 70
rect 622 36 656 70
rect 692 36 726 70
rect 762 36 796 70
rect 832 36 866 70
rect 902 36 936 70
rect 972 36 1006 70
rect 1042 36 1076 70
rect 1112 36 1146 70
rect 1182 36 1216 70
rect 1252 36 1286 70
rect 1321 36 1355 70
rect 1390 36 1424 70
rect 1459 36 1493 70
rect 1528 36 1562 70
rect 1597 36 1631 70
rect 1666 36 1700 70
rect 1735 36 1769 70
rect 1804 36 1838 70
<< mvnsubdiffcont >>
rect 121 2458 155 2492
rect 189 2458 223 2492
rect 257 2458 291 2492
rect 325 2458 359 2492
rect 393 2458 427 2492
rect 461 2458 495 2492
rect 529 2458 563 2492
rect 597 2458 631 2492
rect 665 2458 699 2492
rect 733 2458 767 2492
rect 801 2458 835 2492
rect 869 2458 903 2492
rect 937 2458 971 2492
rect 1005 2458 1039 2492
rect 1073 2458 1107 2492
rect 1141 2458 1175 2492
rect 1209 2458 1243 2492
rect 1277 2458 1311 2492
rect 1345 2458 1379 2492
rect 1413 2458 1447 2492
rect 1481 2458 1515 2492
rect 1549 2458 1583 2492
rect 1617 2458 1651 2492
rect 1685 2458 1719 2492
rect 1753 2458 1787 2492
<< poly >>
rect 780 2384 880 2416
rect 1046 2384 1146 2416
rect 1202 2384 1302 2416
rect 1358 2384 1458 2416
rect 1514 2384 1614 2416
rect 1670 2384 1770 2416
rect 248 2152 348 2184
rect 404 2152 504 2184
rect 248 1520 348 1552
rect 214 1504 348 1520
rect 214 1470 230 1504
rect 264 1470 298 1504
rect 332 1470 348 1504
rect 214 1454 348 1470
rect 404 1520 504 1552
rect 404 1504 538 1520
rect 404 1470 420 1504
rect 454 1470 488 1504
rect 522 1470 538 1504
rect 404 1454 538 1470
rect 780 1352 880 1384
rect 746 1336 880 1352
rect 746 1302 762 1336
rect 796 1302 830 1336
rect 864 1302 880 1336
rect 746 1286 880 1302
rect 1046 1352 1146 1384
rect 1202 1352 1302 1384
rect 1358 1352 1458 1384
rect 1514 1352 1614 1384
rect 1670 1352 1770 1384
rect 1046 1336 1770 1352
rect 1046 1302 1062 1336
rect 1096 1302 1136 1336
rect 1170 1302 1209 1336
rect 1243 1302 1282 1336
rect 1316 1302 1355 1336
rect 1389 1302 1428 1336
rect 1462 1302 1501 1336
rect 1535 1302 1574 1336
rect 1608 1302 1647 1336
rect 1681 1302 1720 1336
rect 1754 1302 1770 1336
rect 1046 1286 1770 1302
rect 90 1228 502 1244
rect 90 1194 106 1228
rect 140 1194 176 1228
rect 210 1194 245 1228
rect 279 1194 314 1228
rect 348 1194 383 1228
rect 417 1194 452 1228
rect 486 1194 502 1228
rect 90 1178 502 1194
rect 90 1146 190 1178
rect 246 1146 346 1178
rect 402 1146 502 1178
rect 558 1228 970 1244
rect 558 1194 574 1228
rect 608 1194 644 1228
rect 678 1194 713 1228
rect 747 1194 782 1228
rect 816 1194 851 1228
rect 885 1194 920 1228
rect 954 1194 970 1228
rect 558 1178 970 1194
rect 1102 1228 1236 1244
rect 1102 1194 1118 1228
rect 1152 1194 1186 1228
rect 1220 1194 1236 1228
rect 1102 1178 1236 1194
rect 558 1146 658 1178
rect 714 1146 814 1178
rect 870 1146 970 1178
rect 1136 1146 1236 1178
rect 1402 1228 1814 1244
rect 1402 1194 1418 1228
rect 1452 1194 1488 1228
rect 1522 1194 1557 1228
rect 1591 1194 1626 1228
rect 1660 1194 1695 1228
rect 1729 1194 1764 1228
rect 1798 1194 1814 1228
rect 1402 1178 1814 1194
rect 1402 1146 1502 1178
rect 1558 1146 1658 1178
rect 1714 1146 1814 1178
rect -224 1038 -90 1054
rect -224 1004 -208 1038
rect -174 1004 -140 1038
rect -106 1004 -90 1038
rect -224 988 -90 1004
rect -190 956 -90 988
rect -190 324 -90 356
rect 1136 514 1236 546
rect 90 114 190 146
rect 246 114 346 146
rect 402 114 502 146
rect 558 114 658 146
rect 714 114 814 146
rect 870 114 970 146
rect 1402 114 1502 146
rect 1558 114 1658 146
rect 1714 114 1814 146
<< polycont >>
rect 230 1470 264 1504
rect 298 1470 332 1504
rect 420 1470 454 1504
rect 488 1470 522 1504
rect 762 1302 796 1336
rect 830 1302 864 1336
rect 1062 1302 1096 1336
rect 1136 1302 1170 1336
rect 1209 1302 1243 1336
rect 1282 1302 1316 1336
rect 1355 1302 1389 1336
rect 1428 1302 1462 1336
rect 1501 1302 1535 1336
rect 1574 1302 1608 1336
rect 1647 1302 1681 1336
rect 1720 1302 1754 1336
rect 106 1194 140 1228
rect 176 1194 210 1228
rect 245 1194 279 1228
rect 314 1194 348 1228
rect 383 1194 417 1228
rect 452 1194 486 1228
rect 574 1194 608 1228
rect 644 1194 678 1228
rect 713 1194 747 1228
rect 782 1194 816 1228
rect 851 1194 885 1228
rect 920 1194 954 1228
rect 1118 1194 1152 1228
rect 1186 1194 1220 1228
rect 1418 1194 1452 1228
rect 1488 1194 1522 1228
rect 1557 1194 1591 1228
rect 1626 1194 1660 1228
rect 1695 1194 1729 1228
rect 1764 1194 1798 1228
rect -208 1004 -174 1038
rect -140 1004 -106 1038
<< locali >>
rect 101 2458 121 2492
rect 176 2458 189 2492
rect 251 2458 257 2492
rect 291 2458 292 2492
rect 359 2458 367 2492
rect 427 2458 442 2492
rect 495 2458 517 2492
rect 563 2458 592 2492
rect 631 2458 665 2492
rect 701 2458 733 2492
rect 776 2458 801 2492
rect 851 2458 869 2492
rect 926 2458 937 2492
rect 1001 2458 1005 2492
rect 1039 2458 1042 2492
rect 1107 2458 1117 2492
rect 1175 2458 1192 2492
rect 1243 2458 1267 2492
rect 1311 2458 1342 2492
rect 1379 2458 1413 2492
rect 1451 2458 1481 2492
rect 1525 2458 1549 2492
rect 1599 2458 1617 2492
rect 1673 2458 1685 2492
rect 1747 2458 1753 2492
rect 735 2314 769 2350
rect 735 2246 769 2278
rect 735 2178 769 2205
rect 735 2110 769 2132
rect 203 2008 237 2040
rect 203 1938 237 1972
rect 203 1870 237 1892
rect 203 1802 237 1810
rect 203 1762 237 1768
rect 203 1680 237 1700
rect 203 1598 237 1632
rect 203 1548 237 1564
rect 359 2008 393 2040
rect 359 1938 393 1972
rect 359 1870 393 1892
rect 359 1802 393 1810
rect 359 1762 393 1768
rect 359 1680 393 1700
rect 359 1598 393 1632
rect 515 2008 549 2040
rect 515 1938 549 1972
rect 515 1870 549 1892
rect 515 1802 549 1810
rect 515 1762 549 1768
rect 515 1680 549 1700
rect 515 1598 549 1632
rect 359 1548 393 1564
rect 436 1521 470 1559
rect 515 1548 549 1564
rect 735 2042 769 2059
rect 735 1974 769 1986
rect 735 1906 769 1913
rect 735 1838 769 1840
rect 735 1801 769 1804
rect 735 1728 769 1736
rect 735 1655 769 1668
rect 735 1582 769 1600
rect 735 1509 769 1532
rect 214 1470 228 1504
rect 264 1470 298 1504
rect 334 1470 348 1504
rect 404 1470 420 1504
rect 470 1487 488 1504
rect 454 1470 488 1487
rect 522 1470 538 1504
rect 735 1430 769 1464
rect 735 1380 769 1396
rect 891 2314 925 2330
rect 891 2257 925 2280
rect 891 2182 925 2212
rect 891 2110 925 2144
rect 891 2042 925 2073
rect 891 1974 925 1998
rect 891 1906 925 1923
rect 891 1838 925 1848
rect 891 1770 925 1773
rect 891 1732 925 1736
rect 891 1657 925 1668
rect 891 1582 925 1600
rect 891 1506 925 1532
rect 891 1430 925 1464
rect 891 1380 925 1396
rect 1001 2314 1035 2330
rect 1001 2246 1035 2280
rect 1001 2178 1035 2211
rect 1001 2110 1035 2137
rect 1001 2042 1035 2063
rect 1001 1974 1035 1989
rect 1001 1906 1035 1915
rect 1001 1838 1035 1841
rect 1001 1801 1035 1804
rect 1001 1727 1035 1736
rect 1001 1653 1035 1668
rect 1001 1579 1035 1600
rect 1001 1505 1035 1532
rect 1001 1430 1035 1464
rect 1001 1380 1035 1396
rect 1157 2314 1191 2350
rect 1157 2246 1191 2276
rect 1157 2178 1191 2202
rect 1157 2110 1191 2128
rect 1157 2042 1191 2054
rect 1157 1974 1191 1980
rect 1157 1866 1191 1872
rect 1157 1792 1191 1804
rect 1157 1718 1191 1736
rect 1157 1644 1191 1668
rect 1157 1570 1191 1600
rect 1157 1498 1191 1532
rect 1157 1430 1191 1464
rect 1157 1380 1191 1396
rect 1313 2314 1347 2330
rect 1313 2246 1347 2280
rect 1313 2178 1347 2211
rect 1313 2110 1347 2137
rect 1313 2042 1347 2063
rect 1313 1974 1347 1989
rect 1313 1906 1347 1915
rect 1313 1838 1347 1841
rect 1313 1801 1347 1804
rect 1313 1727 1347 1736
rect 1313 1653 1347 1668
rect 1313 1579 1347 1600
rect 1313 1505 1347 1532
rect 1313 1430 1347 1464
rect 1313 1380 1347 1396
rect 1469 2314 1503 2350
rect 1469 2246 1503 2276
rect 1469 2178 1503 2202
rect 1469 2110 1503 2128
rect 1469 2042 1503 2054
rect 1469 1974 1503 1980
rect 1469 1866 1503 1872
rect 1469 1792 1503 1804
rect 1469 1718 1503 1736
rect 1469 1644 1503 1668
rect 1469 1570 1503 1600
rect 1469 1498 1503 1532
rect 1469 1430 1503 1464
rect 1469 1380 1503 1396
rect 1625 2314 1659 2330
rect 1625 2246 1659 2280
rect 1625 2178 1659 2211
rect 1625 2110 1659 2137
rect 1625 2042 1659 2063
rect 1625 1974 1659 1989
rect 1625 1906 1659 1915
rect 1625 1838 1659 1841
rect 1625 1801 1659 1804
rect 1625 1727 1659 1736
rect 1625 1653 1659 1668
rect 1625 1579 1659 1600
rect 1625 1505 1659 1532
rect 1625 1430 1659 1464
rect 1625 1380 1659 1396
rect 1781 2314 1815 2350
rect 1781 2246 1815 2276
rect 1781 2178 1815 2202
rect 1781 2110 1815 2128
rect 1781 2042 1815 2054
rect 1781 1974 1815 1980
rect 1781 1866 1815 1872
rect 1781 1792 1815 1804
rect 1781 1718 1815 1736
rect 1781 1644 1815 1668
rect 1781 1570 1815 1600
rect 1781 1498 1815 1532
rect 1781 1430 1815 1464
rect 1781 1380 1815 1396
rect 796 1302 808 1336
rect 864 1302 880 1336
rect 1046 1302 1058 1336
rect 1096 1302 1134 1336
rect 1170 1302 1209 1336
rect 1244 1302 1282 1336
rect 1320 1302 1355 1336
rect 1396 1302 1428 1336
rect 1472 1302 1501 1336
rect 1548 1302 1574 1336
rect 1624 1302 1647 1336
rect 1699 1302 1720 1336
rect 1754 1302 1770 1336
rect 90 1194 102 1228
rect 140 1194 176 1228
rect 221 1194 245 1228
rect 306 1194 314 1228
rect 348 1194 357 1228
rect 417 1194 442 1228
rect 486 1194 502 1228
rect 558 1194 574 1228
rect 608 1194 622 1228
rect 678 1194 703 1228
rect 747 1194 782 1228
rect 818 1194 851 1228
rect 899 1194 920 1228
rect 954 1194 970 1228
rect 1152 1194 1167 1228
rect 1220 1194 1236 1228
rect 1402 1194 1414 1228
rect 1452 1194 1488 1228
rect 1542 1194 1557 1228
rect 1591 1194 1601 1228
rect 1660 1194 1694 1228
rect 1729 1194 1764 1228
rect 1798 1194 1814 1228
rect 45 1076 79 1100
rect -224 1004 -208 1038
rect -174 1004 -140 1038
rect -106 1004 -90 1038
rect 45 1008 79 1025
rect 45 940 79 950
rect -235 882 -201 894
rect -235 810 -201 844
rect -235 742 -201 768
rect -235 674 -201 688
rect -235 606 -201 607
rect -235 560 -201 572
rect -235 479 -201 504
rect -235 402 -201 436
rect -235 352 -201 364
rect -79 882 -45 894
rect -79 810 -45 844
rect -79 742 -45 768
rect -79 674 -45 688
rect -79 606 -45 607
rect -79 560 -45 572
rect -79 479 -45 504
rect -79 402 -45 436
rect -79 352 -45 364
rect 45 872 79 875
rect 45 834 79 838
rect 45 759 79 770
rect 45 684 79 702
rect 45 609 79 634
rect 45 534 79 566
rect 45 464 79 498
rect 45 396 79 425
rect 45 328 79 350
rect 45 260 79 294
rect 45 192 79 226
rect 45 142 79 158
rect 201 1076 235 1092
rect 201 1008 235 1042
rect 201 940 235 964
rect 201 872 235 890
rect 201 804 235 816
rect 201 736 235 742
rect 201 628 235 634
rect 201 554 235 566
rect 201 480 235 498
rect 201 405 235 430
rect 201 330 235 362
rect 201 260 235 294
rect 201 192 235 221
rect 201 142 235 146
rect 357 1076 391 1100
rect 357 1008 391 1025
rect 357 940 391 950
rect 357 872 391 875
rect 357 834 391 838
rect 357 759 391 770
rect 357 684 391 702
rect 357 609 391 634
rect 357 534 391 566
rect 357 464 391 498
rect 357 396 391 425
rect 357 328 391 350
rect 357 260 391 294
rect 357 192 391 226
rect 357 142 391 158
rect 513 1076 547 1092
rect 513 1008 547 1042
rect 513 940 547 964
rect 513 872 547 890
rect 513 804 547 816
rect 513 736 547 742
rect 513 628 547 634
rect 513 554 547 566
rect 513 480 547 498
rect 513 405 547 430
rect 513 330 547 362
rect 513 260 547 294
rect 513 192 547 221
rect 513 142 547 146
rect 669 1076 703 1100
rect 669 1008 703 1025
rect 669 940 703 950
rect 669 872 703 875
rect 669 834 703 838
rect 669 759 703 770
rect 669 684 703 702
rect 669 609 703 634
rect 669 534 703 566
rect 669 464 703 498
rect 669 396 703 425
rect 669 328 703 350
rect 669 260 703 294
rect 669 192 703 226
rect 669 142 703 158
rect 825 1076 859 1092
rect 825 1008 859 1042
rect 825 940 859 964
rect 825 872 859 890
rect 825 804 859 816
rect 825 736 859 742
rect 825 628 859 634
rect 825 554 859 566
rect 825 480 859 498
rect 825 405 859 430
rect 825 330 859 362
rect 825 260 859 294
rect 825 192 859 221
rect 825 142 859 146
rect 981 1076 1015 1100
rect 981 1008 1015 1027
rect 981 940 1015 954
rect 981 872 1015 881
rect 981 804 1015 808
rect 981 769 1015 770
rect 981 696 1015 702
rect 981 623 1015 634
rect 981 550 1015 566
rect 1091 1073 1125 1084
rect 1091 1000 1125 1034
rect 1091 932 1125 959
rect 1091 864 1125 879
rect 1091 796 1125 799
rect 1091 753 1125 762
rect 1091 673 1125 694
rect 1091 592 1125 626
rect 1091 542 1125 558
rect 1247 1068 1281 1093
rect 1247 1000 1281 1017
rect 1247 932 1281 941
rect 1247 864 1281 865
rect 1247 823 1281 830
rect 1247 746 1281 762
rect 1247 669 1281 694
rect 1247 592 1281 626
rect 1247 542 1281 558
rect 1357 1076 1391 1100
rect 1357 1008 1391 1025
rect 1357 940 1391 950
rect 1357 872 1391 875
rect 1357 834 1391 838
rect 1357 759 1391 770
rect 1357 684 1391 702
rect 1357 609 1391 634
rect 981 477 1015 498
rect 981 404 1015 430
rect 981 330 1015 362
rect 981 260 1015 294
rect 981 192 1015 226
rect 981 142 1015 158
rect 1357 534 1391 566
rect 1357 464 1391 498
rect 1357 396 1391 425
rect 1357 328 1391 350
rect 1357 260 1391 294
rect 1357 192 1391 226
rect 1357 142 1391 158
rect 1513 1076 1547 1092
rect 1513 1008 1547 1042
rect 1513 940 1547 946
rect 1513 872 1547 874
rect 1513 836 1547 838
rect 1513 764 1547 770
rect 1513 691 1547 702
rect 1513 618 1547 634
rect 1513 545 1547 566
rect 1513 472 1547 498
rect 1513 399 1547 430
rect 1513 328 1547 362
rect 1513 260 1547 292
rect 1513 192 1547 219
rect 1513 142 1547 146
rect 1669 1076 1703 1100
rect 1669 1008 1703 1025
rect 1669 940 1703 950
rect 1669 872 1703 875
rect 1669 834 1703 838
rect 1669 759 1703 770
rect 1669 684 1703 702
rect 1669 609 1703 634
rect 1669 534 1703 566
rect 1669 464 1703 498
rect 1669 396 1703 425
rect 1669 328 1703 350
rect 1669 260 1703 294
rect 1669 192 1703 226
rect 1669 142 1703 158
rect 1825 1076 1859 1092
rect 1825 1008 1859 1042
rect 1825 940 1859 964
rect 1825 872 1859 890
rect 1825 804 1859 816
rect 1825 736 1859 742
rect 1825 628 1859 634
rect 1825 554 1859 566
rect 1825 480 1859 498
rect 1825 405 1859 430
rect 1825 330 1859 362
rect 1825 260 1859 294
rect 1825 192 1859 221
rect 1825 142 1859 146
rect 96 36 113 70
rect 166 36 188 70
rect 236 36 262 70
rect 306 36 336 70
rect 376 36 410 70
rect 446 36 482 70
rect 518 36 552 70
rect 592 36 622 70
rect 666 36 692 70
rect 740 36 762 70
rect 814 36 832 70
rect 888 36 902 70
rect 962 36 972 70
rect 1036 36 1042 70
rect 1110 36 1112 70
rect 1146 36 1150 70
rect 1216 36 1224 70
rect 1286 36 1298 70
rect 1355 36 1372 70
rect 1424 36 1446 70
rect 1493 36 1520 70
rect 1562 36 1594 70
rect 1631 36 1666 70
rect 1702 36 1735 70
rect 1776 36 1804 70
rect 1850 36 1862 70
<< viali >>
rect 67 2458 101 2492
rect 142 2458 155 2492
rect 155 2458 176 2492
rect 217 2458 223 2492
rect 223 2458 251 2492
rect 292 2458 325 2492
rect 325 2458 326 2492
rect 367 2458 393 2492
rect 393 2458 401 2492
rect 442 2458 461 2492
rect 461 2458 476 2492
rect 517 2458 529 2492
rect 529 2458 551 2492
rect 592 2458 597 2492
rect 597 2458 626 2492
rect 667 2458 699 2492
rect 699 2458 701 2492
rect 742 2458 767 2492
rect 767 2458 776 2492
rect 817 2458 835 2492
rect 835 2458 851 2492
rect 892 2458 903 2492
rect 903 2458 926 2492
rect 967 2458 971 2492
rect 971 2458 1001 2492
rect 1042 2458 1073 2492
rect 1073 2458 1076 2492
rect 1117 2458 1141 2492
rect 1141 2458 1151 2492
rect 1192 2458 1209 2492
rect 1209 2458 1226 2492
rect 1267 2458 1277 2492
rect 1277 2458 1301 2492
rect 1342 2458 1345 2492
rect 1345 2458 1376 2492
rect 1417 2458 1447 2492
rect 1447 2458 1451 2492
rect 1491 2458 1515 2492
rect 1515 2458 1525 2492
rect 1565 2458 1583 2492
rect 1583 2458 1599 2492
rect 1639 2458 1651 2492
rect 1651 2458 1673 2492
rect 1713 2458 1719 2492
rect 1719 2458 1747 2492
rect 1787 2458 1821 2492
rect 735 2350 769 2384
rect 1157 2350 1191 2384
rect 735 2280 769 2312
rect 735 2278 769 2280
rect 735 2212 769 2239
rect 735 2205 769 2212
rect 735 2144 769 2166
rect 735 2132 769 2144
rect 203 2074 237 2090
rect 203 2056 237 2074
rect 203 2006 237 2008
rect 203 1974 237 2006
rect 203 1904 237 1926
rect 203 1892 237 1904
rect 203 1836 237 1844
rect 203 1810 237 1836
rect 203 1734 237 1762
rect 203 1728 237 1734
rect 203 1666 237 1680
rect 203 1646 237 1666
rect 203 1564 237 1598
rect 359 2074 393 2090
rect 359 2056 393 2074
rect 359 2006 393 2008
rect 359 1974 393 2006
rect 359 1904 393 1926
rect 359 1892 393 1904
rect 359 1836 393 1844
rect 359 1810 393 1836
rect 359 1734 393 1762
rect 359 1728 393 1734
rect 359 1666 393 1680
rect 359 1646 393 1666
rect 359 1564 393 1598
rect 515 2074 549 2090
rect 515 2056 549 2074
rect 515 2006 549 2008
rect 515 1974 549 2006
rect 515 1904 549 1926
rect 515 1892 549 1904
rect 515 1836 549 1844
rect 515 1810 549 1836
rect 515 1734 549 1762
rect 515 1728 549 1734
rect 515 1666 549 1680
rect 515 1646 549 1666
rect 436 1559 470 1593
rect 515 1564 549 1598
rect 735 2076 769 2093
rect 735 2059 769 2076
rect 735 2008 769 2020
rect 735 1986 769 2008
rect 735 1940 769 1947
rect 735 1913 769 1940
rect 735 1872 769 1874
rect 735 1840 769 1872
rect 735 1770 769 1801
rect 735 1767 769 1770
rect 735 1702 769 1728
rect 735 1694 769 1702
rect 735 1634 769 1655
rect 735 1621 769 1634
rect 735 1566 769 1582
rect 735 1548 769 1566
rect 436 1504 470 1521
rect 228 1470 230 1504
rect 230 1470 262 1504
rect 300 1470 332 1504
rect 332 1470 334 1504
rect 436 1487 454 1504
rect 454 1487 470 1504
rect 735 1498 769 1509
rect 735 1475 769 1498
rect 891 2246 925 2257
rect 891 2223 925 2246
rect 891 2178 925 2182
rect 891 2148 925 2178
rect 891 2076 925 2107
rect 891 2073 925 2076
rect 891 2008 925 2032
rect 891 1998 925 2008
rect 891 1940 925 1957
rect 891 1923 925 1940
rect 891 1872 925 1882
rect 891 1848 925 1872
rect 891 1804 925 1807
rect 891 1773 925 1804
rect 891 1702 925 1732
rect 891 1698 925 1702
rect 891 1634 925 1657
rect 891 1623 925 1634
rect 891 1566 925 1582
rect 891 1548 925 1566
rect 891 1498 925 1506
rect 891 1472 925 1498
rect 891 1396 925 1430
rect 1001 2212 1035 2245
rect 1001 2211 1035 2212
rect 1001 2144 1035 2171
rect 1001 2137 1035 2144
rect 1001 2076 1035 2097
rect 1001 2063 1035 2076
rect 1001 2008 1035 2023
rect 1001 1989 1035 2008
rect 1001 1940 1035 1949
rect 1001 1915 1035 1940
rect 1001 1872 1035 1875
rect 1001 1841 1035 1872
rect 1001 1770 1035 1801
rect 1001 1767 1035 1770
rect 1001 1702 1035 1727
rect 1001 1693 1035 1702
rect 1001 1634 1035 1653
rect 1001 1619 1035 1634
rect 1001 1566 1035 1579
rect 1001 1545 1035 1566
rect 1001 1498 1035 1505
rect 1001 1471 1035 1498
rect 1001 1396 1035 1430
rect 1469 2350 1503 2384
rect 1157 2280 1191 2310
rect 1157 2276 1191 2280
rect 1157 2212 1191 2236
rect 1157 2202 1191 2212
rect 1157 2144 1191 2162
rect 1157 2128 1191 2144
rect 1157 2076 1191 2088
rect 1157 2054 1191 2076
rect 1157 2008 1191 2014
rect 1157 1980 1191 2008
rect 1157 1906 1191 1940
rect 1157 1838 1191 1866
rect 1157 1832 1191 1838
rect 1157 1770 1191 1792
rect 1157 1758 1191 1770
rect 1157 1702 1191 1718
rect 1157 1684 1191 1702
rect 1157 1634 1191 1644
rect 1157 1610 1191 1634
rect 1157 1566 1191 1570
rect 1157 1536 1191 1566
rect 1313 2212 1347 2245
rect 1313 2211 1347 2212
rect 1313 2144 1347 2171
rect 1313 2137 1347 2144
rect 1313 2076 1347 2097
rect 1313 2063 1347 2076
rect 1313 2008 1347 2023
rect 1313 1989 1347 2008
rect 1313 1940 1347 1949
rect 1313 1915 1347 1940
rect 1313 1872 1347 1875
rect 1313 1841 1347 1872
rect 1313 1770 1347 1801
rect 1313 1767 1347 1770
rect 1313 1702 1347 1727
rect 1313 1693 1347 1702
rect 1313 1634 1347 1653
rect 1313 1619 1347 1634
rect 1313 1566 1347 1579
rect 1313 1545 1347 1566
rect 1313 1498 1347 1505
rect 1313 1471 1347 1498
rect 1313 1396 1347 1430
rect 1781 2350 1815 2384
rect 1469 2280 1503 2310
rect 1469 2276 1503 2280
rect 1469 2212 1503 2236
rect 1469 2202 1503 2212
rect 1469 2144 1503 2162
rect 1469 2128 1503 2144
rect 1469 2076 1503 2088
rect 1469 2054 1503 2076
rect 1469 2008 1503 2014
rect 1469 1980 1503 2008
rect 1469 1906 1503 1940
rect 1469 1838 1503 1866
rect 1469 1832 1503 1838
rect 1469 1770 1503 1792
rect 1469 1758 1503 1770
rect 1469 1702 1503 1718
rect 1469 1684 1503 1702
rect 1469 1634 1503 1644
rect 1469 1610 1503 1634
rect 1469 1566 1503 1570
rect 1469 1536 1503 1566
rect 1625 2212 1659 2245
rect 1625 2211 1659 2212
rect 1625 2144 1659 2171
rect 1625 2137 1659 2144
rect 1625 2076 1659 2097
rect 1625 2063 1659 2076
rect 1625 2008 1659 2023
rect 1625 1989 1659 2008
rect 1625 1940 1659 1949
rect 1625 1915 1659 1940
rect 1625 1872 1659 1875
rect 1625 1841 1659 1872
rect 1625 1770 1659 1801
rect 1625 1767 1659 1770
rect 1625 1702 1659 1727
rect 1625 1693 1659 1702
rect 1625 1634 1659 1653
rect 1625 1619 1659 1634
rect 1625 1566 1659 1579
rect 1625 1545 1659 1566
rect 1625 1498 1659 1505
rect 1625 1471 1659 1498
rect 1625 1396 1659 1430
rect 1781 2280 1815 2310
rect 1781 2276 1815 2280
rect 1781 2212 1815 2236
rect 1781 2202 1815 2212
rect 1781 2144 1815 2162
rect 1781 2128 1815 2144
rect 1781 2076 1815 2088
rect 1781 2054 1815 2076
rect 1781 2008 1815 2014
rect 1781 1980 1815 2008
rect 1781 1906 1815 1940
rect 1781 1838 1815 1866
rect 1781 1832 1815 1838
rect 1781 1770 1815 1792
rect 1781 1758 1815 1770
rect 1781 1702 1815 1718
rect 1781 1684 1815 1702
rect 1781 1634 1815 1644
rect 1781 1610 1815 1634
rect 1781 1566 1815 1570
rect 1781 1536 1815 1566
rect 736 1302 762 1336
rect 762 1302 770 1336
rect 808 1302 830 1336
rect 830 1302 842 1336
rect 1058 1302 1062 1336
rect 1062 1302 1092 1336
rect 1134 1302 1136 1336
rect 1136 1302 1168 1336
rect 1210 1302 1243 1336
rect 1243 1302 1244 1336
rect 1286 1302 1316 1336
rect 1316 1302 1320 1336
rect 1362 1302 1389 1336
rect 1389 1302 1396 1336
rect 1438 1302 1462 1336
rect 1462 1302 1472 1336
rect 1514 1302 1535 1336
rect 1535 1302 1548 1336
rect 1590 1302 1608 1336
rect 1608 1302 1624 1336
rect 1665 1302 1681 1336
rect 1681 1302 1699 1336
rect 102 1194 106 1228
rect 106 1194 136 1228
rect 187 1194 210 1228
rect 210 1194 221 1228
rect 272 1194 279 1228
rect 279 1194 306 1228
rect 357 1194 383 1228
rect 383 1194 391 1228
rect 442 1194 452 1228
rect 452 1194 476 1228
rect 622 1194 644 1228
rect 644 1194 656 1228
rect 703 1194 713 1228
rect 713 1194 737 1228
rect 784 1194 816 1228
rect 816 1194 818 1228
rect 865 1194 885 1228
rect 885 1194 899 1228
rect 1095 1194 1118 1228
rect 1118 1194 1129 1228
rect 1167 1194 1186 1228
rect 1186 1194 1201 1228
rect 1414 1194 1418 1228
rect 1418 1194 1448 1228
rect 1508 1194 1522 1228
rect 1522 1194 1542 1228
rect 1601 1194 1626 1228
rect 1626 1194 1635 1228
rect 1694 1194 1695 1228
rect 1695 1194 1728 1228
rect 45 1100 79 1134
rect 357 1100 391 1134
rect 45 1042 79 1059
rect 45 1025 79 1042
rect 45 974 79 984
rect 45 950 79 974
rect 45 906 79 909
rect -235 878 -201 882
rect -235 848 -201 878
rect -235 776 -201 802
rect -235 768 -201 776
rect -235 708 -201 722
rect -235 688 -201 708
rect -235 640 -201 641
rect -235 607 -201 640
rect -235 538 -201 560
rect -235 526 -201 538
rect -235 470 -201 479
rect -235 445 -201 470
rect -235 368 -201 398
rect -235 364 -201 368
rect -79 878 -45 882
rect -79 848 -45 878
rect -79 776 -45 802
rect -79 768 -45 776
rect -79 708 -45 722
rect -79 688 -45 708
rect -79 640 -45 641
rect -79 607 -45 640
rect -79 538 -45 560
rect -79 526 -45 538
rect -79 470 -45 479
rect -79 445 -45 470
rect -79 368 -45 398
rect -79 364 -45 368
rect 45 875 79 906
rect 45 804 79 834
rect 45 800 79 804
rect 45 736 79 759
rect 45 725 79 736
rect 45 668 79 684
rect 45 650 79 668
rect 45 600 79 609
rect 45 575 79 600
rect 45 532 79 534
rect 45 500 79 532
rect 45 430 79 459
rect 45 425 79 430
rect 45 362 79 384
rect 45 350 79 362
rect 201 974 235 998
rect 201 964 235 974
rect 201 906 235 924
rect 201 890 235 906
rect 201 838 235 850
rect 201 816 235 838
rect 201 770 235 776
rect 201 742 235 770
rect 201 668 235 702
rect 201 600 235 628
rect 201 594 235 600
rect 201 532 235 554
rect 201 520 235 532
rect 201 464 235 480
rect 201 446 235 464
rect 201 396 235 405
rect 201 371 235 396
rect 201 328 235 330
rect 201 296 235 328
rect 201 226 235 255
rect 201 221 235 226
rect 201 158 235 180
rect 201 146 235 158
rect 669 1100 703 1134
rect 357 1042 391 1059
rect 357 1025 391 1042
rect 357 974 391 984
rect 357 950 391 974
rect 357 906 391 909
rect 357 875 391 906
rect 357 804 391 834
rect 357 800 391 804
rect 357 736 391 759
rect 357 725 391 736
rect 357 668 391 684
rect 357 650 391 668
rect 357 600 391 609
rect 357 575 391 600
rect 357 532 391 534
rect 357 500 391 532
rect 357 430 391 459
rect 357 425 391 430
rect 357 362 391 384
rect 357 350 391 362
rect 513 974 547 998
rect 513 964 547 974
rect 513 906 547 924
rect 513 890 547 906
rect 513 838 547 850
rect 513 816 547 838
rect 513 770 547 776
rect 513 742 547 770
rect 513 668 547 702
rect 513 600 547 628
rect 513 594 547 600
rect 513 532 547 554
rect 513 520 547 532
rect 513 464 547 480
rect 513 446 547 464
rect 513 396 547 405
rect 513 371 547 396
rect 513 328 547 330
rect 513 296 547 328
rect 513 226 547 255
rect 513 221 547 226
rect 513 158 547 180
rect 513 146 547 158
rect 981 1100 1015 1134
rect 669 1042 703 1059
rect 669 1025 703 1042
rect 669 974 703 984
rect 669 950 703 974
rect 669 906 703 909
rect 669 875 703 906
rect 669 804 703 834
rect 669 800 703 804
rect 669 736 703 759
rect 669 725 703 736
rect 669 668 703 684
rect 669 650 703 668
rect 669 600 703 609
rect 669 575 703 600
rect 669 532 703 534
rect 669 500 703 532
rect 669 430 703 459
rect 669 425 703 430
rect 669 362 703 384
rect 669 350 703 362
rect 825 974 859 998
rect 825 964 859 974
rect 825 906 859 924
rect 825 890 859 906
rect 825 838 859 850
rect 825 816 859 838
rect 825 770 859 776
rect 825 742 859 770
rect 825 668 859 702
rect 825 600 859 628
rect 825 594 859 600
rect 825 532 859 554
rect 825 520 859 532
rect 825 464 859 480
rect 825 446 859 464
rect 825 396 859 405
rect 825 371 859 396
rect 825 328 859 330
rect 825 296 859 328
rect 825 226 859 255
rect 825 221 859 226
rect 825 158 859 180
rect 825 146 859 158
rect 1247 1093 1281 1127
rect 981 1042 1015 1061
rect 981 1027 1015 1042
rect 981 974 1015 988
rect 981 954 1015 974
rect 981 906 1015 915
rect 981 881 1015 906
rect 981 838 1015 842
rect 981 808 1015 838
rect 981 736 1015 769
rect 981 735 1015 736
rect 981 668 1015 696
rect 981 662 1015 668
rect 981 600 1015 623
rect 981 589 1015 600
rect 981 532 1015 550
rect 1091 1068 1125 1073
rect 1091 1039 1125 1068
rect 1091 966 1125 993
rect 1091 959 1125 966
rect 1091 898 1125 913
rect 1091 879 1125 898
rect 1091 830 1125 833
rect 1091 799 1125 830
rect 1091 728 1125 753
rect 1091 719 1125 728
rect 1091 660 1125 673
rect 1091 639 1125 660
rect 1091 558 1125 592
rect 1247 1034 1281 1051
rect 1247 1017 1281 1034
rect 1247 966 1281 975
rect 1247 941 1281 966
rect 1247 898 1281 899
rect 1247 865 1281 898
rect 1247 796 1281 823
rect 1247 789 1281 796
rect 1247 728 1281 746
rect 1247 712 1281 728
rect 1247 660 1281 669
rect 1247 635 1281 660
rect 1247 558 1281 592
rect 1357 1100 1391 1134
rect 1669 1100 1703 1134
rect 1357 1042 1391 1059
rect 1357 1025 1391 1042
rect 1357 974 1391 984
rect 1357 950 1391 974
rect 1357 906 1391 909
rect 1357 875 1391 906
rect 1357 804 1391 834
rect 1357 800 1391 804
rect 1357 736 1391 759
rect 1357 725 1391 736
rect 1357 668 1391 684
rect 1357 650 1391 668
rect 1357 600 1391 609
rect 1357 575 1391 600
rect 981 516 1015 532
rect 981 464 1015 477
rect 981 443 1015 464
rect 981 396 1015 404
rect 981 370 1015 396
rect 981 328 1015 330
rect 981 296 1015 328
rect 1357 532 1391 534
rect 1357 500 1391 532
rect 1357 430 1391 459
rect 1357 425 1391 430
rect 1357 362 1391 384
rect 1357 350 1391 362
rect 1513 974 1547 980
rect 1513 946 1547 974
rect 1513 906 1547 908
rect 1513 874 1547 906
rect 1513 804 1547 836
rect 1513 802 1547 804
rect 1513 736 1547 764
rect 1513 730 1547 736
rect 1513 668 1547 691
rect 1513 657 1547 668
rect 1513 600 1547 618
rect 1513 584 1547 600
rect 1513 532 1547 545
rect 1513 511 1547 532
rect 1513 464 1547 472
rect 1513 438 1547 464
rect 1513 396 1547 399
rect 1513 365 1547 396
rect 1513 294 1547 326
rect 1513 292 1547 294
rect 1513 226 1547 253
rect 1513 219 1547 226
rect 1513 158 1547 180
rect 1513 146 1547 158
rect 1669 1042 1703 1059
rect 1669 1025 1703 1042
rect 1669 974 1703 984
rect 1669 950 1703 974
rect 1669 906 1703 909
rect 1669 875 1703 906
rect 1669 804 1703 834
rect 1669 800 1703 804
rect 1669 736 1703 759
rect 1669 725 1703 736
rect 1669 668 1703 684
rect 1669 650 1703 668
rect 1669 600 1703 609
rect 1669 575 1703 600
rect 1669 532 1703 534
rect 1669 500 1703 532
rect 1669 430 1703 459
rect 1669 425 1703 430
rect 1669 362 1703 384
rect 1669 350 1703 362
rect 1825 974 1859 998
rect 1825 964 1859 974
rect 1825 906 1859 924
rect 1825 890 1859 906
rect 1825 838 1859 850
rect 1825 816 1859 838
rect 1825 770 1859 776
rect 1825 742 1859 770
rect 1825 668 1859 702
rect 1825 600 1859 628
rect 1825 594 1859 600
rect 1825 532 1859 554
rect 1825 520 1859 532
rect 1825 464 1859 480
rect 1825 446 1859 464
rect 1825 396 1859 405
rect 1825 371 1859 396
rect 1825 328 1859 330
rect 1825 296 1859 328
rect 1825 226 1859 255
rect 1825 221 1859 226
rect 1825 158 1859 180
rect 1825 146 1859 158
rect 38 36 62 70
rect 62 36 72 70
rect 113 36 132 70
rect 132 36 147 70
rect 188 36 202 70
rect 202 36 222 70
rect 262 36 272 70
rect 272 36 296 70
rect 336 36 342 70
rect 342 36 370 70
rect 410 36 412 70
rect 412 36 444 70
rect 484 36 516 70
rect 516 36 518 70
rect 558 36 586 70
rect 586 36 592 70
rect 632 36 656 70
rect 656 36 666 70
rect 706 36 726 70
rect 726 36 740 70
rect 780 36 796 70
rect 796 36 814 70
rect 854 36 866 70
rect 866 36 888 70
rect 928 36 936 70
rect 936 36 962 70
rect 1002 36 1006 70
rect 1006 36 1036 70
rect 1076 36 1110 70
rect 1150 36 1182 70
rect 1182 36 1184 70
rect 1224 36 1252 70
rect 1252 36 1258 70
rect 1298 36 1321 70
rect 1321 36 1332 70
rect 1372 36 1390 70
rect 1390 36 1406 70
rect 1446 36 1459 70
rect 1459 36 1480 70
rect 1520 36 1528 70
rect 1528 36 1554 70
rect 1594 36 1597 70
rect 1597 36 1628 70
rect 1668 36 1700 70
rect 1700 36 1702 70
rect 1742 36 1769 70
rect 1769 36 1776 70
rect 1816 36 1838 70
rect 1838 36 1850 70
<< metal1 >>
rect 55 2492 1833 2498
rect 55 2458 67 2492
rect 101 2458 142 2492
rect 176 2458 217 2492
rect 251 2458 292 2492
rect 326 2458 367 2492
rect 401 2458 442 2492
rect 476 2458 517 2492
rect 551 2458 592 2492
rect 626 2458 667 2492
rect 701 2458 742 2492
rect 776 2458 817 2492
rect 851 2458 892 2492
rect 926 2458 967 2492
rect 1001 2458 1042 2492
rect 1076 2458 1117 2492
rect 1151 2458 1192 2492
rect 1226 2458 1267 2492
rect 1301 2458 1342 2492
rect 1376 2458 1417 2492
rect 1451 2458 1491 2492
rect 1525 2458 1565 2492
rect 1599 2458 1639 2492
rect 1673 2458 1713 2492
rect 1747 2458 1787 2492
rect 1821 2458 1833 2492
rect 55 2384 1833 2458
rect 55 2350 735 2384
rect 769 2350 1157 2384
rect 1191 2350 1469 2384
rect 1503 2350 1781 2384
rect 1815 2350 1833 2384
rect 55 2312 1833 2350
rect 55 2298 735 2312
tri 319 2278 339 2298 ne
rect 339 2278 413 2298
tri 413 2278 433 2298 nw
tri 695 2278 715 2298 ne
rect 715 2278 735 2298
rect 769 2310 1833 2312
rect 769 2298 1157 2310
rect 769 2278 787 2298
tri 339 2276 341 2278 ne
rect 341 2276 411 2278
tri 411 2276 413 2278 nw
tri 715 2276 717 2278 ne
rect 717 2276 787 2278
tri 787 2276 809 2298 nw
tri 1117 2276 1139 2298 ne
rect 1139 2276 1157 2298
rect 1191 2298 1469 2310
rect 1191 2276 1209 2298
tri 1209 2276 1231 2298 nw
tri 1429 2276 1451 2298 ne
rect 1451 2276 1469 2298
rect 1503 2298 1781 2310
rect 1503 2276 1521 2298
tri 1521 2276 1543 2298 nw
tri 1741 2276 1763 2298 ne
rect 1763 2276 1781 2298
rect 1815 2298 1833 2310
rect 1815 2276 1821 2298
tri 1821 2286 1833 2298 nw
tri 341 2264 353 2276 ne
rect 194 2090 246 2102
rect 194 2056 203 2090
rect 237 2056 246 2090
rect 194 2008 246 2056
rect 194 1974 203 2008
rect 237 1974 246 2008
rect 194 1926 246 1974
rect 194 1892 203 1926
rect 237 1892 246 1926
rect 194 1844 246 1892
rect 194 1810 203 1844
rect 237 1810 246 1844
rect 194 1762 246 1810
rect 194 1728 203 1762
rect 237 1728 246 1762
rect 194 1689 246 1728
rect 194 1618 246 1637
rect 194 1564 203 1566
rect 237 1564 246 1566
rect 194 1552 246 1564
rect 353 2090 399 2276
tri 399 2264 411 2276 nw
tri 717 2264 729 2276 ne
rect 729 2269 780 2276
tri 780 2269 787 2276 nw
tri 1139 2269 1146 2276 ne
rect 1146 2269 1197 2276
rect 729 2239 775 2269
tri 775 2264 780 2269 nw
rect 729 2205 735 2239
rect 769 2205 775 2239
rect 729 2166 775 2205
rect 729 2132 735 2166
rect 769 2132 775 2166
rect 353 2056 359 2090
rect 393 2056 399 2090
rect 353 2008 399 2056
rect 353 1974 359 2008
rect 393 1974 399 2008
rect 353 1926 399 1974
rect 353 1892 359 1926
rect 393 1892 399 1926
rect 353 1844 399 1892
rect 353 1810 359 1844
rect 393 1810 399 1844
rect 353 1762 399 1810
rect 353 1728 359 1762
rect 393 1728 399 1762
rect 353 1680 399 1728
rect 353 1646 359 1680
rect 393 1646 399 1680
rect 353 1598 399 1646
rect 507 2090 559 2102
rect 507 2056 515 2090
rect 549 2056 559 2090
rect 507 2008 559 2056
rect 507 1974 515 2008
rect 549 1974 559 2008
rect 507 1926 559 1974
rect 507 1892 515 1926
rect 549 1892 559 1926
rect 507 1844 559 1892
rect 507 1810 515 1844
rect 549 1810 559 1844
rect 507 1762 559 1810
rect 507 1728 515 1762
rect 549 1728 559 1762
rect 507 1680 559 1728
rect 507 1674 515 1680
rect 549 1674 559 1680
rect 507 1610 559 1622
rect 353 1564 359 1598
rect 393 1564 399 1598
rect 353 1552 399 1564
rect 427 1604 479 1610
rect 427 1533 479 1552
rect 216 1504 346 1510
rect 216 1470 228 1504
rect 262 1470 300 1504
rect 334 1470 346 1504
rect 427 1475 479 1481
rect 216 1430 346 1470
tri 346 1430 374 1458 sw
tri 479 1430 507 1458 se
rect 507 1430 559 1558
rect 729 2093 775 2132
rect 729 2059 735 2093
rect 769 2059 775 2093
rect 729 2020 775 2059
rect 729 1986 735 2020
rect 769 1986 775 2020
rect 729 1947 775 1986
rect 729 1913 735 1947
rect 769 1913 775 1947
rect 729 1874 775 1913
rect 729 1840 735 1874
rect 769 1840 775 1874
rect 729 1801 775 1840
rect 729 1767 735 1801
rect 769 1767 775 1801
rect 729 1728 775 1767
rect 729 1694 735 1728
rect 769 1694 775 1728
rect 729 1655 775 1694
rect 729 1621 735 1655
rect 769 1621 775 1655
rect 729 1582 775 1621
rect 729 1548 735 1582
rect 769 1548 775 1582
rect 729 1509 775 1548
rect 729 1475 735 1509
rect 769 1475 775 1509
rect 729 1463 775 1475
rect 885 2257 931 2269
tri 1146 2264 1151 2269 ne
rect 885 2223 891 2257
rect 925 2223 931 2257
rect 885 2182 931 2223
rect 885 2148 891 2182
rect 925 2148 931 2182
rect 885 2107 931 2148
rect 885 2073 891 2107
rect 925 2073 931 2107
rect 885 2032 931 2073
rect 885 1998 891 2032
rect 925 1998 931 2032
rect 885 1957 931 1998
rect 885 1923 891 1957
rect 925 1923 931 1957
rect 885 1882 931 1923
rect 885 1848 891 1882
rect 925 1848 931 1882
rect 885 1807 931 1848
rect 885 1773 891 1807
rect 925 1773 931 1807
rect 885 1732 931 1773
rect 885 1698 891 1732
rect 925 1698 931 1732
rect 885 1657 931 1698
rect 885 1623 891 1657
rect 925 1623 931 1657
rect 885 1582 931 1623
rect 885 1548 891 1582
rect 925 1548 931 1582
rect 885 1506 931 1548
rect 885 1472 891 1506
rect 925 1472 931 1506
tri 559 1430 587 1458 sw
rect 885 1430 931 1472
rect 216 1424 374 1430
tri 374 1424 380 1430 sw
tri 473 1424 479 1430 se
rect 479 1424 587 1430
tri 587 1424 593 1430 sw
rect 216 1416 626 1424
tri 626 1416 634 1424 sw
rect 216 1396 634 1416
tri 634 1396 654 1416 sw
rect 885 1396 891 1430
rect 925 1396 931 1430
rect 216 1372 654 1396
tri 604 1344 632 1372 ne
rect 632 1346 654 1372
tri 654 1346 704 1396 sw
rect 885 1362 931 1396
rect 995 2245 1041 2257
rect 995 2211 1001 2245
rect 1035 2211 1041 2245
rect 995 2171 1041 2211
rect 995 2137 1001 2171
rect 1035 2137 1041 2171
rect 995 2097 1041 2137
rect 995 2063 1001 2097
rect 1035 2063 1041 2097
rect 995 2023 1041 2063
rect 995 1989 1001 2023
rect 1035 1989 1041 2023
rect 995 1949 1041 1989
rect 995 1915 1001 1949
rect 1035 1915 1041 1949
rect 995 1875 1041 1915
rect 995 1841 1001 1875
rect 1035 1841 1041 1875
rect 995 1801 1041 1841
rect 995 1767 1001 1801
rect 1035 1767 1041 1801
rect 995 1727 1041 1767
rect 995 1693 1001 1727
rect 1035 1693 1041 1727
rect 995 1653 1041 1693
rect 995 1619 1001 1653
rect 1035 1619 1041 1653
rect 995 1579 1041 1619
rect 995 1545 1001 1579
rect 1035 1545 1041 1579
rect 995 1505 1041 1545
rect 1151 2236 1197 2269
tri 1197 2264 1209 2276 nw
tri 1451 2264 1463 2276 ne
rect 1151 2202 1157 2236
rect 1191 2202 1197 2236
rect 1151 2162 1197 2202
rect 1151 2128 1157 2162
rect 1191 2128 1197 2162
rect 1151 2088 1197 2128
rect 1151 2054 1157 2088
rect 1191 2054 1197 2088
rect 1151 2014 1197 2054
rect 1151 1980 1157 2014
rect 1191 1980 1197 2014
rect 1151 1940 1197 1980
rect 1151 1906 1157 1940
rect 1191 1906 1197 1940
rect 1151 1866 1197 1906
rect 1151 1832 1157 1866
rect 1191 1832 1197 1866
rect 1151 1792 1197 1832
rect 1151 1758 1157 1792
rect 1191 1758 1197 1792
rect 1151 1718 1197 1758
rect 1151 1684 1157 1718
rect 1191 1684 1197 1718
rect 1151 1644 1197 1684
rect 1151 1610 1157 1644
rect 1191 1610 1197 1644
rect 1151 1570 1197 1610
rect 1151 1536 1157 1570
rect 1191 1536 1197 1570
rect 1151 1524 1197 1536
rect 1307 2245 1353 2257
rect 1307 2211 1313 2245
rect 1347 2211 1353 2245
rect 1307 2171 1353 2211
rect 1307 2137 1313 2171
rect 1347 2137 1353 2171
rect 1307 2097 1353 2137
rect 1307 2063 1313 2097
rect 1347 2063 1353 2097
rect 1307 2023 1353 2063
rect 1307 1989 1313 2023
rect 1347 1989 1353 2023
rect 1307 1949 1353 1989
rect 1307 1915 1313 1949
rect 1347 1915 1353 1949
rect 1307 1875 1353 1915
rect 1307 1841 1313 1875
rect 1347 1841 1353 1875
rect 1307 1801 1353 1841
rect 1307 1767 1313 1801
rect 1347 1767 1353 1801
rect 1307 1727 1353 1767
rect 1307 1693 1313 1727
rect 1347 1693 1353 1727
rect 1307 1653 1353 1693
rect 1307 1619 1313 1653
rect 1347 1619 1353 1653
rect 1307 1579 1353 1619
rect 1307 1545 1313 1579
rect 1347 1545 1353 1579
tri 1041 1505 1054 1518 sw
tri 1294 1505 1307 1518 se
rect 1307 1505 1353 1545
rect 1463 2236 1509 2276
tri 1509 2264 1521 2276 nw
tri 1763 2264 1775 2276 ne
rect 1463 2202 1469 2236
rect 1503 2202 1509 2236
rect 1463 2162 1509 2202
rect 1463 2128 1469 2162
rect 1503 2128 1509 2162
rect 1463 2088 1509 2128
rect 1463 2054 1469 2088
rect 1503 2054 1509 2088
rect 1463 2014 1509 2054
rect 1463 1980 1469 2014
rect 1503 1980 1509 2014
rect 1463 1940 1509 1980
rect 1463 1906 1469 1940
rect 1503 1906 1509 1940
rect 1463 1866 1509 1906
rect 1463 1832 1469 1866
rect 1503 1832 1509 1866
rect 1463 1792 1509 1832
rect 1463 1758 1469 1792
rect 1503 1758 1509 1792
rect 1463 1718 1509 1758
rect 1463 1684 1469 1718
rect 1503 1684 1509 1718
rect 1463 1644 1509 1684
rect 1463 1610 1469 1644
rect 1503 1610 1509 1644
rect 1463 1570 1509 1610
rect 1463 1536 1469 1570
rect 1503 1536 1509 1570
rect 1463 1524 1509 1536
rect 1619 2245 1665 2257
rect 1619 2211 1625 2245
rect 1659 2211 1665 2245
rect 1619 2171 1665 2211
rect 1619 2137 1625 2171
rect 1659 2137 1665 2171
rect 1619 2097 1665 2137
rect 1619 2063 1625 2097
rect 1659 2063 1665 2097
rect 1619 2023 1665 2063
rect 1619 1989 1625 2023
rect 1659 1989 1665 2023
rect 1619 1949 1665 1989
rect 1619 1915 1625 1949
rect 1659 1915 1665 1949
rect 1619 1875 1665 1915
rect 1619 1841 1625 1875
rect 1659 1841 1665 1875
rect 1619 1801 1665 1841
rect 1619 1767 1625 1801
rect 1659 1767 1665 1801
rect 1619 1727 1665 1767
rect 1619 1693 1625 1727
rect 1659 1693 1665 1727
rect 1619 1653 1665 1693
rect 1619 1619 1625 1653
rect 1659 1619 1665 1653
rect 1619 1579 1665 1619
rect 1619 1545 1625 1579
rect 1659 1545 1665 1579
tri 1353 1505 1366 1518 sw
tri 1606 1505 1619 1518 se
rect 1619 1505 1665 1545
rect 1775 2236 1821 2276
rect 1775 2202 1781 2236
rect 1815 2202 1821 2236
rect 1775 2162 1821 2202
rect 1775 2128 1781 2162
rect 1815 2128 1821 2162
rect 1775 2088 1821 2128
rect 1775 2054 1781 2088
rect 1815 2054 1821 2088
rect 1775 2014 1821 2054
rect 1775 1980 1781 2014
rect 1815 1980 1821 2014
rect 1775 1940 1821 1980
rect 1775 1906 1781 1940
rect 1815 1906 1821 1940
rect 1775 1866 1821 1906
rect 1775 1832 1781 1866
rect 1815 1832 1821 1866
rect 1775 1792 1821 1832
rect 1775 1758 1781 1792
rect 1815 1758 1821 1792
rect 1775 1718 1821 1758
rect 1775 1684 1781 1718
rect 1815 1684 1821 1718
rect 1775 1644 1821 1684
rect 1775 1610 1781 1644
rect 1815 1610 1821 1644
rect 1775 1570 1821 1610
rect 1775 1536 1781 1570
rect 1815 1536 1821 1570
rect 1775 1524 1821 1536
rect 995 1471 1001 1505
rect 1035 1484 1054 1505
tri 1054 1484 1075 1505 sw
tri 1273 1484 1294 1505 se
rect 1294 1484 1313 1505
rect 1035 1471 1313 1484
rect 1347 1484 1366 1505
tri 1366 1484 1387 1505 sw
tri 1585 1484 1606 1505 se
rect 1606 1484 1625 1505
rect 1347 1471 1625 1484
rect 1659 1484 1665 1505
tri 1665 1484 1699 1518 sw
rect 1659 1471 1903 1484
rect 995 1430 1903 1471
rect 995 1396 1001 1430
rect 1035 1396 1313 1430
rect 1347 1396 1625 1430
rect 1659 1396 1903 1430
tri 885 1346 901 1362 ne
rect 901 1346 931 1362
tri 931 1346 971 1386 sw
rect 995 1384 1903 1396
tri 1761 1350 1795 1384 ne
rect 632 1344 704 1346
tri 704 1344 706 1346 sw
tri 901 1344 903 1346 ne
rect 903 1344 1740 1346
rect 0 1336 523 1344
tri 523 1336 531 1344 sw
tri 632 1342 634 1344 ne
rect 634 1342 706 1344
tri 706 1342 708 1344 sw
tri 903 1342 905 1344 ne
rect 905 1342 1740 1344
tri 634 1336 640 1342 ne
rect 640 1336 854 1342
tri 905 1336 911 1342 ne
rect 911 1336 1740 1342
rect 0 1316 531 1336
tri 531 1316 551 1336 sw
tri 640 1316 660 1336 ne
rect 660 1316 736 1336
rect 0 1311 551 1316
tri 551 1311 556 1316 sw
tri 660 1311 665 1316 ne
rect 665 1311 736 1316
rect 0 1302 556 1311
tri 556 1302 565 1311 sw
tri 665 1302 674 1311 ne
rect 674 1302 736 1311
rect 770 1302 808 1336
rect 842 1302 854 1336
tri 911 1316 931 1336 ne
rect 931 1316 1058 1336
tri 931 1302 945 1316 ne
rect 945 1302 1058 1316
rect 1092 1302 1134 1336
rect 1168 1302 1210 1336
rect 1244 1302 1286 1336
rect 1320 1302 1362 1336
rect 1396 1302 1438 1336
rect 1472 1302 1514 1336
rect 1548 1302 1590 1336
rect 1624 1302 1665 1336
rect 1699 1302 1740 1336
rect 0 1296 565 1302
tri 565 1296 571 1302 sw
tri 674 1296 680 1302 ne
rect 680 1296 854 1302
tri 945 1296 951 1302 ne
rect 951 1296 1740 1302
rect 0 1292 571 1296
tri 501 1240 553 1292 ne
rect 553 1240 571 1292
rect 0 1228 488 1240
tri 553 1237 556 1240 ne
rect 556 1237 571 1240
tri 571 1237 630 1296 sw
tri 680 1290 686 1296 ne
rect 686 1290 854 1296
tri 1207 1290 1213 1296 ne
rect 1213 1290 1740 1296
tri 1213 1262 1241 1290 ne
tri 556 1234 559 1237 ne
rect 559 1234 911 1237
tri 559 1228 565 1234 ne
rect 565 1228 911 1234
rect 0 1194 102 1228
rect 136 1194 187 1228
rect 221 1194 272 1228
rect 306 1194 357 1228
rect 391 1194 442 1228
rect 476 1194 488 1228
tri 565 1194 599 1228 ne
rect 599 1194 622 1228
rect 656 1194 703 1228
rect 737 1194 784 1228
rect 818 1194 865 1228
rect 899 1194 911 1228
rect 0 1188 488 1194
tri 599 1188 605 1194 ne
rect 605 1188 911 1194
tri 605 1185 608 1188 ne
rect 608 1185 911 1188
rect 977 1228 1213 1234
rect 977 1194 1095 1228
rect 1129 1194 1167 1228
rect 1201 1194 1213 1228
rect 977 1188 1213 1194
rect 1241 1228 1740 1290
rect 1241 1194 1414 1228
rect 1448 1194 1508 1228
rect 1542 1194 1601 1228
rect 1635 1194 1694 1228
rect 1728 1194 1740 1228
rect 1241 1188 1740 1194
rect 977 1185 1052 1188
tri 1052 1185 1055 1188 nw
tri 943 1146 977 1180 se
rect 977 1146 1021 1185
tri 1021 1154 1052 1185 nw
rect 39 1134 117 1146
rect 39 1100 45 1134
rect 79 1100 117 1134
rect 39 1094 117 1100
rect 169 1094 188 1146
rect 240 1094 350 1146
rect 402 1094 421 1146
rect 473 1094 479 1146
rect 39 1086 479 1094
rect 507 1094 513 1146
rect 565 1094 583 1146
rect 635 1134 1021 1146
rect 635 1100 669 1134
rect 703 1100 981 1134
rect 1015 1100 1021 1134
rect 635 1094 1021 1100
rect 507 1086 1021 1094
rect 39 1073 106 1086
tri 106 1073 119 1086 nw
tri 317 1073 330 1086 ne
rect 330 1073 418 1086
tri 418 1073 431 1086 nw
tri 629 1073 642 1086 ne
rect 642 1073 730 1086
tri 730 1073 743 1086 nw
tri 941 1073 954 1086 ne
rect 954 1073 1021 1086
rect 1241 1127 1287 1188
tri 1287 1154 1321 1188 nw
tri 1769 1154 1795 1180 se
rect 1795 1154 1903 1384
tri 1761 1146 1769 1154 se
rect 1769 1146 1903 1154
rect 1241 1093 1247 1127
rect 1281 1093 1287 1127
rect 39 1061 94 1073
tri 94 1061 106 1073 nw
tri 330 1061 342 1073 ne
rect 342 1061 406 1073
tri 406 1061 418 1073 nw
tri 642 1061 654 1073 ne
rect 654 1061 718 1073
tri 718 1061 730 1073 nw
tri 954 1061 966 1073 ne
rect 966 1061 1021 1073
rect 39 1059 92 1061
tri 92 1059 94 1061 nw
tri 342 1059 344 1061 ne
rect 344 1059 404 1061
tri 404 1059 406 1061 nw
tri 654 1059 656 1061 ne
rect 656 1059 712 1061
rect -169 995 -94 1047
rect 39 1025 45 1059
rect 79 1025 85 1059
tri 85 1052 92 1059 nw
tri 344 1052 351 1059 ne
rect 39 984 85 1025
rect 351 1025 357 1059
rect 391 1055 400 1059
tri 400 1055 404 1059 nw
tri 656 1055 660 1059 ne
rect 391 1025 397 1055
tri 397 1052 400 1055 nw
rect 39 950 45 984
rect 79 950 85 984
rect -457 924 -298 933
tri -298 924 -289 933 sw
rect -457 909 -289 924
tri -289 909 -274 924 sw
rect 39 909 85 950
rect -457 894 -274 909
tri -274 894 -259 909 sw
rect -457 882 -195 894
rect -457 848 -235 882
rect -201 848 -195 882
rect -457 802 -195 848
rect -457 768 -235 802
rect -201 768 -195 802
rect -457 722 -195 768
rect -457 688 -235 722
rect -201 688 -195 722
rect -457 641 -195 688
rect -457 607 -235 641
rect -201 607 -195 641
rect -457 560 -195 607
rect -457 526 -235 560
rect -201 526 -195 560
rect -457 479 -195 526
rect -457 445 -235 479
rect -201 445 -195 479
rect -457 398 -195 445
rect -457 364 -235 398
rect -201 364 -195 398
rect -457 230 -195 364
rect -88 882 -36 894
rect -88 848 -79 882
rect -45 848 -36 882
rect -88 802 -36 848
rect -88 768 -79 802
rect -45 768 -36 802
rect -88 740 -36 768
rect -88 676 -36 688
rect -88 607 -79 624
rect -45 607 -36 624
rect -88 560 -36 607
rect -88 526 -79 560
rect -45 526 -36 560
rect -88 479 -36 526
rect -88 445 -79 479
rect -45 445 -36 479
rect -88 398 -36 445
rect -88 364 -79 398
rect -45 364 -36 398
rect -88 352 -36 364
rect 39 875 45 909
rect 79 875 85 909
rect 39 834 85 875
rect 39 800 45 834
rect 79 800 85 834
rect 39 759 85 800
rect 39 725 45 759
rect 79 725 85 759
rect 39 684 85 725
rect 39 650 45 684
rect 79 650 85 684
rect 39 609 85 650
rect 39 575 45 609
rect 79 575 85 609
rect 39 534 85 575
rect 39 500 45 534
rect 79 500 85 534
rect 39 459 85 500
rect 39 425 45 459
rect 79 425 85 459
rect 39 384 85 425
rect 39 350 45 384
rect 79 350 85 384
rect 39 338 85 350
rect 195 998 241 1010
rect 195 964 201 998
rect 235 964 241 998
rect 195 924 241 964
rect 195 890 201 924
rect 235 890 241 924
rect 195 850 241 890
rect 195 816 201 850
rect 235 816 241 850
rect 195 776 241 816
rect 195 742 201 776
rect 235 742 241 776
rect 195 702 241 742
rect 195 668 201 702
rect 235 668 241 702
rect 195 628 241 668
rect 195 594 201 628
rect 235 594 241 628
rect 195 554 241 594
rect 195 520 201 554
rect 235 520 241 554
rect 195 480 241 520
rect 195 446 201 480
rect 235 446 241 480
rect 195 405 241 446
rect 195 371 201 405
rect 235 371 241 405
rect 195 330 241 371
rect 351 984 397 1025
rect 660 1025 669 1059
rect 703 1025 712 1059
tri 712 1055 718 1061 nw
tri 966 1055 972 1061 ne
rect 972 1055 981 1061
tri 972 1052 975 1055 ne
rect 351 950 357 984
rect 391 950 397 984
rect 351 909 397 950
rect 351 875 357 909
rect 391 875 397 909
rect 351 834 397 875
rect 351 800 357 834
rect 391 800 397 834
rect 351 759 397 800
rect 351 725 357 759
rect 391 725 397 759
rect 351 684 397 725
rect 351 650 357 684
rect 391 650 397 684
rect 351 609 397 650
rect 351 575 357 609
rect 391 575 397 609
rect 351 534 397 575
rect 351 500 357 534
rect 391 500 397 534
rect 351 459 397 500
rect 351 425 357 459
rect 391 425 397 459
rect 351 384 397 425
rect 351 350 357 384
rect 391 350 397 384
rect 351 338 397 350
rect 507 998 553 1010
rect 507 964 513 998
rect 547 964 553 998
rect 507 924 553 964
rect 507 890 513 924
rect 547 890 553 924
rect 507 850 553 890
rect 507 816 513 850
rect 547 816 553 850
rect 507 776 553 816
rect 507 742 513 776
rect 547 742 553 776
rect 507 702 553 742
rect 507 668 513 702
rect 547 668 553 702
rect 507 628 553 668
rect 507 594 513 628
rect 547 594 553 628
rect 507 554 553 594
rect 507 520 513 554
rect 547 520 553 554
rect 507 480 553 520
rect 507 446 513 480
rect 547 446 553 480
rect 507 405 553 446
rect 507 371 513 405
rect 547 371 553 405
rect 195 296 201 330
rect 235 296 241 330
tri 186 255 195 264 se
rect 195 255 241 296
rect 507 330 553 371
rect 660 984 712 1025
rect 975 1027 981 1055
rect 1015 1027 1021 1061
rect 660 950 669 984
rect 703 950 712 984
rect 660 909 712 950
rect 660 875 669 909
rect 703 875 712 909
rect 660 834 712 875
rect 660 800 669 834
rect 703 800 712 834
rect 660 759 712 800
rect 660 740 669 759
rect 703 740 712 759
rect 660 684 712 688
rect 660 676 669 684
rect 703 676 712 684
rect 660 609 712 624
rect 660 575 669 609
rect 703 575 712 609
rect 660 534 712 575
rect 660 500 669 534
rect 703 500 712 534
rect 660 459 712 500
rect 660 425 669 459
rect 703 425 712 459
rect 660 384 712 425
rect 660 350 669 384
rect 703 350 712 384
rect 660 338 712 350
rect 819 998 865 1010
rect 819 964 825 998
rect 859 964 865 998
rect 819 924 865 964
rect 819 890 825 924
rect 859 890 865 924
rect 819 850 865 890
rect 819 816 825 850
rect 859 816 865 850
rect 819 776 865 816
rect 819 742 825 776
rect 859 742 865 776
rect 819 702 865 742
rect 819 668 825 702
rect 859 668 865 702
rect 819 628 865 668
rect 819 594 825 628
rect 859 594 865 628
rect 819 554 865 594
rect 819 520 825 554
rect 859 520 865 554
rect 819 480 865 520
rect 819 446 825 480
rect 859 446 865 480
rect 819 405 865 446
rect 819 371 825 405
rect 859 371 865 405
rect 507 296 513 330
rect 547 296 553 330
tri 241 255 250 264 sw
tri 498 255 507 264 se
rect 507 255 553 296
rect 819 330 865 371
rect 819 296 825 330
rect 859 296 865 330
tri 553 255 562 264 sw
tri 810 255 819 264 se
rect 819 255 865 296
rect 975 988 1021 1027
rect 975 954 981 988
rect 1015 954 1021 988
rect 975 915 1021 954
rect 975 881 981 915
rect 1015 881 1021 915
rect 975 842 1021 881
rect 975 808 981 842
rect 1015 808 1021 842
rect 975 769 1021 808
rect 975 735 981 769
rect 1015 735 1021 769
rect 975 696 1021 735
rect 975 662 981 696
rect 1015 662 1021 696
rect 975 623 1021 662
rect 975 589 981 623
rect 1015 589 1021 623
rect 975 550 1021 589
rect 975 516 981 550
rect 1015 516 1021 550
rect 975 477 1021 516
rect 975 443 981 477
rect 1015 443 1021 477
rect 975 404 1021 443
rect 975 370 981 404
rect 1015 370 1021 404
rect 975 330 1021 370
rect 975 296 981 330
rect 1015 296 1021 330
rect 975 284 1021 296
rect 1085 1073 1131 1085
rect 1085 1039 1091 1073
rect 1125 1039 1131 1073
rect 1085 993 1131 1039
rect 1085 959 1091 993
rect 1125 959 1131 993
rect 1085 913 1131 959
rect 1085 879 1091 913
rect 1125 879 1131 913
rect 1085 833 1131 879
rect 1085 799 1091 833
rect 1125 799 1131 833
rect 1085 753 1131 799
rect 1085 719 1091 753
rect 1125 719 1131 753
rect 1085 673 1131 719
rect 1085 639 1091 673
rect 1125 639 1131 673
rect 1085 592 1131 639
rect 1085 558 1091 592
rect 1125 558 1131 592
tri 865 255 874 264 sw
tri 1076 255 1085 264 se
rect 1085 255 1131 558
rect 1241 1051 1287 1093
rect 1241 1017 1247 1051
rect 1281 1017 1287 1051
rect 1241 975 1287 1017
rect 1241 941 1247 975
rect 1281 941 1287 975
rect 1241 899 1287 941
rect 1241 865 1247 899
rect 1281 865 1287 899
rect 1241 823 1287 865
rect 1241 789 1247 823
rect 1281 789 1287 823
rect 1241 746 1287 789
rect 1241 712 1247 746
rect 1281 712 1287 746
rect 1241 669 1287 712
rect 1241 635 1247 669
rect 1281 635 1287 669
rect 1241 592 1287 635
rect 1241 558 1247 592
rect 1281 558 1287 592
rect 1241 546 1287 558
rect 1351 1134 1903 1146
rect 1351 1100 1357 1134
rect 1391 1100 1669 1134
rect 1703 1100 1903 1134
rect 1351 1059 1903 1100
rect 1351 1025 1357 1059
rect 1391 1038 1669 1059
rect 1391 1025 1418 1038
tri 1418 1025 1431 1038 nw
tri 1629 1025 1642 1038 ne
rect 1642 1025 1669 1038
rect 1703 1038 1903 1059
rect 1703 1025 1715 1038
rect 1351 984 1397 1025
tri 1397 1004 1418 1025 nw
tri 1642 1004 1663 1025 ne
rect 1663 1010 1715 1025
tri 1715 1010 1743 1038 nw
rect 1351 950 1357 984
rect 1391 950 1397 984
rect 1351 909 1397 950
rect 1351 875 1357 909
rect 1391 875 1397 909
rect 1351 834 1397 875
rect 1351 800 1357 834
rect 1391 800 1397 834
rect 1351 759 1397 800
rect 1351 725 1357 759
rect 1391 725 1397 759
rect 1351 684 1397 725
rect 1351 650 1357 684
rect 1391 650 1397 684
rect 1351 609 1397 650
rect 1351 575 1357 609
rect 1391 575 1397 609
rect 1351 534 1397 575
rect 1351 500 1357 534
rect 1391 500 1397 534
rect 1351 459 1397 500
rect 1351 425 1357 459
rect 1391 425 1397 459
rect 1351 384 1397 425
rect 1351 350 1357 384
rect 1391 350 1397 384
rect 1351 338 1397 350
rect 1507 980 1553 992
rect 1507 946 1513 980
rect 1547 946 1553 980
rect 1507 908 1553 946
rect 1507 874 1513 908
rect 1547 874 1553 908
rect 1507 836 1553 874
rect 1507 802 1513 836
rect 1547 802 1553 836
rect 1507 764 1553 802
rect 1507 730 1513 764
rect 1547 730 1553 764
rect 1507 691 1553 730
rect 1507 657 1513 691
rect 1547 657 1553 691
rect 1507 618 1553 657
rect 1507 584 1513 618
rect 1547 584 1553 618
rect 1507 545 1553 584
rect 1507 511 1513 545
rect 1547 511 1553 545
rect 1507 472 1553 511
rect 1507 438 1513 472
rect 1547 438 1553 472
rect 1507 399 1553 438
rect 1507 365 1513 399
rect 1547 365 1553 399
rect 1507 326 1553 365
rect 1663 984 1709 1010
tri 1709 1004 1715 1010 nw
rect 1663 950 1669 984
rect 1703 950 1709 984
rect 1663 909 1709 950
rect 1663 875 1669 909
rect 1703 875 1709 909
rect 1663 834 1709 875
rect 1663 800 1669 834
rect 1703 800 1709 834
rect 1663 759 1709 800
rect 1663 725 1669 759
rect 1703 725 1709 759
rect 1663 684 1709 725
rect 1663 650 1669 684
rect 1703 650 1709 684
rect 1663 609 1709 650
rect 1663 575 1669 609
rect 1703 575 1709 609
rect 1663 534 1709 575
rect 1663 500 1669 534
rect 1703 500 1709 534
rect 1663 459 1709 500
rect 1663 425 1669 459
rect 1703 425 1709 459
rect 1663 384 1709 425
rect 1663 350 1669 384
rect 1703 350 1709 384
rect 1663 338 1709 350
rect 1819 998 1865 1010
rect 1819 964 1825 998
rect 1859 964 1865 998
rect 1819 924 1865 964
rect 1819 890 1825 924
rect 1859 890 1865 924
rect 1819 850 1865 890
rect 1819 816 1825 850
rect 1859 816 1865 850
rect 1819 776 1865 816
rect 1819 742 1825 776
rect 1859 742 1865 776
rect 1819 702 1865 742
rect 1819 668 1825 702
rect 1859 668 1865 702
rect 1819 628 1865 668
rect 1819 594 1825 628
rect 1859 594 1865 628
rect 1819 554 1865 594
rect 1819 520 1825 554
rect 1859 520 1865 554
rect 1819 480 1865 520
rect 1819 446 1825 480
rect 1859 446 1865 480
rect 1819 405 1865 446
rect 1819 371 1825 405
rect 1859 371 1865 405
rect 1507 292 1513 326
rect 1547 292 1553 326
tri 1131 255 1140 264 sw
tri 1498 255 1507 264 se
rect 1507 255 1553 292
rect 1819 330 1865 371
rect 1819 296 1825 330
rect 1859 296 1865 330
tri 1553 255 1562 264 sw
tri 1810 255 1819 264 se
rect 1819 255 1865 296
tri 181 250 186 255 se
rect 186 250 201 255
tri -195 230 -175 250 sw
tri 161 230 181 250 se
rect 181 230 201 250
rect -457 221 201 230
rect 235 230 250 255
tri 250 230 275 255 sw
tri 473 230 498 255 se
rect 498 230 513 255
rect 235 221 513 230
rect 547 230 562 255
tri 562 230 587 255 sw
tri 785 230 810 255 se
rect 810 230 825 255
rect 547 221 825 230
rect 859 253 874 255
tri 874 253 876 255 sw
tri 1074 253 1076 255 se
rect 1076 253 1140 255
tri 1140 253 1142 255 sw
tri 1496 253 1498 255 se
rect 1498 253 1562 255
rect 859 230 876 253
tri 876 230 899 253 sw
tri 1051 230 1074 253 se
rect 1074 230 1142 253
tri 1142 230 1165 253 sw
tri 1473 230 1496 253 se
rect 1496 230 1513 253
rect 859 221 1513 230
rect -457 219 1513 221
rect 1547 230 1562 253
tri 1562 230 1587 255 sw
tri 1785 230 1810 255 se
rect 1810 230 1825 255
rect 1547 221 1825 230
rect 1859 230 1865 255
tri 1865 230 1899 264 sw
rect 1859 221 1903 230
rect 1547 219 1903 221
rect -457 180 1903 219
rect -457 146 201 180
rect 235 146 513 180
rect 547 146 825 180
rect 859 146 1513 180
rect 1547 146 1825 180
rect 1859 146 1903 180
rect -457 70 1903 146
rect -457 36 38 70
rect 72 36 113 70
rect 147 36 188 70
rect 222 36 262 70
rect 296 36 336 70
rect 370 36 410 70
rect 444 36 484 70
rect 518 36 558 70
rect 592 36 632 70
rect 666 36 706 70
rect 740 36 780 70
rect 814 36 854 70
rect 888 36 928 70
rect 962 36 1002 70
rect 1036 36 1076 70
rect 1110 36 1150 70
rect 1184 36 1224 70
rect 1258 36 1298 70
rect 1332 36 1372 70
rect 1406 36 1446 70
rect 1480 36 1520 70
rect 1554 36 1594 70
rect 1628 36 1668 70
rect 1702 36 1742 70
rect 1776 36 1816 70
rect 1850 36 1903 70
rect -457 30 1903 36
<< via1 >>
rect 194 1680 246 1689
rect 194 1646 203 1680
rect 203 1646 237 1680
rect 237 1646 246 1680
rect 194 1637 246 1646
rect 194 1598 246 1618
rect 194 1566 203 1598
rect 203 1566 237 1598
rect 237 1566 246 1598
rect 507 1646 515 1674
rect 515 1646 549 1674
rect 549 1646 559 1674
rect 507 1622 559 1646
rect 427 1593 479 1604
rect 427 1559 436 1593
rect 436 1559 470 1593
rect 470 1559 479 1593
rect 427 1552 479 1559
rect 427 1521 479 1533
rect 427 1487 436 1521
rect 436 1487 470 1521
rect 470 1487 479 1521
rect 427 1481 479 1487
rect 507 1598 559 1610
rect 507 1564 515 1598
rect 515 1564 549 1598
rect 549 1564 559 1598
rect 507 1558 559 1564
rect 117 1094 169 1146
rect 188 1094 240 1146
rect 350 1134 402 1146
rect 350 1100 357 1134
rect 357 1100 391 1134
rect 391 1100 402 1134
rect 350 1094 402 1100
rect 421 1094 473 1146
rect 513 1094 565 1146
rect 583 1094 635 1146
rect -88 722 -36 740
rect -88 688 -79 722
rect -79 688 -45 722
rect -45 688 -36 722
rect -88 641 -36 676
rect -88 624 -79 641
rect -79 624 -45 641
rect -45 624 -36 641
rect 660 725 669 740
rect 669 725 703 740
rect 703 725 712 740
rect 660 688 712 725
rect 660 650 669 676
rect 669 650 703 676
rect 703 650 712 676
rect 660 624 712 650
<< metal2 >>
rect 194 1689 246 1695
rect 194 1618 246 1637
rect 507 1674 559 1680
rect 507 1610 559 1622
tri 160 1146 194 1180 se
rect 194 1146 246 1566
rect 427 1604 479 1610
rect 427 1533 479 1552
tri 393 1146 427 1180 se
rect 427 1146 479 1481
rect 111 1094 117 1146
rect 169 1094 188 1146
rect 240 1094 246 1146
rect 344 1094 350 1146
rect 402 1094 421 1146
rect 473 1094 479 1146
rect 507 1146 559 1558
tri 559 1146 593 1180 sw
rect 507 1094 513 1146
rect 565 1094 583 1146
rect 635 1094 641 1146
rect -88 740 712 746
rect -36 688 660 740
rect -88 676 712 688
rect -36 624 660 676
rect -88 618 712 624
use sky130_fd_pr__nfet_01v8__example_55959141808550  sky130_fd_pr__nfet_01v8__example_55959141808550_2
timestamp 1619862920
transform 1 0 1402 0 1 146
box -28 0 440 471
use sky130_fd_pr__nfet_01v8__example_55959141808550  sky130_fd_pr__nfet_01v8__example_55959141808550_1
timestamp 1619862920
transform 1 0 558 0 1 146
box -28 0 440 471
use sky130_fd_pr__nfet_01v8__example_55959141808550  sky130_fd_pr__nfet_01v8__example_55959141808550_0
timestamp 1619862920
transform 1 0 90 0 1 146
box -28 0 440 471
use sky130_fd_pr__nfet_01v8__example_55959141808528  sky130_fd_pr__nfet_01v8__example_55959141808528_1
timestamp 1619862920
transform 1 0 1136 0 1 546
box -28 0 128 267
use sky130_fd_pr__nfet_01v8__example_55959141808528  sky130_fd_pr__nfet_01v8__example_55959141808528_0
timestamp 1619862920
transform 1 0 -190 0 1 356
box -28 0 128 267
use sky130_fd_pr__pfet_01v8__example_55959141808537  sky130_fd_pr__pfet_01v8__example_55959141808537_0
timestamp 1619862920
transform 1 0 1046 0 1 1384
box -28 0 752 471
use sky130_fd_pr__pfet_01v8__example_55959141808548  sky130_fd_pr__pfet_01v8__example_55959141808548_0
timestamp 1619862920
transform 1 0 780 0 1 1384
box -28 0 128 471
use sky130_fd_pr__pfet_01v8__example_55959141808549  sky130_fd_pr__pfet_01v8__example_55959141808549_1
timestamp 1619862920
transform 1 0 404 0 1 1552
box -28 0 128 267
use sky130_fd_pr__pfet_01v8__example_55959141808549  sky130_fd_pr__pfet_01v8__example_55959141808549_0
timestamp 1619862920
transform 1 0 248 0 1 1552
box -28 0 128 267
<< labels >>
flabel metal1 s 0 1188 67 1240 3 FreeSans 520 0 0 0 IN
port 1 nsew
flabel metal1 s 0 1292 56 1344 3 FreeSans 520 0 0 0 INB
port 2 nsew
flabel metal1 s 64 2315 228 2452 3 FreeSans 520 0 0 0 VDDIO_Q
port 3 nsew
flabel metal1 s 12 47 95 123 3 FreeSans 520 0 0 0 VSSD
port 4 nsew
flabel metal1 s 1843 1228 1888 1353 3 FreeSans 520 0 0 0 OUT
port 5 nsew
flabel metal1 s 1421 1260 1570 1319 3 FreeSans 520 0 0 0 OUT_B
port 6 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 36244536
string GDS_START 36200720
<< end >>
