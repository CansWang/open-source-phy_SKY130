magic
tech sky130A
magscale 1 2
timestamp 1619862920
<< checkpaint >>
rect -1288 -1260 1388 1345
use sky130_fd_pr__hvdfm1sd__example_55959141808242  sky130_fd_pr__hvdfm1sd__example_55959141808242_0
timestamp 1619862920
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808242  sky130_fd_pr__hvdfm1sd__example_55959141808242_1
timestamp 1619862920
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 128 85 128 85 0 FreeSans 300 0 0 0 D
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 665896
string GDS_START 664970
<< end >>
