magic
tech sky130A
magscale 1 2
timestamp 1619240079
<< error_p >>
rect 254 37537 320 40000
rect 15000 37537 15066 40000
<< error_s >>
rect 254 35157 320 37537
rect 15000 35157 15066 37537
rect 2114 34342 2196 34375
rect 2054 34282 2213 34315
rect 1985 34250 1987 34274
rect 1925 34138 1938 34214
rect 1985 34153 1998 34250
rect 2198 34153 2213 34282
rect 1856 34084 1938 34138
rect 2258 34100 2273 34364
rect 12709 34100 12725 34364
rect 12786 34342 12868 34375
rect 12769 34282 12928 34315
rect 12769 34153 12785 34282
rect 12995 34250 12997 34274
rect 12984 34153 12997 34250
rect 2258 34082 2342 34100
rect 12640 34082 12725 34100
rect 13044 34138 13057 34214
rect 13044 34084 13126 34138
rect 2258 34079 2355 34082
rect 12627 34079 12725 34082
rect 1796 34024 1998 34078
rect 1670 33814 1692 33917
rect 1567 33787 1692 33814
rect 1730 33814 1752 33977
rect 2110 33850 2155 34078
rect 2170 34019 2295 34040
rect 12687 34019 12812 34040
rect 2170 33910 2215 34019
rect 12767 33910 12812 34019
rect 12827 33850 12872 34078
rect 12984 34024 13186 34078
rect 13230 33814 13252 33977
rect 1730 33812 1891 33814
rect 13091 33812 13252 33814
rect 1730 33778 2037 33812
rect 12945 33778 13252 33812
rect 13290 33814 13312 33917
rect 13290 33787 13415 33814
rect 1507 33727 1831 33754
rect 1670 33718 1831 33727
rect 1346 33494 1364 33589
rect 1239 33459 1364 33494
rect 1406 33494 1424 33636
rect 1792 33562 1831 33718
rect 1852 33718 1977 33752
rect 13005 33718 13130 33752
rect 1852 33622 1891 33718
rect 13091 33622 13130 33718
rect 13151 33727 13475 33754
rect 13151 33718 13312 33727
rect 13151 33562 13190 33718
rect 13558 33494 13576 33636
rect 1406 33487 1571 33494
rect 13411 33487 13576 33494
rect 1406 33454 1712 33487
rect 13270 33454 13576 33487
rect 13618 33494 13636 33589
rect 13618 33459 13743 33494
rect 1179 33399 1511 33434
rect 1346 33394 1511 33399
rect 1467 33237 1511 33394
rect 1527 33394 1652 33427
rect 13330 33394 13455 33427
rect 1527 33297 1571 33394
rect 13411 33297 13455 33394
rect 13471 33399 13803 33434
rect 13471 33394 13636 33399
rect 13471 33237 13515 33394
rect 1086 33134 1511 33168
rect 13471 33134 13896 33168
rect 1026 33107 1484 33108
rect 1029 33074 1484 33107
rect 13498 33107 13956 33108
rect 13498 33074 13953 33107
rect 7594 27865 7649 29187
rect 1235 20874 1579 20885
rect 1063 20852 1579 20874
rect 1454 20840 1579 20852
rect 13403 20882 13747 20885
rect 13772 20882 13959 20907
rect 13403 20852 13959 20882
rect 13403 20840 13528 20852
rect 1123 20792 1248 20814
rect 1234 20684 1248 20792
rect 1294 20792 1639 20825
rect 1294 20643 1308 20792
rect 1394 20780 1639 20792
rect 13343 20792 13688 20825
rect 13343 20780 13588 20792
rect 1675 20565 1719 20722
rect 1554 20560 1719 20565
rect 1387 20525 1719 20560
rect 1735 20565 1779 20662
rect 13203 20565 13247 20662
rect 1735 20532 1860 20565
rect 13122 20532 13247 20565
rect 13263 20565 13307 20722
rect 13642 20585 13688 20792
rect 13702 20792 13826 20822
rect 13702 20645 13748 20792
rect 13772 20657 13826 20792
rect 13832 20792 13899 20847
rect 13832 20750 13886 20792
rect 13832 20717 13899 20750
rect 13263 20560 13428 20565
rect 13263 20525 13595 20560
rect 1447 20465 1572 20500
rect 1554 20370 1572 20465
rect 1614 20472 1920 20505
rect 13062 20472 13368 20505
rect 1614 20465 1779 20472
rect 13203 20465 13368 20472
rect 1614 20323 1632 20465
rect 2000 20241 2039 20397
rect 1878 20232 2039 20241
rect 1715 20205 2039 20232
rect 2060 20241 2099 20337
rect 12883 20241 12922 20337
rect 2060 20207 2185 20241
rect 12797 20207 12922 20241
rect 12943 20241 12982 20397
rect 13350 20323 13368 20465
rect 13410 20465 13535 20500
rect 13410 20370 13428 20465
rect 12943 20232 13104 20241
rect 12943 20205 13267 20232
rect 1775 20145 1900 20172
rect 1878 20042 1900 20145
rect 1938 20147 2245 20181
rect 12737 20147 13044 20181
rect 1938 20145 2092 20147
rect 12890 20145 13044 20147
rect 1938 19982 1960 20145
rect 12072 19904 12118 19986
rect 2056 19883 2272 19891
rect 2056 19881 2301 19883
rect 12028 19856 12118 19904
rect 12132 19904 12178 20046
rect 13022 19982 13044 20145
rect 13082 20145 13207 20172
rect 13082 20042 13104 20145
rect 12132 19883 12544 19904
rect 12619 19891 12767 19904
rect 12619 19881 12926 19891
rect 2116 19821 2241 19831
rect 11968 19823 12707 19844
rect 11968 19796 12178 19823
rect 12559 19821 12707 19823
rect 11825 19547 11876 19706
rect 11885 19544 11936 19766
rect 12681 19641 12707 19821
rect 12741 19821 12866 19831
rect 12741 19701 12767 19821
rect 254 14007 320 18997
rect 15000 14007 15066 18997
rect 254 12837 320 13687
rect 15000 12837 15066 13687
rect 254 11667 320 12517
rect 15000 11667 15066 12517
rect 254 9547 320 11347
rect 15000 9547 15066 11347
rect 254 8337 320 9227
rect 15000 8337 15066 9227
rect 254 7368 320 8017
rect 15000 7368 15066 8017
rect 254 6397 320 7047
rect 15000 6397 15066 7047
rect 254 5187 320 6077
rect 15000 5187 15066 6077
rect 254 3977 320 4867
rect 15000 3977 15066 4867
rect 0 3007 320 3657
rect 14807 3007 15127 3657
rect 254 1797 320 2687
rect 15000 1797 15066 2687
rect 254 427 320 1477
rect 15000 427 15066 1477
<< metal3 >>
rect 5078 0 9858 391
<< metal4 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 19000
rect 14746 14007 15000 19000
rect 0 12817 254 13707
rect 14746 12817 15000 13707
rect 0 11647 254 12537
rect 14746 11647 15000 12537
rect 0 11281 254 11347
rect 14746 11281 15000 11347
rect 0 10625 254 11221
rect 14746 10625 15000 11221
rect 0 10329 254 10565
rect 14746 10329 15000 10565
rect 0 9673 254 10269
rect 14746 9673 15000 10269
rect 0 9547 254 9613
rect 14746 9547 15000 9613
rect 0 8317 254 9247
rect 14746 8317 15000 9247
rect 0 7347 254 8037
rect 14746 7347 15000 8037
rect 0 6377 254 7067
rect 14746 6377 15000 7067
rect 0 5167 254 6097
rect 14746 5167 15000 6097
rect 0 3957 254 4887
rect 14746 3957 15000 4887
rect 0 2987 193 3677
rect 14807 2987 15000 3677
rect 0 1777 254 2707
rect 14746 1777 15000 2707
rect 0 407 254 1497
rect 14746 407 15000 1497
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 7329 27865 7594 29187
rect 0 14007 254 18997
rect 14746 14007 15000 18997
rect 0 12837 254 13687
rect 14746 12837 15000 13687
rect 0 11667 254 12517
rect 14746 11667 15000 12517
rect 0 9547 254 11347
rect 14746 9547 15000 11347
rect 0 8337 254 9227
rect 14746 8337 15000 9227
rect 0 7368 254 8017
rect 14746 7368 15000 8017
rect 0 6397 254 7047
rect 14746 6397 15000 7047
rect 0 5187 254 6077
rect 14746 5187 15000 6077
rect 0 3977 254 4867
rect 14746 3977 15000 4867
rect 0 3007 193 3657
rect 14807 3007 15000 3657
rect 0 1797 254 2687
rect 14746 1797 15000 2687
rect 0 427 254 1477
rect 14746 427 15000 1477
use sky130_fd_io__simple_pad_and_busses  sky130_fd_io__simple_pad_and_busses_0
timestamp 1619240079
transform 1 0 -8 0 1 -1
box 8 1 14858 36278
<< labels >>
flabel metal3 s 5078 0 9858 391 0 FreeSans 3125 0 0 0 P_CORE
flabel metal4 s 0 7347 254 8037 3 FreeSans 812 0 0 0 VSSA
flabel metal4 s 0 11281 254 11347 3 FreeSans 812 0 0 0 VSSA
flabel metal4 s 0 9547 254 9613 3 FreeSans 812 0 0 0 VSSA
flabel metal4 s 0 10329 254 10565 3 FreeSans 812 0 0 0 VSSA
flabel metal4 s 14746 7347 15000 8037 3 FreeSans 812 180 0 0 VSSA
flabel metal4 s 14746 11281 15000 11347 3 FreeSans 812 180 0 0 VSSA
flabel metal4 s 14746 9547 15000 9613 3 FreeSans 812 180 0 0 VSSA
flabel metal4 s 14746 10329 15000 10565 3 FreeSans 812 180 0 0 VSSA
flabel metal5 s 14746 7368 15000 8017 3 FreeSans 812 180 0 0 VSSA
flabel metal5 s 0 9547 254 11347 3 FreeSans 812 0 0 0 VSSA
flabel metal5 s 0 7368 254 8017 3 FreeSans 812 0 0 0 VSSA
flabel metal5 s 14746 9547 15000 11347 3 FreeSans 812 180 0 0 VSSA
flabel metal4 s 0 8317 254 9247 3 FreeSans 812 0 0 0 VSSD
flabel metal4 s 14746 8317 15000 9247 3 FreeSans 812 180 0 0 VSSD
flabel metal5 s 0 8337 254 9227 3 FreeSans 812 0 0 0 VSSD
flabel metal5 s 14746 8337 15000 9227 3 FreeSans 812 180 0 0 VSSD
flabel metal4 s 0 9673 254 10269 3 FreeSans 812 0 0 0 AMUXBUS_B
flabel metal4 s 14746 9673 15000 10269 3 FreeSans 812 180 0 0 AMUXBUS_B
flabel metal4 s 0 10625 254 11221 3 FreeSans 812 0 0 0 AMUXBUS_A
flabel metal4 s 14746 10625 15000 11221 3 FreeSans 812 180 0 0 AMUXBUS_A
flabel metal4 s 0 12817 254 13707 3 FreeSans 812 0 0 0 VDDIO_Q
flabel metal4 s 14746 12817 15000 13707 3 FreeSans 812 180 0 0 VDDIO_Q
flabel metal5 s 14746 12837 15000 13687 3 FreeSans 812 180 0 0 VDDIO_Q
flabel metal5 s 0 12837 254 13687 3 FreeSans 812 0 0 0 VDDIO_Q
flabel metal4 s 0 14007 254 19000 3 FreeSans 812 0 0 0 VDDIO
flabel metal4 s 0 3957 254 4887 3 FreeSans 812 0 0 0 VDDIO
flabel metal4 s 14746 14007 15000 19000 3 FreeSans 812 180 0 0 VDDIO
flabel metal4 s 14746 3957 15000 4887 3 FreeSans 812 180 0 0 VDDIO
flabel metal5 s 0 3977 254 4867 3 FreeSans 812 0 0 0 VDDIO
flabel metal5 s 0 14007 254 18997 3 FreeSans 812 0 0 0 VDDIO
flabel metal5 s 14746 3977 15000 4867 3 FreeSans 812 180 0 0 VDDIO
flabel metal5 s 14746 14007 15000 18997 3 FreeSans 812 180 0 0 VDDIO
flabel metal4 s 0 6377 254 7067 3 FreeSans 812 0 0 0 VSWITCH
flabel metal4 s 14746 6377 15000 7067 3 FreeSans 812 180 0 0 VSWITCH
flabel metal5 s 14746 6397 15000 7047 3 FreeSans 812 180 0 0 VSWITCH
flabel metal5 s 0 6397 254 7047 3 FreeSans 812 0 0 0 VSWITCH
flabel metal4 s 0 5167 254 6097 3 FreeSans 812 0 0 0 VSSIO
flabel metal4 s 14746 5167 15000 6097 3 FreeSans 812 180 0 0 VSSIO
flabel metal4 s 0 35157 254 40000 3 FreeSans 812 0 0 0 VSSIO
flabel metal4 s 127 38321 127 38321 3 FreeSans 812 0 0 0 VSSIO
flabel metal4 s 14746 35157 15000 40000 3 FreeSans 812 180 0 0 VSSIO
flabel metal4 s 14873 38321 14873 38321 3 FreeSans 812 180 0 0 VSSIO
flabel metal5 s 14746 5187 15000 6077 3 FreeSans 812 180 0 0 VSSIO
flabel metal5 s 14746 35157 15000 40000 3 FreeSans 812 180 0 0 VSSIO
flabel metal5 s 0 35157 254 40000 3 FreeSans 812 0 0 0 VSSIO
flabel metal5 s 0 5187 254 6077 3 FreeSans 812 0 0 0 VSSIO
flabel metal4 s 0 2987 193 3677 3 FreeSans 812 0 0 0 VDDA
flabel metal4 s 14807 2987 15000 3677 3 FreeSans 812 180 0 0 VDDA
flabel metal5 s 0 3007 193 3657 3 FreeSans 812 0 0 0 VDDA
flabel metal5 s 14807 3007 15000 3657 3 FreeSans 812 180 0 0 VDDA
flabel metal4 s 0 1777 254 2707 3 FreeSans 812 0 0 0 VCCD
flabel metal4 s 14746 1777 15000 2707 3 FreeSans 812 180 0 0 VCCD
flabel metal5 s 0 1797 254 2687 3 FreeSans 812 0 0 0 VCCD
flabel metal5 s 14746 1797 15000 2687 3 FreeSans 812 180 0 0 VCCD
flabel metal4 s 0 407 254 1497 3 FreeSans 812 0 0 0 VCCHIB
flabel metal4 s 14746 407 15000 1497 3 FreeSans 812 180 0 0 VCCHIB
flabel metal5 s 0 427 254 1477 3 FreeSans 812 0 0 0 VCCHIB
flabel metal5 s 14746 427 15000 1477 3 FreeSans 812 180 0 0 VCCHIB
flabel metal4 s 0 11647 254 12537 3 FreeSans 812 0 0 0 VSSIO_Q
flabel metal4 s 14746 11647 15000 12537 3 FreeSans 812 180 0 0 VSSIO_Q
flabel metal5 s 14746 11667 15000 12517 3 FreeSans 812 180 0 0 VSSIO_Q
flabel metal5 s 0 11667 254 12517 3 FreeSans 812 0 0 0 VSSIO_Q
flabel metal5 s 7329 27865 7594 29187 0 FreeSans 3125 0 0 0 P_PAD
<< end >>
