magic
tech sky130A
magscale 1 2
timestamp 1619862920
<< checkpaint >>
rect -3455 -3444 18488 40846
<< metal1 >>
rect 15240 14945 17187 15070
rect 15240 9453 15341 14945
rect 17057 9453 17187 14945
rect 15240 7473 17187 9453
rect 15240 5437 15324 7473
rect 17104 5437 17187 7473
rect 5101 -7 5685 83
rect 4185 -163 11313 -7
rect 15240 -163 17187 5437
rect 4185 -1384 17187 -163
rect 4185 -2184 16387 -1384
tri 16387 -2184 17187 -1384 nw
<< via1 >>
rect 15341 9453 17057 14945
rect 15324 5437 17104 7473
<< metal2 >>
rect 15240 39515 17187 39586
rect 15240 34819 15307 39515
rect 17123 34819 17187 39515
rect 15240 14945 17187 34819
rect 15240 9453 15341 14945
rect 17057 9453 17187 14945
rect 15240 9312 17187 9453
rect -2195 8794 100 8833
rect -2195 7938 -2136 8794
rect -240 7938 100 8794
rect -2195 7903 100 7938
rect 14940 8802 17228 8840
rect 14940 7946 15165 8802
rect 16181 7946 17228 8802
rect 14940 7910 17228 7946
rect 15240 7473 17187 7560
rect 15240 5613 15324 7473
rect 17104 5613 17187 7473
rect 15240 4837 15298 5613
rect 17114 4837 17187 5613
rect 15240 4678 17187 4837
<< via2 >>
rect 15307 34819 17123 39515
rect -2136 7938 -240 8794
rect 15165 7946 16181 8802
rect 15298 5437 15324 5613
rect 15324 5437 17104 5613
rect 17104 5437 17114 5613
rect 15298 4837 17114 5437
<< metal3 >>
rect 15240 39519 17187 39586
rect 15240 34815 15303 39519
rect 17127 34815 17187 39519
rect 15240 34743 17187 34815
rect -2195 8797 -179 8833
rect -2195 7933 -2141 8797
rect -237 7933 -179 8797
rect -2195 7903 -179 7933
rect 15121 8806 17228 8840
rect 15121 8802 15181 8806
rect 15121 7946 15165 8802
rect 15121 7942 15181 7946
rect 17165 7942 17228 8806
rect 15121 7910 17228 7942
rect 15240 5617 17187 5683
rect 15240 4833 15294 5617
rect 17118 4833 17187 5617
rect 15240 4753 17187 4833
rect 5228 2223 7341 2269
rect 5228 1439 5252 2223
rect 7316 1439 7341 2223
rect 5228 1394 7341 1439
rect 7705 2221 9818 2267
rect 7705 1437 7729 2221
rect 9793 1437 9818 2221
rect 7705 1392 9818 1437
<< via3 >>
rect 15303 39515 17127 39519
rect 15303 34819 15307 39515
rect 15307 34819 17123 39515
rect 17123 34819 17127 39515
rect 15303 34815 17127 34819
rect -2141 8794 -237 8797
rect -2141 7938 -2136 8794
rect -2136 7938 -240 8794
rect -240 7938 -237 8794
rect -2141 7933 -237 7938
rect 15181 8802 17165 8806
rect 15181 7946 16181 8802
rect 16181 7946 17165 8802
rect 15181 7942 17165 7946
rect 15294 5613 17118 5617
rect 15294 4837 15298 5613
rect 15298 4837 17114 5613
rect 17114 4837 17118 5613
rect 15294 4833 17118 4837
rect 5252 1439 7316 2223
rect 7729 1437 9793 2221
<< metal4 >>
rect 14957 39519 17187 39586
rect 14957 34815 15303 39519
rect 17127 34815 17187 39519
rect 14957 34743 17187 34815
rect -2195 8797 14 8833
rect -2195 7933 -2141 8797
rect -237 7933 14 8797
rect -2195 7903 14 7933
rect 14940 8806 17228 8840
rect 14940 7942 15181 8806
rect 17165 7942 17228 8806
rect 14940 7910 17228 7942
rect 14987 5617 17187 5683
rect 14987 4833 15294 5617
rect 17118 4833 17187 5617
rect 14987 4753 17187 4833
rect 5228 2223 7341 2269
rect 5228 1439 5252 2223
rect 7316 1439 7341 2223
rect 5228 1394 7341 1439
rect 7705 2221 9818 2267
rect 7705 1437 7729 2221
rect 9793 1437 9818 2221
rect 7705 1392 9818 1437
<< properties >>
string FIXED_BBOX 0 -7 15000 39593
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_END 1204620
string GDS_START 700240
<< end >>
