magic
tech sky130A
magscale 1 2
timestamp 1619862920
<< checkpaint >>
rect -1288 -1260 1408 1731
use sky130_fd_pr__hvdfl1sd__example_5595914180851  sky130_fd_pr__hvdfl1sd__example_5595914180851_0
timestamp 1619862920
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_5595914180851  sky130_fd_pr__hvdfl1sd__example_5595914180851_1
timestamp 1619862920
transform 1 0 120 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 148 471 148 471 0 FreeSans 300 0 0 0 D
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 3520886
string GDS_START 3519960
<< end >>
