module phase_interpolator (
    input [3:0] l_con,
    input [3:0] r_con,
    output pasheout
);
    
// Buffer to avoid load the osc core overly



endmodule