magic
tech sky130A
magscale 1 2
timestamp 1619862920
<< checkpaint >>
rect 3035 -7162 28233 18845
<< dnwell >>
rect 4795 4227 6256 11135
<< nwell >>
rect 4710 10929 6283 11231
rect 4710 4433 5012 10929
rect 4710 4131 6283 4433
<< pwell >>
rect 5072 10715 5850 10869
rect 5072 4668 5226 10715
rect 5696 4668 5850 10715
rect 5072 4514 5850 4668
<< psubdiff >>
rect 5098 4927 5200 4956
rect 5098 4655 5200 4689
rect 5132 4642 5200 4655
rect 5132 4621 5166 4642
rect 5098 4540 5166 4621
rect 5676 4608 5722 4642
rect 5676 4574 5824 4608
rect 5676 4540 5710 4574
rect 5744 4540 5824 4574
<< mvpsubdiff >>
rect 5098 10809 5174 10843
rect 5208 10809 5314 10843
rect 5098 10775 5314 10809
rect 5200 10741 5314 10775
rect 5756 10762 5824 10843
rect 5756 10741 5790 10762
rect 5722 10728 5790 10741
rect 5722 10694 5824 10728
rect 5098 4956 5200 4961
<< mvnsubdiff >>
rect 4776 11097 4844 11165
rect 4810 11063 4844 11097
rect 5286 11131 5321 11165
rect 5355 11131 5390 11165
rect 5424 11131 5459 11165
rect 5493 11131 5528 11165
rect 5562 11131 5597 11165
rect 5631 11131 5666 11165
rect 5700 11131 5735 11165
rect 5769 11131 5804 11165
rect 5838 11131 5873 11165
rect 5907 11131 5942 11165
rect 5976 11131 6011 11165
rect 6045 11131 6080 11165
rect 6114 11131 6149 11165
rect 6183 11131 6217 11165
rect 5286 11097 6217 11131
rect 5286 11063 5321 11097
rect 5355 11063 5390 11097
rect 5424 11063 5459 11097
rect 5493 11063 5528 11097
rect 5562 11063 5597 11097
rect 5631 11063 5666 11097
rect 5700 11063 5735 11097
rect 5769 11063 5804 11097
rect 5838 11063 5873 11097
rect 5907 11063 5942 11097
rect 5976 11063 6011 11097
rect 6045 11063 6080 11097
rect 6114 11063 6149 11097
rect 6183 11063 6217 11097
rect 4776 11028 4912 11063
rect 4810 10994 4844 11028
rect 4878 10995 4912 11028
rect 5286 11029 6217 11063
rect 5286 10995 5321 11029
rect 5355 10995 5390 11029
rect 5424 10995 5459 11029
rect 5493 10995 5528 11029
rect 5562 10995 5597 11029
rect 5631 10995 5666 11029
rect 5700 10995 5735 11029
rect 5769 10995 5804 11029
rect 5838 10995 5873 11029
rect 5907 10995 5942 11029
rect 5976 10995 6011 11029
rect 6045 10995 6080 11029
rect 6114 10995 6149 11029
rect 6183 10995 6217 11029
rect 4878 10994 4946 10995
rect 4776 10960 4946 10994
rect 4776 10959 4912 10960
rect 4810 10925 4844 10959
rect 4878 10926 4912 10959
rect 4878 10925 4946 10926
rect 4776 10891 4946 10925
rect 4776 10890 4912 10891
rect 4810 10856 4844 10890
rect 4878 10857 4912 10890
rect 4878 10856 4946 10857
rect 4776 10822 4946 10856
rect 4776 10821 4912 10822
rect 4810 10787 4844 10821
rect 4878 10788 4912 10821
rect 4878 10787 4946 10788
rect 4776 10753 4946 10787
rect 4776 10752 4912 10753
rect 4810 10718 4844 10752
rect 4878 10719 4912 10752
rect 4878 10718 4946 10719
rect 4776 10684 4946 10718
rect 4776 10683 4912 10684
rect 4810 10649 4844 10683
rect 4878 10650 4912 10683
rect 4878 10649 4946 10650
rect 4776 10615 4946 10649
rect 4776 10614 4912 10615
rect 4810 10580 4844 10614
rect 4878 10581 4912 10614
rect 4878 10580 4946 10581
rect 4776 10546 4946 10580
rect 4776 10545 4912 10546
rect 4810 10511 4844 10545
rect 4878 10512 4912 10545
rect 4878 10511 4946 10512
rect 4776 10477 4946 10511
rect 4776 10476 4912 10477
rect 4810 10442 4844 10476
rect 4878 10443 4912 10476
rect 4878 10442 4946 10443
rect 4776 10408 4946 10442
rect 4776 10407 4912 10408
rect 4810 10373 4844 10407
rect 4878 10374 4912 10407
rect 4878 10373 4946 10374
rect 4776 10339 4946 10373
rect 4776 10338 4912 10339
rect 4810 10304 4844 10338
rect 4878 10305 4912 10338
rect 4878 10304 4946 10305
rect 4776 10270 4946 10304
rect 4776 10269 4912 10270
rect 4810 10235 4844 10269
rect 4878 10236 4912 10269
rect 4878 10235 4946 10236
rect 4776 10201 4946 10235
rect 4776 10200 4912 10201
rect 4810 10166 4844 10200
rect 4878 10167 4912 10200
rect 4878 10166 4946 10167
rect 4776 10132 4946 10166
rect 4776 10131 4912 10132
rect 4810 10097 4844 10131
rect 4878 10098 4912 10131
rect 4878 10097 4946 10098
rect 4776 10063 4946 10097
rect 4776 10062 4912 10063
rect 4810 10028 4844 10062
rect 4878 10029 4912 10062
rect 4878 10028 4946 10029
rect 4776 9994 4946 10028
rect 4776 9993 4912 9994
rect 4810 9959 4844 9993
rect 4878 9960 4912 9993
rect 4878 9959 4946 9960
rect 4776 9925 4946 9959
rect 4776 9924 4912 9925
rect 4810 9890 4844 9924
rect 4878 9891 4912 9924
rect 4878 9890 4946 9891
rect 4776 9856 4946 9890
rect 4776 9855 4912 9856
rect 4810 9821 4844 9855
rect 4878 9822 4912 9855
rect 4878 9821 4946 9822
rect 4776 9787 4946 9821
rect 4776 9786 4912 9787
rect 4810 9752 4844 9786
rect 4878 9753 4912 9786
rect 4878 9752 4946 9753
rect 4776 9718 4946 9752
rect 4776 9717 4912 9718
rect 4810 9683 4844 9717
rect 4878 9684 4912 9717
rect 4878 9683 4946 9684
rect 4776 9649 4946 9683
rect 4776 9648 4912 9649
rect 4810 9614 4844 9648
rect 4878 9615 4912 9648
rect 4878 9614 4946 9615
rect 4776 9580 4946 9614
rect 4776 9579 4912 9580
rect 4810 9545 4844 9579
rect 4878 9546 4912 9579
rect 4878 9545 4946 9546
rect 4776 9511 4946 9545
rect 4776 9510 4912 9511
rect 4810 9476 4844 9510
rect 4878 9477 4912 9510
rect 4878 9476 4946 9477
rect 4776 9442 4946 9476
rect 4776 9441 4912 9442
rect 4810 9407 4844 9441
rect 4878 9408 4912 9441
rect 4878 9407 4946 9408
rect 4776 9373 4946 9407
rect 4776 9372 4912 9373
rect 4810 9338 4844 9372
rect 4878 9339 4912 9372
rect 4878 9338 4946 9339
rect 4776 9304 4946 9338
rect 4776 9303 4912 9304
rect 4810 9269 4844 9303
rect 4878 9270 4912 9303
rect 4878 9269 4946 9270
rect 4776 9235 4946 9269
rect 4776 9234 4912 9235
rect 4810 9200 4844 9234
rect 4878 9201 4912 9234
rect 4878 9200 4946 9201
rect 4776 9166 4946 9200
rect 4776 9165 4912 9166
rect 4810 9131 4844 9165
rect 4878 9132 4912 9165
rect 4878 9131 4946 9132
rect 4776 9097 4946 9131
rect 4776 9096 4912 9097
rect 4810 9062 4844 9096
rect 4878 9063 4912 9096
rect 4878 9062 4946 9063
rect 4776 9028 4946 9062
rect 4776 9027 4912 9028
rect 4810 8993 4844 9027
rect 4878 8994 4912 9027
rect 4878 8993 4946 8994
rect 4776 8959 4946 8993
rect 4776 8958 4912 8959
rect 4810 8924 4844 8958
rect 4878 8925 4912 8958
rect 4878 8924 4946 8925
rect 4776 8890 4946 8924
rect 4776 8889 4912 8890
rect 4810 8855 4844 8889
rect 4878 8856 4912 8889
rect 4878 8855 4946 8856
rect 4776 8821 4946 8855
rect 4776 8820 4912 8821
rect 4810 8786 4844 8820
rect 4878 8787 4912 8820
rect 4878 8786 4946 8787
rect 4776 8752 4946 8786
rect 4776 8751 4912 8752
rect 4810 8717 4844 8751
rect 4878 8718 4912 8751
rect 4878 8717 4946 8718
rect 4776 8683 4946 8717
rect 4776 8682 4912 8683
rect 4810 8648 4844 8682
rect 4878 8649 4912 8682
rect 4878 8648 4946 8649
rect 4776 8614 4946 8648
rect 4776 8613 4912 8614
rect 4810 8579 4844 8613
rect 4878 8580 4912 8613
rect 4878 8579 4946 8580
rect 4776 8545 4946 8579
rect 4776 8544 4912 8545
rect 4810 8510 4844 8544
rect 4878 8511 4912 8544
rect 4878 8510 4946 8511
rect 4776 8476 4946 8510
rect 4776 8475 4912 8476
rect 4810 8441 4844 8475
rect 4878 8442 4912 8475
rect 4878 8441 4946 8442
rect 4776 8407 4946 8441
rect 4776 8406 4912 8407
rect 4810 8372 4844 8406
rect 4878 8373 4912 8406
rect 4878 8372 4946 8373
rect 4776 8338 4946 8372
rect 4776 8337 4912 8338
rect 4810 8303 4844 8337
rect 4878 8304 4912 8337
rect 4878 8303 4946 8304
rect 4776 8269 4946 8303
rect 4776 8268 4912 8269
rect 4810 8234 4844 8268
rect 4878 8235 4912 8268
rect 4878 8234 4946 8235
rect 4776 8200 4946 8234
rect 4776 8199 4912 8200
rect 4810 8165 4844 8199
rect 4878 8166 4912 8199
rect 4878 8165 4946 8166
rect 4776 8131 4946 8165
rect 4776 8130 4912 8131
rect 4810 8096 4844 8130
rect 4878 8097 4912 8130
rect 4878 8096 4946 8097
rect 4776 8062 4946 8096
rect 4776 8061 4912 8062
rect 4810 8027 4844 8061
rect 4878 8028 4912 8061
rect 4878 8027 4946 8028
rect 4776 7993 4946 8027
rect 4776 7992 4912 7993
rect 4810 7958 4844 7992
rect 4878 7959 4912 7992
rect 4878 7958 4946 7959
rect 4776 7924 4946 7958
rect 4776 7923 4912 7924
rect 4810 7889 4844 7923
rect 4878 7890 4912 7923
rect 4878 7889 4946 7890
rect 4776 7855 4946 7889
rect 4776 7854 4912 7855
rect 4810 7820 4844 7854
rect 4878 7821 4912 7854
rect 4878 7820 4946 7821
rect 4776 7786 4946 7820
rect 4776 7785 4912 7786
rect 4810 7751 4844 7785
rect 4878 7752 4912 7785
rect 4878 7751 4946 7752
rect 4776 7717 4946 7751
rect 4776 7716 4912 7717
rect 4810 7682 4844 7716
rect 4878 7683 4912 7716
rect 4878 7682 4946 7683
rect 4776 7648 4946 7682
rect 4776 7647 4912 7648
rect 4810 7613 4844 7647
rect 4878 7614 4912 7647
rect 4878 7613 4946 7614
rect 4776 7579 4946 7613
rect 4776 7578 4912 7579
rect 4810 7544 4844 7578
rect 4878 7545 4912 7578
rect 4878 7544 4946 7545
rect 4776 7510 4946 7544
rect 4776 7509 4912 7510
rect 4810 7475 4844 7509
rect 4878 7476 4912 7509
rect 4878 7475 4946 7476
rect 4776 7441 4946 7475
rect 4776 7440 4912 7441
rect 4810 7406 4844 7440
rect 4878 7407 4912 7440
rect 4878 7406 4946 7407
rect 4776 7372 4946 7406
rect 4776 7371 4912 7372
rect 4810 7337 4844 7371
rect 4878 7338 4912 7371
rect 4878 7337 4946 7338
rect 4776 7303 4946 7337
rect 4776 7302 4912 7303
rect 4810 7268 4844 7302
rect 4878 7269 4912 7302
rect 4878 7268 4946 7269
rect 4776 7234 4946 7268
rect 4776 7233 4912 7234
rect 4810 7199 4844 7233
rect 4878 7200 4912 7233
rect 4878 7199 4946 7200
rect 4776 7165 4946 7199
rect 4776 7164 4912 7165
rect 4810 7130 4844 7164
rect 4878 7131 4912 7164
rect 4878 7130 4946 7131
rect 4776 7096 4946 7130
rect 4776 7095 4912 7096
rect 4810 7061 4844 7095
rect 4878 7062 4912 7095
rect 4878 7061 4946 7062
rect 4776 7027 4946 7061
rect 4776 7026 4912 7027
rect 4810 6992 4844 7026
rect 4878 6993 4912 7026
rect 4878 6992 4946 6993
rect 4776 6958 4946 6992
rect 4776 6957 4912 6958
rect 4810 6923 4844 6957
rect 4878 6924 4912 6957
rect 4878 6923 4946 6924
rect 4776 6889 4946 6923
rect 4776 6888 4912 6889
rect 4810 6854 4844 6888
rect 4878 6855 4912 6888
rect 4878 6854 4946 6855
rect 4776 6820 4946 6854
rect 4776 6819 4912 6820
rect 4810 6785 4844 6819
rect 4878 6786 4912 6819
rect 4878 6785 4946 6786
rect 4776 6751 4946 6785
rect 4776 6750 4912 6751
rect 4810 6716 4844 6750
rect 4878 6717 4912 6750
rect 4878 6716 4946 6717
rect 4776 6682 4946 6716
rect 4776 6681 4912 6682
rect 4810 6647 4844 6681
rect 4878 6648 4912 6681
rect 4878 6647 4946 6648
rect 4776 6613 4946 6647
rect 4776 6612 4912 6613
rect 4810 6578 4844 6612
rect 4878 6579 4912 6612
rect 4878 6578 4946 6579
rect 4776 6544 4946 6578
rect 4776 6543 4912 6544
rect 4878 6510 4912 6543
rect 4878 6475 4946 6510
rect 4946 4333 4981 4367
rect 5015 4333 5050 4367
rect 5084 4333 5119 4367
rect 5153 4333 5188 4367
rect 5222 4333 5257 4367
rect 5291 4333 5326 4367
rect 5360 4333 5395 4367
rect 5429 4333 5464 4367
rect 5498 4333 5533 4367
rect 5567 4333 5602 4367
rect 5636 4333 5671 4367
rect 5705 4333 5740 4367
rect 5774 4333 5809 4367
rect 4878 4299 5809 4333
rect 4878 4265 4913 4299
rect 4947 4265 4982 4299
rect 5016 4265 5051 4299
rect 5085 4265 5120 4299
rect 5154 4265 5189 4299
rect 5223 4265 5258 4299
rect 5292 4265 5327 4299
rect 5361 4265 5396 4299
rect 5430 4265 5465 4299
rect 5499 4265 5534 4299
rect 5568 4265 5603 4299
rect 5637 4265 5672 4299
rect 5706 4265 5741 4299
rect 4776 4231 5741 4265
rect 4776 4197 4844 4231
rect 4878 4197 4913 4231
rect 4947 4197 4982 4231
rect 5016 4197 5051 4231
rect 5085 4197 5120 4231
rect 5154 4197 5189 4231
rect 5223 4197 5258 4231
rect 5292 4197 5327 4231
rect 5361 4197 5396 4231
rect 5430 4197 5465 4231
rect 5499 4197 5534 4231
rect 5568 4197 5603 4231
rect 5637 4197 5672 4231
rect 5706 4197 5741 4231
rect 6183 4197 6217 4367
<< psubdiffcont >>
rect 5098 4689 5200 4927
rect 5098 4621 5132 4655
rect 5166 4540 5676 4642
rect 5722 4608 5824 4956
rect 5710 4540 5744 4574
<< mvpsubdiffcont >>
rect 5174 10809 5208 10843
rect 5098 4961 5200 10775
rect 5314 10741 5756 10843
rect 5790 10728 5824 10762
rect 5722 4956 5824 10694
<< mvnsubdiffcont >>
rect 4776 11063 4810 11097
rect 4844 11063 5286 11165
rect 5321 11131 5355 11165
rect 5390 11131 5424 11165
rect 5459 11131 5493 11165
rect 5528 11131 5562 11165
rect 5597 11131 5631 11165
rect 5666 11131 5700 11165
rect 5735 11131 5769 11165
rect 5804 11131 5838 11165
rect 5873 11131 5907 11165
rect 5942 11131 5976 11165
rect 6011 11131 6045 11165
rect 6080 11131 6114 11165
rect 6149 11131 6183 11165
rect 5321 11063 5355 11097
rect 5390 11063 5424 11097
rect 5459 11063 5493 11097
rect 5528 11063 5562 11097
rect 5597 11063 5631 11097
rect 5666 11063 5700 11097
rect 5735 11063 5769 11097
rect 5804 11063 5838 11097
rect 5873 11063 5907 11097
rect 5942 11063 5976 11097
rect 6011 11063 6045 11097
rect 6080 11063 6114 11097
rect 6149 11063 6183 11097
rect 4776 10994 4810 11028
rect 4844 10994 4878 11028
rect 4912 10995 5286 11063
rect 5321 10995 5355 11029
rect 5390 10995 5424 11029
rect 5459 10995 5493 11029
rect 5528 10995 5562 11029
rect 5597 10995 5631 11029
rect 5666 10995 5700 11029
rect 5735 10995 5769 11029
rect 5804 10995 5838 11029
rect 5873 10995 5907 11029
rect 5942 10995 5976 11029
rect 6011 10995 6045 11029
rect 6080 10995 6114 11029
rect 6149 10995 6183 11029
rect 4776 10925 4810 10959
rect 4844 10925 4878 10959
rect 4912 10926 4946 10960
rect 4776 10856 4810 10890
rect 4844 10856 4878 10890
rect 4912 10857 4946 10891
rect 4776 10787 4810 10821
rect 4844 10787 4878 10821
rect 4912 10788 4946 10822
rect 4776 10718 4810 10752
rect 4844 10718 4878 10752
rect 4912 10719 4946 10753
rect 4776 10649 4810 10683
rect 4844 10649 4878 10683
rect 4912 10650 4946 10684
rect 4776 10580 4810 10614
rect 4844 10580 4878 10614
rect 4912 10581 4946 10615
rect 4776 10511 4810 10545
rect 4844 10511 4878 10545
rect 4912 10512 4946 10546
rect 4776 10442 4810 10476
rect 4844 10442 4878 10476
rect 4912 10443 4946 10477
rect 4776 10373 4810 10407
rect 4844 10373 4878 10407
rect 4912 10374 4946 10408
rect 4776 10304 4810 10338
rect 4844 10304 4878 10338
rect 4912 10305 4946 10339
rect 4776 10235 4810 10269
rect 4844 10235 4878 10269
rect 4912 10236 4946 10270
rect 4776 10166 4810 10200
rect 4844 10166 4878 10200
rect 4912 10167 4946 10201
rect 4776 10097 4810 10131
rect 4844 10097 4878 10131
rect 4912 10098 4946 10132
rect 4776 10028 4810 10062
rect 4844 10028 4878 10062
rect 4912 10029 4946 10063
rect 4776 9959 4810 9993
rect 4844 9959 4878 9993
rect 4912 9960 4946 9994
rect 4776 9890 4810 9924
rect 4844 9890 4878 9924
rect 4912 9891 4946 9925
rect 4776 9821 4810 9855
rect 4844 9821 4878 9855
rect 4912 9822 4946 9856
rect 4776 9752 4810 9786
rect 4844 9752 4878 9786
rect 4912 9753 4946 9787
rect 4776 9683 4810 9717
rect 4844 9683 4878 9717
rect 4912 9684 4946 9718
rect 4776 9614 4810 9648
rect 4844 9614 4878 9648
rect 4912 9615 4946 9649
rect 4776 9545 4810 9579
rect 4844 9545 4878 9579
rect 4912 9546 4946 9580
rect 4776 9476 4810 9510
rect 4844 9476 4878 9510
rect 4912 9477 4946 9511
rect 4776 9407 4810 9441
rect 4844 9407 4878 9441
rect 4912 9408 4946 9442
rect 4776 9338 4810 9372
rect 4844 9338 4878 9372
rect 4912 9339 4946 9373
rect 4776 9269 4810 9303
rect 4844 9269 4878 9303
rect 4912 9270 4946 9304
rect 4776 9200 4810 9234
rect 4844 9200 4878 9234
rect 4912 9201 4946 9235
rect 4776 9131 4810 9165
rect 4844 9131 4878 9165
rect 4912 9132 4946 9166
rect 4776 9062 4810 9096
rect 4844 9062 4878 9096
rect 4912 9063 4946 9097
rect 4776 8993 4810 9027
rect 4844 8993 4878 9027
rect 4912 8994 4946 9028
rect 4776 8924 4810 8958
rect 4844 8924 4878 8958
rect 4912 8925 4946 8959
rect 4776 8855 4810 8889
rect 4844 8855 4878 8889
rect 4912 8856 4946 8890
rect 4776 8786 4810 8820
rect 4844 8786 4878 8820
rect 4912 8787 4946 8821
rect 4776 8717 4810 8751
rect 4844 8717 4878 8751
rect 4912 8718 4946 8752
rect 4776 8648 4810 8682
rect 4844 8648 4878 8682
rect 4912 8649 4946 8683
rect 4776 8579 4810 8613
rect 4844 8579 4878 8613
rect 4912 8580 4946 8614
rect 4776 8510 4810 8544
rect 4844 8510 4878 8544
rect 4912 8511 4946 8545
rect 4776 8441 4810 8475
rect 4844 8441 4878 8475
rect 4912 8442 4946 8476
rect 4776 8372 4810 8406
rect 4844 8372 4878 8406
rect 4912 8373 4946 8407
rect 4776 8303 4810 8337
rect 4844 8303 4878 8337
rect 4912 8304 4946 8338
rect 4776 8234 4810 8268
rect 4844 8234 4878 8268
rect 4912 8235 4946 8269
rect 4776 8165 4810 8199
rect 4844 8165 4878 8199
rect 4912 8166 4946 8200
rect 4776 8096 4810 8130
rect 4844 8096 4878 8130
rect 4912 8097 4946 8131
rect 4776 8027 4810 8061
rect 4844 8027 4878 8061
rect 4912 8028 4946 8062
rect 4776 7958 4810 7992
rect 4844 7958 4878 7992
rect 4912 7959 4946 7993
rect 4776 7889 4810 7923
rect 4844 7889 4878 7923
rect 4912 7890 4946 7924
rect 4776 7820 4810 7854
rect 4844 7820 4878 7854
rect 4912 7821 4946 7855
rect 4776 7751 4810 7785
rect 4844 7751 4878 7785
rect 4912 7752 4946 7786
rect 4776 7682 4810 7716
rect 4844 7682 4878 7716
rect 4912 7683 4946 7717
rect 4776 7613 4810 7647
rect 4844 7613 4878 7647
rect 4912 7614 4946 7648
rect 4776 7544 4810 7578
rect 4844 7544 4878 7578
rect 4912 7545 4946 7579
rect 4776 7475 4810 7509
rect 4844 7475 4878 7509
rect 4912 7476 4946 7510
rect 4776 7406 4810 7440
rect 4844 7406 4878 7440
rect 4912 7407 4946 7441
rect 4776 7337 4810 7371
rect 4844 7337 4878 7371
rect 4912 7338 4946 7372
rect 4776 7268 4810 7302
rect 4844 7268 4878 7302
rect 4912 7269 4946 7303
rect 4776 7199 4810 7233
rect 4844 7199 4878 7233
rect 4912 7200 4946 7234
rect 4776 7130 4810 7164
rect 4844 7130 4878 7164
rect 4912 7131 4946 7165
rect 4776 7061 4810 7095
rect 4844 7061 4878 7095
rect 4912 7062 4946 7096
rect 4776 6992 4810 7026
rect 4844 6992 4878 7026
rect 4912 6993 4946 7027
rect 4776 6923 4810 6957
rect 4844 6923 4878 6957
rect 4912 6924 4946 6958
rect 4776 6854 4810 6888
rect 4844 6854 4878 6888
rect 4912 6855 4946 6889
rect 4776 6785 4810 6819
rect 4844 6785 4878 6819
rect 4912 6786 4946 6820
rect 4776 6716 4810 6750
rect 4844 6716 4878 6750
rect 4912 6717 4946 6751
rect 4776 6647 4810 6681
rect 4844 6647 4878 6681
rect 4912 6648 4946 6682
rect 4776 6578 4810 6612
rect 4844 6578 4878 6612
rect 4912 6579 4946 6613
rect 4776 6475 4878 6543
rect 4912 6510 4946 6544
rect 4776 4333 4946 6475
rect 4981 4333 5015 4367
rect 5050 4333 5084 4367
rect 5119 4333 5153 4367
rect 5188 4333 5222 4367
rect 5257 4333 5291 4367
rect 5326 4333 5360 4367
rect 5395 4333 5429 4367
rect 5464 4333 5498 4367
rect 5533 4333 5567 4367
rect 5602 4333 5636 4367
rect 5671 4333 5705 4367
rect 5740 4333 5774 4367
rect 4776 4265 4878 4333
rect 5809 4299 6183 4367
rect 4913 4265 4947 4299
rect 4982 4265 5016 4299
rect 5051 4265 5085 4299
rect 5120 4265 5154 4299
rect 5189 4265 5223 4299
rect 5258 4265 5292 4299
rect 5327 4265 5361 4299
rect 5396 4265 5430 4299
rect 5465 4265 5499 4299
rect 5534 4265 5568 4299
rect 5603 4265 5637 4299
rect 5672 4265 5706 4299
rect 4844 4197 4878 4231
rect 4913 4197 4947 4231
rect 4982 4197 5016 4231
rect 5051 4197 5085 4231
rect 5120 4197 5154 4231
rect 5189 4197 5223 4231
rect 5258 4197 5292 4231
rect 5327 4197 5361 4231
rect 5396 4197 5430 4231
rect 5465 4197 5499 4231
rect 5534 4197 5568 4231
rect 5603 4197 5637 4231
rect 5672 4197 5706 4231
rect 5741 4197 6183 4299
<< poly >>
rect 5282 10582 5433 10605
rect 5282 10548 5298 10582
rect 5332 10548 5366 10582
rect 5400 10548 5433 10582
rect 5282 10525 5433 10548
rect 5489 10582 5640 10605
rect 5489 10548 5522 10582
rect 5556 10548 5590 10582
rect 5624 10548 5640 10582
rect 5489 10525 5640 10548
rect 5282 9850 5433 9873
rect 5282 9816 5298 9850
rect 5332 9816 5366 9850
rect 5400 9816 5433 9850
rect 5282 9793 5433 9816
rect 5489 9850 5640 9873
rect 5489 9816 5522 9850
rect 5556 9816 5590 9850
rect 5624 9816 5640 9850
rect 5489 9793 5640 9816
rect 5282 9118 5433 9141
rect 5282 9084 5298 9118
rect 5332 9084 5366 9118
rect 5400 9084 5433 9118
rect 5282 9061 5433 9084
rect 5489 9118 5640 9141
rect 5489 9084 5522 9118
rect 5556 9084 5590 9118
rect 5624 9084 5640 9118
rect 5489 9061 5640 9084
rect 5282 8386 5433 8409
rect 5282 8352 5298 8386
rect 5332 8352 5366 8386
rect 5400 8352 5433 8386
rect 5282 8329 5433 8352
rect 5489 8386 5640 8409
rect 5489 8352 5522 8386
rect 5556 8352 5590 8386
rect 5624 8352 5640 8386
rect 5489 8329 5640 8352
rect 5282 7654 5433 7677
rect 5282 7620 5298 7654
rect 5332 7620 5366 7654
rect 5400 7620 5433 7654
rect 5282 7597 5433 7620
rect 5489 7654 5640 7677
rect 5489 7620 5522 7654
rect 5556 7620 5590 7654
rect 5624 7620 5640 7654
rect 5489 7597 5640 7620
rect 5282 6922 5433 6945
rect 5282 6888 5298 6922
rect 5332 6888 5366 6922
rect 5400 6888 5433 6922
rect 5282 6865 5433 6888
rect 5489 6922 5640 6945
rect 5489 6888 5522 6922
rect 5556 6888 5590 6922
rect 5624 6888 5640 6922
rect 5489 6865 5640 6888
rect 5282 6190 5433 6213
rect 5282 6156 5298 6190
rect 5332 6156 5366 6190
rect 5400 6156 5433 6190
rect 5282 6133 5433 6156
rect 5489 6190 5640 6213
rect 5489 6156 5522 6190
rect 5556 6156 5590 6190
rect 5624 6156 5640 6190
rect 5489 6133 5640 6156
rect 5289 367 5545 383
rect 5289 333 5305 367
rect 5339 333 5400 367
rect 5434 333 5495 367
rect 5529 333 5545 367
rect 5289 317 5545 333
rect 5732 367 5988 383
rect 5732 333 5748 367
rect 5782 333 5843 367
rect 5877 333 5938 367
rect 5972 333 5988 367
rect 5732 317 5988 333
rect 5289 -432 5545 -409
rect 5289 -466 5305 -432
rect 5339 -466 5400 -432
rect 5434 -466 5495 -432
rect 5529 -466 5545 -432
rect 5289 -489 5545 -466
rect 5732 -432 5988 -409
rect 5732 -466 5748 -432
rect 5782 -466 5843 -432
rect 5877 -466 5938 -432
rect 5972 -466 5988 -432
rect 5732 -489 5988 -466
rect 5289 -1238 5545 -1215
rect 5289 -1272 5305 -1238
rect 5339 -1272 5400 -1238
rect 5434 -1272 5495 -1238
rect 5529 -1272 5545 -1238
rect 5289 -1295 5545 -1272
rect 5732 -1238 5988 -1215
rect 5732 -1272 5748 -1238
rect 5782 -1272 5843 -1238
rect 5877 -1272 5938 -1238
rect 5972 -1272 5988 -1238
rect 5732 -1295 5988 -1272
rect 5289 -2034 5545 -2011
rect 5289 -2068 5305 -2034
rect 5339 -2068 5400 -2034
rect 5434 -2068 5495 -2034
rect 5529 -2068 5545 -2034
rect 5289 -2091 5545 -2068
<< polycont >>
rect 5298 10548 5332 10582
rect 5366 10548 5400 10582
rect 5522 10548 5556 10582
rect 5590 10548 5624 10582
rect 5298 9816 5332 9850
rect 5366 9816 5400 9850
rect 5522 9816 5556 9850
rect 5590 9816 5624 9850
rect 5298 9084 5332 9118
rect 5366 9084 5400 9118
rect 5522 9084 5556 9118
rect 5590 9084 5624 9118
rect 5298 8352 5332 8386
rect 5366 8352 5400 8386
rect 5522 8352 5556 8386
rect 5590 8352 5624 8386
rect 5298 7620 5332 7654
rect 5366 7620 5400 7654
rect 5522 7620 5556 7654
rect 5590 7620 5624 7654
rect 5298 6888 5332 6922
rect 5366 6888 5400 6922
rect 5522 6888 5556 6922
rect 5590 6888 5624 6922
rect 5298 6156 5332 6190
rect 5366 6156 5400 6190
rect 5522 6156 5556 6190
rect 5590 6156 5624 6190
rect 5305 333 5339 367
rect 5400 333 5434 367
rect 5495 333 5529 367
rect 5748 333 5782 367
rect 5843 333 5877 367
rect 5938 333 5972 367
rect 5305 -466 5339 -432
rect 5400 -466 5434 -432
rect 5495 -466 5529 -432
rect 5748 -466 5782 -432
rect 5843 -466 5877 -432
rect 5938 -466 5972 -432
rect 5305 -1272 5339 -1238
rect 5400 -1272 5434 -1238
rect 5495 -1272 5529 -1238
rect 5748 -1272 5782 -1238
rect 5843 -1272 5877 -1238
rect 5938 -1272 5972 -1238
rect 5305 -2068 5339 -2034
rect 5400 -2068 5434 -2034
rect 5495 -2068 5529 -2034
<< locali >>
rect 4766 11169 6238 11175
rect 4766 11165 4845 11169
rect 4879 11165 4918 11169
rect 4952 11165 4991 11169
rect 5025 11165 5064 11169
rect 5098 11165 5137 11169
rect 5171 11165 5210 11169
rect 5244 11165 5284 11169
rect 5318 11165 5358 11169
rect 5392 11165 5432 11169
rect 5466 11165 5506 11169
rect 5540 11165 5580 11169
rect 5614 11165 5654 11169
rect 5688 11165 5728 11169
rect 5762 11165 5802 11169
rect 5836 11165 5876 11169
rect 5910 11165 5950 11169
rect 5984 11165 6024 11169
rect 6058 11165 6098 11169
rect 6132 11165 6172 11169
rect 4766 11097 4844 11165
rect 5318 11135 5321 11165
rect 5286 11131 5321 11135
rect 5355 11135 5358 11165
rect 5424 11135 5432 11165
rect 5493 11135 5506 11165
rect 5562 11135 5580 11165
rect 5631 11135 5654 11165
rect 5700 11135 5728 11165
rect 5769 11135 5802 11165
rect 5355 11131 5390 11135
rect 5424 11131 5459 11135
rect 5493 11131 5528 11135
rect 5562 11131 5597 11135
rect 5631 11131 5666 11135
rect 5700 11131 5735 11135
rect 5769 11131 5804 11135
rect 5838 11131 5873 11165
rect 5910 11135 5942 11165
rect 5984 11135 6011 11165
rect 6058 11135 6080 11165
rect 6132 11135 6149 11165
rect 6206 11135 6238 11169
rect 5907 11131 5942 11135
rect 5976 11131 6011 11135
rect 6045 11131 6080 11135
rect 6114 11131 6149 11135
rect 6183 11131 6238 11135
rect 5286 11097 6238 11131
rect 4766 11063 4772 11097
rect 4810 11063 4844 11097
rect 5318 11063 5321 11097
rect 5355 11063 5358 11097
rect 5424 11063 5432 11097
rect 5493 11063 5506 11097
rect 5562 11063 5580 11097
rect 5631 11063 5654 11097
rect 5700 11063 5728 11097
rect 5769 11063 5802 11097
rect 5838 11063 5873 11097
rect 5910 11063 5942 11097
rect 5984 11063 6011 11097
rect 6058 11063 6080 11097
rect 6132 11063 6149 11097
rect 6206 11063 6238 11097
rect 4766 11028 4912 11063
rect 4766 11024 4776 11028
rect 4766 10990 4772 11024
rect 4810 10994 4844 11028
rect 4878 10995 4912 11028
rect 5286 11029 6238 11063
rect 5286 11025 5321 11029
rect 5318 10995 5321 11025
rect 5355 11025 5390 11029
rect 5424 11025 5459 11029
rect 5493 11025 5528 11029
rect 5562 11025 5597 11029
rect 5631 11025 5666 11029
rect 5700 11025 5735 11029
rect 5769 11025 5804 11029
rect 5355 10995 5358 11025
rect 5424 10995 5432 11025
rect 5493 10995 5506 11025
rect 5562 10995 5580 11025
rect 5631 10995 5654 11025
rect 5700 10995 5728 11025
rect 5769 10995 5802 11025
rect 5838 10995 5873 11029
rect 5907 11025 5942 11029
rect 5976 11025 6011 11029
rect 6045 11025 6080 11029
rect 6114 11025 6149 11029
rect 6183 11025 6238 11029
rect 5910 10995 5942 11025
rect 5984 10995 6011 11025
rect 6058 10995 6080 11025
rect 6132 10995 6149 11025
rect 4806 10990 4844 10994
rect 4878 10991 4916 10995
rect 4950 10991 4989 10995
rect 5023 10991 5062 10995
rect 5096 10991 5136 10995
rect 5170 10991 5210 10995
rect 5244 10991 5284 10995
rect 5318 10991 5358 10995
rect 5392 10991 5432 10995
rect 5466 10991 5506 10995
rect 5540 10991 5580 10995
rect 5614 10991 5654 10995
rect 5688 10991 5728 10995
rect 5762 10991 5802 10995
rect 5836 10991 5876 10995
rect 5910 10991 5950 10995
rect 5984 10991 6024 10995
rect 6058 10991 6098 10995
rect 6132 10991 6172 10995
rect 6206 10991 6238 11025
rect 4878 10990 6238 10991
rect 4766 10985 6238 10990
rect 4766 10960 4956 10985
rect 4766 10959 4912 10960
rect 4766 10951 4776 10959
rect 4766 10917 4772 10951
rect 4810 10925 4844 10959
rect 4878 10926 4912 10959
rect 4946 10952 4956 10960
rect 4806 10917 4844 10925
rect 4878 10918 4916 10926
rect 4950 10918 4956 10952
rect 4878 10917 4956 10918
rect 4766 10891 4956 10917
rect 4766 10890 4912 10891
rect 4766 10878 4776 10890
rect 4766 10844 4772 10878
rect 4810 10856 4844 10890
rect 4878 10857 4912 10890
rect 4946 10879 4956 10891
rect 4806 10844 4844 10856
rect 4878 10845 4916 10857
rect 4950 10845 4956 10879
rect 4878 10844 4956 10845
rect 4766 10822 4956 10844
rect 4766 10821 4912 10822
rect 4766 10805 4776 10821
rect 4766 10771 4772 10805
rect 4810 10787 4844 10821
rect 4878 10788 4912 10821
rect 4946 10806 4956 10822
rect 4806 10771 4844 10787
rect 4878 10772 4916 10788
rect 4950 10772 4956 10806
rect 4878 10771 4956 10772
rect 4766 10753 4956 10771
rect 4766 10752 4912 10753
rect 4766 10732 4776 10752
rect 4766 10698 4772 10732
rect 4810 10718 4844 10752
rect 4878 10719 4912 10752
rect 4946 10733 4956 10753
rect 4806 10698 4844 10718
rect 4878 10699 4916 10719
rect 4950 10699 4956 10733
rect 4878 10698 4956 10699
rect 4766 10684 4956 10698
rect 4766 10683 4912 10684
rect 4766 10659 4776 10683
rect 4766 10625 4772 10659
rect 4810 10649 4844 10683
rect 4878 10650 4912 10683
rect 4946 10660 4956 10684
rect 4806 10625 4844 10649
rect 4878 10626 4916 10650
rect 4950 10626 4956 10660
rect 4878 10625 4956 10626
rect 4766 10615 4956 10625
rect 4766 10614 4912 10615
rect 4766 10586 4776 10614
rect 4766 10552 4772 10586
rect 4810 10580 4844 10614
rect 4878 10581 4912 10614
rect 4946 10587 4956 10615
rect 4806 10552 4844 10580
rect 4878 10553 4916 10581
rect 4950 10553 4956 10587
rect 4878 10552 4956 10553
rect 4766 10546 4956 10552
rect 4766 10545 4912 10546
rect 4766 10513 4776 10545
rect 4766 10479 4772 10513
rect 4810 10511 4844 10545
rect 4878 10512 4912 10545
rect 4946 10514 4956 10546
rect 4806 10479 4844 10511
rect 4878 10480 4916 10512
rect 4950 10480 4956 10514
rect 4878 10479 4956 10480
rect 4766 10477 4956 10479
rect 4766 10476 4912 10477
rect 4766 10442 4776 10476
rect 4810 10442 4844 10476
rect 4878 10443 4912 10476
rect 4946 10443 4956 10477
rect 4878 10442 4956 10443
rect 4766 10441 4956 10442
rect 4766 10440 4916 10441
rect 4766 10406 4772 10440
rect 4806 10407 4844 10440
rect 4878 10408 4916 10440
rect 4766 10373 4776 10406
rect 4810 10373 4844 10407
rect 4878 10374 4912 10408
rect 4950 10407 4956 10441
rect 4946 10374 4956 10407
rect 4878 10373 4956 10374
rect 4766 10368 4956 10373
rect 4766 10367 4916 10368
rect 4766 10333 4772 10367
rect 4806 10338 4844 10367
rect 4878 10339 4916 10367
rect 4766 10304 4776 10333
rect 4810 10304 4844 10338
rect 4878 10305 4912 10339
rect 4950 10334 4956 10368
rect 4946 10305 4956 10334
rect 4878 10304 4956 10305
rect 4766 10295 4956 10304
rect 4766 10294 4916 10295
rect 4766 10260 4772 10294
rect 4806 10269 4844 10294
rect 4878 10270 4916 10294
rect 4766 10235 4776 10260
rect 4810 10235 4844 10269
rect 4878 10236 4912 10270
rect 4950 10261 4956 10295
rect 4946 10236 4956 10261
rect 4878 10235 4956 10236
rect 4766 10222 4956 10235
rect 4766 10221 4916 10222
rect 4766 10187 4772 10221
rect 4806 10200 4844 10221
rect 4878 10201 4916 10221
rect 4766 10166 4776 10187
rect 4810 10166 4844 10200
rect 4878 10167 4912 10201
rect 4950 10188 4956 10222
rect 4946 10167 4956 10188
rect 4878 10166 4956 10167
rect 4766 10149 4956 10166
rect 4766 10148 4916 10149
rect 4766 10114 4772 10148
rect 4806 10131 4844 10148
rect 4878 10132 4916 10148
rect 4766 10097 4776 10114
rect 4810 10097 4844 10131
rect 4878 10098 4912 10132
rect 4950 10115 4956 10149
rect 4946 10098 4956 10115
rect 4878 10097 4956 10098
rect 4766 10076 4956 10097
rect 4766 10075 4916 10076
rect 4766 10041 4772 10075
rect 4806 10062 4844 10075
rect 4878 10063 4916 10075
rect 4766 10028 4776 10041
rect 4810 10028 4844 10062
rect 4878 10029 4912 10063
rect 4950 10042 4956 10076
rect 4946 10029 4956 10042
rect 4878 10028 4956 10029
rect 4766 10003 4956 10028
rect 4766 10002 4916 10003
rect 4766 9968 4772 10002
rect 4806 9993 4844 10002
rect 4878 9994 4916 10002
rect 4766 9959 4776 9968
rect 4810 9959 4844 9993
rect 4878 9960 4912 9994
rect 4950 9969 4956 10003
rect 4946 9960 4956 9969
rect 4878 9959 4956 9960
rect 4766 9930 4956 9959
rect 4766 9929 4916 9930
rect 4766 9895 4772 9929
rect 4806 9924 4844 9929
rect 4878 9925 4916 9929
rect 4766 9890 4776 9895
rect 4810 9890 4844 9924
rect 4878 9891 4912 9925
rect 4950 9896 4956 9930
rect 4946 9891 4956 9896
rect 4878 9890 4956 9891
rect 4766 9857 4956 9890
rect 4766 9856 4916 9857
rect 4766 9822 4772 9856
rect 4806 9855 4844 9856
rect 4766 9821 4776 9822
rect 4810 9821 4844 9855
rect 4878 9822 4912 9856
rect 4950 9823 4956 9857
rect 4946 9822 4956 9823
rect 4878 9821 4956 9822
rect 4766 9787 4956 9821
rect 4766 9786 4912 9787
rect 4766 9783 4776 9786
rect 4766 9749 4772 9783
rect 4810 9752 4844 9786
rect 4878 9753 4912 9786
rect 4946 9784 4956 9787
rect 4806 9749 4844 9752
rect 4878 9750 4916 9753
rect 4950 9750 4956 9784
rect 4878 9749 4956 9750
rect 4766 9718 4956 9749
rect 4766 9717 4912 9718
rect 4766 9710 4776 9717
rect 4766 9676 4772 9710
rect 4810 9683 4844 9717
rect 4878 9684 4912 9717
rect 4946 9711 4956 9718
rect 4806 9676 4844 9683
rect 4878 9677 4916 9684
rect 4950 9677 4956 9711
rect 4878 9676 4956 9677
rect 4766 9649 4956 9676
rect 4766 9648 4912 9649
rect 4766 9637 4776 9648
rect 4766 9603 4772 9637
rect 4810 9614 4844 9648
rect 4878 9615 4912 9648
rect 4946 9638 4956 9649
rect 4806 9603 4844 9614
rect 4878 9604 4916 9615
rect 4950 9604 4956 9638
rect 4878 9603 4956 9604
rect 4766 9580 4956 9603
rect 4766 9579 4912 9580
rect 4766 9564 4776 9579
rect 4766 9530 4772 9564
rect 4810 9545 4844 9579
rect 4878 9546 4912 9579
rect 4946 9565 4956 9580
rect 4806 9530 4844 9545
rect 4878 9531 4916 9546
rect 4950 9531 4956 9565
rect 4878 9530 4956 9531
rect 4766 9511 4956 9530
rect 4766 9510 4912 9511
rect 4766 9491 4776 9510
rect 4766 9457 4772 9491
rect 4810 9476 4844 9510
rect 4878 9477 4912 9510
rect 4946 9492 4956 9511
rect 4806 9457 4844 9476
rect 4878 9458 4916 9477
rect 4950 9458 4956 9492
rect 4878 9457 4956 9458
rect 4766 9442 4956 9457
rect 4766 9441 4912 9442
rect 4766 9418 4776 9441
rect 4766 9384 4772 9418
rect 4810 9407 4844 9441
rect 4878 9408 4912 9441
rect 4946 9419 4956 9442
rect 4806 9384 4844 9407
rect 4878 9385 4916 9408
rect 4950 9385 4956 9419
rect 4878 9384 4956 9385
rect 4766 9373 4956 9384
rect 4766 9372 4912 9373
rect 4766 9345 4776 9372
rect 4766 9311 4772 9345
rect 4810 9338 4844 9372
rect 4878 9339 4912 9372
rect 4946 9346 4956 9373
rect 4806 9311 4844 9338
rect 4878 9312 4916 9339
rect 4950 9312 4956 9346
rect 4878 9311 4956 9312
rect 4766 9304 4956 9311
rect 4766 9303 4912 9304
rect 4766 9272 4776 9303
rect 4766 9238 4772 9272
rect 4810 9269 4844 9303
rect 4878 9270 4912 9303
rect 4946 9273 4956 9304
rect 4806 9238 4844 9269
rect 4878 9239 4916 9270
rect 4950 9239 4956 9273
rect 4878 9238 4956 9239
rect 4766 9235 4956 9238
rect 4766 9234 4912 9235
rect 4766 9200 4776 9234
rect 4810 9200 4844 9234
rect 4878 9201 4912 9234
rect 4946 9201 4956 9235
rect 4878 9200 4956 9201
rect 4766 9199 4916 9200
rect 4766 9165 4772 9199
rect 4806 9165 4844 9199
rect 4878 9166 4916 9199
rect 4950 9166 4956 9200
rect 4766 9131 4776 9165
rect 4810 9131 4844 9165
rect 4878 9132 4912 9166
rect 4946 9132 4956 9166
rect 4878 9131 4956 9132
rect 4766 9127 4956 9131
rect 4766 9126 4916 9127
rect 4766 9092 4772 9126
rect 4806 9096 4844 9126
rect 4878 9097 4916 9126
rect 4766 9062 4776 9092
rect 4810 9062 4844 9096
rect 4878 9063 4912 9097
rect 4950 9093 4956 9127
rect 4946 9063 4956 9093
rect 4878 9062 4956 9063
rect 4766 9054 4956 9062
rect 4766 9053 4916 9054
rect 4766 9019 4772 9053
rect 4806 9027 4844 9053
rect 4878 9028 4916 9053
rect 4766 8993 4776 9019
rect 4810 8993 4844 9027
rect 4878 8994 4912 9028
rect 4950 9020 4956 9054
rect 4946 8994 4956 9020
rect 4878 8993 4956 8994
rect 4766 8981 4956 8993
rect 4766 8980 4916 8981
rect 4766 8946 4772 8980
rect 4806 8958 4844 8980
rect 4878 8959 4916 8980
rect 4766 8924 4776 8946
rect 4810 8924 4844 8958
rect 4878 8925 4912 8959
rect 4950 8947 4956 8981
rect 4946 8925 4956 8947
rect 4878 8924 4956 8925
rect 4766 8908 4956 8924
rect 4766 8907 4916 8908
rect 4766 8873 4772 8907
rect 4806 8889 4844 8907
rect 4878 8890 4916 8907
rect 4766 8855 4776 8873
rect 4810 8855 4844 8889
rect 4878 8856 4912 8890
rect 4950 8874 4956 8908
rect 4946 8856 4956 8874
rect 4878 8855 4956 8856
rect 4766 8835 4956 8855
rect 4766 8834 4916 8835
rect 4766 4264 4772 8834
rect 4878 8821 4916 8834
rect 4878 8787 4912 8821
rect 4950 8801 4956 8835
rect 4946 8787 4956 8801
rect 4878 8762 4956 8787
rect 4950 4376 4956 8762
rect 5090 10845 5832 10851
rect 5090 10809 5174 10845
rect 5208 10811 5252 10845
rect 5286 10843 5330 10845
rect 5364 10843 5408 10845
rect 5442 10843 5486 10845
rect 5520 10843 5564 10845
rect 5598 10843 5642 10845
rect 5676 10843 5720 10845
rect 5754 10843 5832 10845
rect 5286 10811 5314 10843
rect 5208 10809 5314 10811
rect 5090 10775 5314 10809
rect 5090 10773 5098 10775
rect 5200 10773 5314 10775
rect 5756 10773 5832 10843
rect 5090 10739 5096 10773
rect 5202 10739 5252 10773
rect 5286 10741 5314 10773
rect 5286 10739 5330 10741
rect 5364 10739 5408 10741
rect 5442 10739 5486 10741
rect 5520 10739 5564 10741
rect 5598 10739 5642 10741
rect 5676 10739 5720 10741
rect 5090 10700 5098 10739
rect 5200 10733 5720 10739
rect 5200 10700 5208 10733
rect 5090 10666 5096 10700
rect 5202 10666 5208 10700
rect 5090 10627 5098 10666
rect 5200 10627 5208 10666
rect 5090 10593 5096 10627
rect 5202 10593 5208 10627
rect 5090 10554 5098 10593
rect 5200 10554 5208 10593
rect 5714 10667 5720 10733
rect 5826 10667 5832 10773
rect 5714 10628 5722 10667
rect 5824 10628 5832 10667
rect 5714 10594 5720 10628
rect 5826 10594 5832 10628
rect 5090 10520 5096 10554
rect 5202 10520 5208 10554
rect 5282 10582 5416 10589
rect 5282 10548 5298 10582
rect 5332 10548 5366 10582
rect 5282 10541 5366 10548
rect 5090 10481 5098 10520
rect 5200 10481 5208 10520
rect 5090 10447 5096 10481
rect 5202 10447 5208 10481
rect 5400 10541 5416 10582
rect 5506 10582 5640 10589
rect 5506 10541 5522 10582
rect 5556 10548 5590 10582
rect 5624 10548 5640 10582
rect 5366 10499 5400 10537
rect 5556 10541 5640 10548
rect 5714 10555 5722 10594
rect 5824 10555 5832 10594
rect 5522 10499 5556 10537
rect 5714 10521 5720 10555
rect 5826 10521 5832 10555
rect 5714 10482 5722 10521
rect 5824 10482 5832 10521
rect 5090 10408 5098 10447
rect 5200 10408 5208 10447
rect 5090 10374 5096 10408
rect 5202 10374 5208 10408
rect 5090 10335 5098 10374
rect 5200 10335 5208 10374
rect 5090 10301 5096 10335
rect 5202 10301 5208 10335
rect 5090 10262 5098 10301
rect 5200 10262 5208 10301
rect 5090 10228 5096 10262
rect 5202 10228 5208 10262
rect 5090 10189 5098 10228
rect 5200 10189 5208 10228
rect 5090 10155 5096 10189
rect 5202 10155 5208 10189
rect 5090 10116 5098 10155
rect 5200 10116 5208 10155
rect 5090 4610 5096 10116
rect 5202 4650 5208 10116
rect 5714 10448 5720 10482
rect 5826 10448 5832 10482
rect 5714 10409 5722 10448
rect 5824 10409 5832 10448
rect 5714 10375 5720 10409
rect 5826 10375 5832 10409
rect 5714 10336 5722 10375
rect 5824 10336 5832 10375
rect 5714 10302 5720 10336
rect 5826 10302 5832 10336
rect 5714 10263 5722 10302
rect 5824 10263 5832 10302
rect 5714 10229 5720 10263
rect 5826 10229 5832 10263
rect 5714 10190 5722 10229
rect 5824 10190 5832 10229
rect 5714 10156 5720 10190
rect 5826 10156 5832 10190
rect 5714 10117 5722 10156
rect 5824 10117 5832 10156
rect 5714 10083 5720 10117
rect 5826 10083 5832 10117
rect 5714 10044 5722 10083
rect 5824 10044 5832 10083
rect 5714 10010 5720 10044
rect 5826 10010 5832 10044
rect 5714 9971 5722 10010
rect 5824 9971 5832 10010
rect 5714 9937 5720 9971
rect 5826 9937 5832 9971
rect 5714 9898 5722 9937
rect 5824 9898 5832 9937
rect 5282 9852 5366 9857
rect 5400 9852 5416 9857
rect 5282 9850 5416 9852
rect 5282 9816 5298 9850
rect 5332 9816 5366 9850
rect 5400 9816 5416 9850
rect 5282 9814 5416 9816
rect 5282 9809 5366 9814
rect 5400 9809 5416 9814
rect 5506 9852 5522 9857
rect 5714 9864 5720 9898
rect 5826 9864 5832 9898
rect 5556 9852 5640 9857
rect 5506 9850 5640 9852
rect 5506 9816 5522 9850
rect 5556 9816 5590 9850
rect 5624 9816 5640 9850
rect 5506 9814 5640 9816
rect 5506 9809 5522 9814
rect 5556 9809 5640 9814
rect 5714 9825 5722 9864
rect 5824 9825 5832 9864
rect 5714 9791 5720 9825
rect 5826 9791 5832 9825
rect 5714 9752 5722 9791
rect 5824 9752 5832 9791
rect 5714 9718 5720 9752
rect 5826 9718 5832 9752
rect 5714 9679 5722 9718
rect 5824 9679 5832 9718
rect 5714 9645 5720 9679
rect 5826 9645 5832 9679
rect 5714 9606 5722 9645
rect 5824 9606 5832 9645
rect 5714 9572 5720 9606
rect 5826 9572 5832 9606
rect 5714 9533 5722 9572
rect 5824 9533 5832 9572
rect 5714 9499 5720 9533
rect 5826 9499 5832 9533
rect 5714 9460 5722 9499
rect 5824 9460 5832 9499
rect 5714 9426 5720 9460
rect 5826 9426 5832 9460
rect 5714 9387 5722 9426
rect 5824 9387 5832 9426
rect 5714 9353 5720 9387
rect 5826 9353 5832 9387
rect 5714 9314 5722 9353
rect 5824 9314 5832 9353
rect 5714 9280 5720 9314
rect 5826 9280 5832 9314
rect 5714 9216 5722 9280
rect 5824 9216 5832 9280
rect 5714 9182 5720 9216
rect 5826 9182 5832 9216
rect 5282 9120 5366 9125
rect 5400 9120 5416 9125
rect 5282 9118 5416 9120
rect 5282 9084 5298 9118
rect 5332 9084 5366 9118
rect 5400 9084 5416 9118
rect 5282 9082 5416 9084
rect 5282 9077 5366 9082
rect 5400 9077 5416 9082
rect 5506 9120 5522 9125
rect 5714 9143 5722 9182
rect 5824 9143 5832 9182
rect 5556 9120 5640 9125
rect 5506 9118 5640 9120
rect 5506 9084 5522 9118
rect 5556 9084 5590 9118
rect 5624 9084 5640 9118
rect 5506 9082 5640 9084
rect 5506 9077 5522 9082
rect 5556 9077 5640 9082
rect 5714 9109 5720 9143
rect 5826 9109 5832 9143
rect 5714 9070 5722 9109
rect 5824 9070 5832 9109
rect 5714 9036 5720 9070
rect 5826 9036 5832 9070
rect 5714 8997 5722 9036
rect 5824 8997 5832 9036
rect 5714 8963 5720 8997
rect 5826 8963 5832 8997
rect 5714 8924 5722 8963
rect 5824 8924 5832 8963
rect 5714 8890 5720 8924
rect 5826 8890 5832 8924
rect 5714 8851 5722 8890
rect 5824 8851 5832 8890
rect 5714 8817 5720 8851
rect 5826 8817 5832 8851
rect 5714 8778 5722 8817
rect 5824 8778 5832 8817
rect 5714 8744 5720 8778
rect 5826 8744 5832 8778
rect 5714 8705 5722 8744
rect 5824 8705 5832 8744
rect 5714 8671 5720 8705
rect 5826 8671 5832 8705
rect 5714 8632 5722 8671
rect 5824 8632 5832 8671
rect 5714 8598 5720 8632
rect 5826 8598 5832 8632
rect 5714 8559 5722 8598
rect 5824 8559 5832 8598
rect 5714 8525 5720 8559
rect 5826 8525 5832 8559
rect 5714 8486 5722 8525
rect 5824 8486 5832 8525
rect 5714 8452 5720 8486
rect 5826 8452 5832 8486
rect 5282 8388 5366 8393
rect 5400 8388 5416 8393
rect 5282 8386 5416 8388
rect 5282 8352 5298 8386
rect 5332 8352 5366 8386
rect 5400 8352 5416 8386
rect 5282 8350 5416 8352
rect 5282 8345 5366 8350
rect 5400 8345 5416 8350
rect 5506 8388 5522 8393
rect 5714 8413 5722 8452
rect 5824 8413 5832 8452
rect 5556 8388 5640 8393
rect 5506 8386 5640 8388
rect 5506 8352 5522 8386
rect 5556 8352 5590 8386
rect 5624 8352 5640 8386
rect 5506 8350 5640 8352
rect 5506 8345 5522 8350
rect 5556 8345 5640 8350
rect 5714 8379 5720 8413
rect 5826 8379 5832 8413
rect 5714 8340 5722 8379
rect 5824 8340 5832 8379
rect 5714 8306 5720 8340
rect 5826 8306 5832 8340
rect 5714 8267 5722 8306
rect 5824 8267 5832 8306
rect 5714 8233 5720 8267
rect 5826 8233 5832 8267
rect 5714 8194 5722 8233
rect 5824 8194 5832 8233
rect 5714 8160 5720 8194
rect 5826 8160 5832 8194
rect 5714 8121 5722 8160
rect 5824 8121 5832 8160
rect 5714 8087 5720 8121
rect 5826 8087 5832 8121
rect 5714 8048 5722 8087
rect 5824 8048 5832 8087
rect 5714 8014 5720 8048
rect 5826 8014 5832 8048
rect 5714 7975 5722 8014
rect 5824 7975 5832 8014
rect 5714 7941 5720 7975
rect 5826 7941 5832 7975
rect 5714 7902 5722 7941
rect 5824 7902 5832 7941
rect 5714 7868 5720 7902
rect 5826 7868 5832 7902
rect 5714 7829 5722 7868
rect 5824 7829 5832 7868
rect 5714 7795 5720 7829
rect 5826 7795 5832 7829
rect 5714 7756 5722 7795
rect 5824 7756 5832 7795
rect 5714 7722 5720 7756
rect 5826 7722 5832 7756
rect 5282 7656 5366 7661
rect 5400 7656 5416 7661
rect 5282 7654 5416 7656
rect 5282 7620 5298 7654
rect 5332 7620 5366 7654
rect 5400 7620 5416 7654
rect 5282 7618 5416 7620
rect 5282 7613 5366 7618
rect 5400 7613 5416 7618
rect 5506 7656 5522 7661
rect 5714 7683 5722 7722
rect 5824 7683 5832 7722
rect 5556 7656 5640 7661
rect 5506 7654 5640 7656
rect 5506 7620 5522 7654
rect 5556 7620 5590 7654
rect 5624 7620 5640 7654
rect 5506 7618 5640 7620
rect 5506 7613 5522 7618
rect 5556 7613 5640 7618
rect 5714 7649 5720 7683
rect 5826 7649 5832 7683
rect 5714 7610 5722 7649
rect 5824 7610 5832 7649
rect 5714 7576 5720 7610
rect 5826 7576 5832 7610
rect 5714 7537 5722 7576
rect 5824 7537 5832 7576
rect 5714 7503 5720 7537
rect 5826 7503 5832 7537
rect 5714 7464 5722 7503
rect 5824 7464 5832 7503
rect 5714 7430 5720 7464
rect 5826 7430 5832 7464
rect 5714 7391 5722 7430
rect 5824 7391 5832 7430
rect 5714 7357 5720 7391
rect 5826 7357 5832 7391
rect 5714 7318 5722 7357
rect 5824 7318 5832 7357
rect 5714 7284 5720 7318
rect 5826 7284 5832 7318
rect 5714 7245 5722 7284
rect 5824 7245 5832 7284
rect 5714 7211 5720 7245
rect 5826 7211 5832 7245
rect 5714 7172 5722 7211
rect 5824 7172 5832 7211
rect 5714 7138 5720 7172
rect 5826 7138 5832 7172
rect 5714 7099 5722 7138
rect 5824 7099 5832 7138
rect 5714 7065 5720 7099
rect 5826 7065 5832 7099
rect 5714 7026 5722 7065
rect 5824 7026 5832 7065
rect 5714 6992 5720 7026
rect 5826 6992 5832 7026
rect 5282 6924 5366 6929
rect 5400 6924 5416 6929
rect 5282 6922 5416 6924
rect 5282 6888 5298 6922
rect 5332 6888 5366 6922
rect 5400 6888 5416 6922
rect 5282 6886 5416 6888
rect 5282 6881 5366 6886
rect 5400 6881 5416 6886
rect 5506 6924 5522 6929
rect 5714 6953 5722 6992
rect 5824 6953 5832 6992
rect 5556 6924 5640 6929
rect 5506 6922 5640 6924
rect 5506 6888 5522 6922
rect 5556 6888 5590 6922
rect 5624 6888 5640 6922
rect 5506 6886 5640 6888
rect 5506 6881 5522 6886
rect 5556 6881 5640 6886
rect 5714 6919 5720 6953
rect 5826 6919 5832 6953
rect 5714 6880 5722 6919
rect 5824 6880 5832 6919
rect 5714 6846 5720 6880
rect 5826 6846 5832 6880
rect 5714 6807 5722 6846
rect 5824 6807 5832 6846
rect 5714 6773 5720 6807
rect 5826 6773 5832 6807
rect 5714 6734 5722 6773
rect 5824 6734 5832 6773
rect 5714 6700 5720 6734
rect 5826 6700 5832 6734
rect 5714 6661 5722 6700
rect 5824 6661 5832 6700
rect 5282 6192 5366 6197
rect 5400 6192 5416 6197
rect 5282 6190 5416 6192
rect 5282 6156 5298 6190
rect 5332 6156 5366 6190
rect 5400 6156 5416 6190
rect 5282 6154 5416 6156
rect 5282 6149 5366 6154
rect 5400 6149 5416 6154
rect 5506 6192 5522 6197
rect 5556 6192 5640 6197
rect 5506 6190 5640 6192
rect 5506 6156 5522 6190
rect 5556 6156 5590 6190
rect 5624 6156 5640 6190
rect 5506 6154 5640 6156
rect 5506 6149 5522 6154
rect 5556 6149 5640 6154
rect 5714 4683 5720 6661
rect 5826 4683 5832 6661
rect 5714 4650 5722 4683
rect 5202 4644 5722 4650
rect 5202 4642 5244 4644
rect 5278 4642 5320 4644
rect 5354 4642 5395 4644
rect 5429 4642 5470 4644
rect 5504 4642 5545 4644
rect 5579 4642 5620 4644
rect 5654 4642 5695 4644
rect 5676 4610 5695 4642
rect 5090 4540 5166 4610
rect 5676 4608 5722 4610
rect 5824 4608 5832 4683
rect 5676 4595 5832 4608
rect 5676 4574 5792 4595
rect 5676 4540 5710 4574
rect 5744 4572 5792 4574
rect 5748 4561 5792 4572
rect 5826 4561 5832 4595
rect 5090 4538 5168 4540
rect 5202 4538 5246 4540
rect 5280 4538 5324 4540
rect 5358 4538 5402 4540
rect 5436 4538 5480 4540
rect 5514 4538 5558 4540
rect 5592 4538 5636 4540
rect 5670 4538 5714 4540
rect 5748 4538 5832 4561
rect 5090 4532 5832 4538
rect 4950 4370 6238 4376
rect 4950 4367 4990 4370
rect 5024 4367 5064 4370
rect 5098 4367 5138 4370
rect 5172 4367 5212 4370
rect 5246 4367 5286 4370
rect 5320 4367 5360 4370
rect 4950 4336 4981 4367
rect 5024 4336 5050 4367
rect 5098 4336 5119 4367
rect 5172 4336 5188 4367
rect 5246 4336 5257 4367
rect 5320 4336 5326 4367
rect 4946 4333 4981 4336
rect 5015 4333 5050 4336
rect 5084 4333 5119 4336
rect 5153 4333 5188 4336
rect 5222 4333 5257 4336
rect 5291 4333 5326 4336
rect 5394 4367 5434 4370
rect 5468 4367 5508 4370
rect 5542 4367 5582 4370
rect 5616 4367 5656 4370
rect 5690 4367 5730 4370
rect 5764 4367 5804 4370
rect 5838 4367 5878 4370
rect 5912 4367 5952 4370
rect 5986 4367 6026 4370
rect 6060 4367 6099 4370
rect 6133 4367 6172 4370
rect 5394 4336 5395 4367
rect 5360 4333 5395 4336
rect 5429 4336 5434 4367
rect 5498 4336 5508 4367
rect 5567 4336 5582 4367
rect 5636 4336 5656 4367
rect 5705 4336 5730 4367
rect 5774 4336 5804 4367
rect 6206 4336 6238 4370
rect 5429 4333 5464 4336
rect 5498 4333 5533 4336
rect 5567 4333 5602 4336
rect 5636 4333 5671 4336
rect 5705 4333 5740 4336
rect 5774 4333 5809 4336
rect 4878 4299 5809 4333
rect 4878 4265 4913 4299
rect 4947 4298 4982 4299
rect 5016 4298 5051 4299
rect 5085 4298 5120 4299
rect 5154 4298 5189 4299
rect 5223 4298 5258 4299
rect 5292 4298 5327 4299
rect 4952 4265 4982 4298
rect 5026 4265 5051 4298
rect 5100 4265 5120 4298
rect 5174 4265 5189 4298
rect 5248 4265 5258 4298
rect 5322 4265 5327 4298
rect 5361 4298 5396 4299
rect 5361 4265 5362 4298
rect 4878 4264 4918 4265
rect 4952 4264 4992 4265
rect 5026 4264 5066 4265
rect 5100 4264 5140 4265
rect 5174 4264 5214 4265
rect 5248 4264 5288 4265
rect 5322 4264 5362 4265
rect 5430 4298 5465 4299
rect 5499 4298 5534 4299
rect 5568 4298 5603 4299
rect 5637 4298 5672 4299
rect 5706 4298 5741 4299
rect 6183 4298 6238 4336
rect 5430 4265 5436 4298
rect 5499 4265 5510 4298
rect 5568 4265 5584 4298
rect 5637 4265 5658 4298
rect 5706 4265 5732 4298
rect 5396 4264 5436 4265
rect 5470 4264 5510 4265
rect 5544 4264 5584 4265
rect 5618 4264 5658 4265
rect 5692 4264 5732 4265
rect 6206 4264 6238 4298
rect 4766 4231 5741 4264
rect 4766 4192 4844 4231
rect 4878 4197 4913 4231
rect 4947 4226 4982 4231
rect 5016 4226 5051 4231
rect 5085 4226 5120 4231
rect 5154 4226 5189 4231
rect 5223 4226 5258 4231
rect 5292 4226 5327 4231
rect 4952 4197 4982 4226
rect 5026 4197 5051 4226
rect 5100 4197 5120 4226
rect 5174 4197 5189 4226
rect 5248 4197 5258 4226
rect 5322 4197 5327 4226
rect 5361 4226 5396 4231
rect 5361 4197 5362 4226
rect 4878 4192 4918 4197
rect 4952 4192 4992 4197
rect 5026 4192 5066 4197
rect 5100 4192 5140 4197
rect 5174 4192 5214 4197
rect 5248 4192 5288 4197
rect 5322 4192 5362 4197
rect 5430 4226 5465 4231
rect 5499 4226 5534 4231
rect 5568 4226 5603 4231
rect 5637 4226 5672 4231
rect 5706 4226 5741 4231
rect 6183 4226 6238 4264
rect 5430 4197 5436 4226
rect 5499 4197 5510 4226
rect 5568 4197 5584 4226
rect 5637 4197 5658 4226
rect 5706 4197 5732 4226
rect 5396 4192 5436 4197
rect 5470 4192 5510 4197
rect 5544 4192 5584 4197
rect 5618 4192 5658 4197
rect 5692 4192 5732 4197
rect 5766 4192 5806 4197
rect 5840 4192 5880 4197
rect 5914 4192 5953 4197
rect 5987 4192 6026 4197
rect 6060 4192 6099 4197
rect 6133 4192 6172 4197
rect 6206 4192 6238 4226
rect 4766 4186 6238 4192
rect 5289 333 5301 367
rect 5339 333 5382 367
rect 5434 333 5462 367
rect 5529 333 5542 367
rect 5576 333 5622 367
rect 5656 333 5702 367
rect 5736 333 5748 367
rect 5816 333 5843 367
rect 5896 333 5938 367
rect 5976 333 5988 367
rect 5244 159 5278 198
rect 5244 85 5278 125
rect 5535 159 5569 198
rect 5535 85 5569 125
rect 5687 18 5721 93
rect 5999 18 6033 93
rect 5400 -81 5434 -43
rect 5843 -242 5877 -204
rect 5289 -432 5545 -425
rect 5732 -432 5988 -425
rect 5289 -466 5301 -432
rect 5339 -466 5382 -432
rect 5434 -466 5462 -432
rect 5529 -466 5542 -432
rect 5576 -466 5622 -432
rect 5656 -466 5702 -432
rect 5736 -466 5748 -432
rect 5816 -466 5843 -432
rect 5896 -466 5938 -432
rect 5976 -466 5988 -432
rect 5289 -473 5545 -466
rect 5732 -473 5988 -466
rect 5244 -602 5278 -563
rect 5244 -676 5278 -636
rect 5556 -602 5590 -563
rect 5556 -676 5590 -636
rect 5687 -602 5721 -563
rect 5687 -676 5721 -636
rect 5999 -602 6033 -563
rect 5999 -676 6033 -636
rect 5400 -863 5434 -825
rect 5843 -949 5877 -911
rect 5289 -1238 5545 -1231
rect 5732 -1238 5988 -1231
rect 5289 -1272 5301 -1238
rect 5339 -1272 5382 -1238
rect 5434 -1272 5462 -1238
rect 5529 -1272 5542 -1238
rect 5576 -1272 5622 -1238
rect 5656 -1272 5702 -1238
rect 5736 -1272 5748 -1238
rect 5816 -1272 5843 -1238
rect 5896 -1272 5938 -1238
rect 5976 -1272 5988 -1238
rect 5289 -1279 5545 -1272
rect 5732 -1279 5988 -1272
rect 5244 -1396 5278 -1357
rect 5244 -1470 5278 -1430
rect 5556 -1396 5590 -1357
rect 5556 -1470 5590 -1430
rect 5687 -1396 5721 -1357
rect 5687 -1470 5721 -1430
rect 5999 -1396 6033 -1357
rect 5999 -1470 6033 -1430
rect 5400 -1659 5434 -1621
rect 5843 -1745 5877 -1707
rect 5289 -2034 5545 -2027
rect 5289 -2068 5301 -2034
rect 5339 -2068 5400 -2034
rect 5434 -2068 5495 -2034
rect 5533 -2068 5545 -2034
rect 5289 -2075 5545 -2068
rect 5244 -2204 5278 -2165
rect 5244 -2278 5278 -2238
rect 5556 -2204 5590 -2165
rect 5556 -2278 5590 -2238
rect 5400 -2440 5434 -2402
<< viali >>
rect 4845 11165 4879 11169
rect 4918 11165 4952 11169
rect 4991 11165 5025 11169
rect 5064 11165 5098 11169
rect 5137 11165 5171 11169
rect 5210 11165 5244 11169
rect 5284 11165 5318 11169
rect 5358 11165 5392 11169
rect 5432 11165 5466 11169
rect 5506 11165 5540 11169
rect 5580 11165 5614 11169
rect 5654 11165 5688 11169
rect 5728 11165 5762 11169
rect 5802 11165 5836 11169
rect 5876 11165 5910 11169
rect 5950 11165 5984 11169
rect 6024 11165 6058 11169
rect 6098 11165 6132 11169
rect 6172 11165 6206 11169
rect 4845 11135 4879 11165
rect 4918 11135 4952 11165
rect 4991 11135 5025 11165
rect 5064 11135 5098 11165
rect 5137 11135 5171 11165
rect 5210 11135 5244 11165
rect 5284 11135 5286 11165
rect 5286 11135 5318 11165
rect 5358 11135 5390 11165
rect 5390 11135 5392 11165
rect 5432 11135 5459 11165
rect 5459 11135 5466 11165
rect 5506 11135 5528 11165
rect 5528 11135 5540 11165
rect 5580 11135 5597 11165
rect 5597 11135 5614 11165
rect 5654 11135 5666 11165
rect 5666 11135 5688 11165
rect 5728 11135 5735 11165
rect 5735 11135 5762 11165
rect 5802 11135 5804 11165
rect 5804 11135 5836 11165
rect 5876 11135 5907 11165
rect 5907 11135 5910 11165
rect 5950 11135 5976 11165
rect 5976 11135 5984 11165
rect 6024 11135 6045 11165
rect 6045 11135 6058 11165
rect 6098 11135 6114 11165
rect 6114 11135 6132 11165
rect 6172 11135 6183 11165
rect 6183 11135 6206 11165
rect 4772 11063 4776 11097
rect 4776 11063 4806 11097
rect 4844 11063 4878 11097
rect 4918 11063 4952 11097
rect 4991 11063 5025 11097
rect 5064 11063 5098 11097
rect 5137 11063 5171 11097
rect 5210 11063 5244 11097
rect 5284 11063 5286 11097
rect 5286 11063 5318 11097
rect 5358 11063 5390 11097
rect 5390 11063 5392 11097
rect 5432 11063 5459 11097
rect 5459 11063 5466 11097
rect 5506 11063 5528 11097
rect 5528 11063 5540 11097
rect 5580 11063 5597 11097
rect 5597 11063 5614 11097
rect 5654 11063 5666 11097
rect 5666 11063 5688 11097
rect 5728 11063 5735 11097
rect 5735 11063 5762 11097
rect 5802 11063 5804 11097
rect 5804 11063 5836 11097
rect 5876 11063 5907 11097
rect 5907 11063 5910 11097
rect 5950 11063 5976 11097
rect 5976 11063 5984 11097
rect 6024 11063 6045 11097
rect 6045 11063 6058 11097
rect 6098 11063 6114 11097
rect 6114 11063 6132 11097
rect 6172 11063 6183 11097
rect 6183 11063 6206 11097
rect 4772 10994 4776 11024
rect 4776 10994 4806 11024
rect 4844 10994 4878 11024
rect 4916 10995 4950 11025
rect 4989 10995 5023 11025
rect 5062 10995 5096 11025
rect 5136 10995 5170 11025
rect 5210 10995 5244 11025
rect 5284 10995 5286 11025
rect 5286 10995 5318 11025
rect 5358 10995 5390 11025
rect 5390 10995 5392 11025
rect 5432 10995 5459 11025
rect 5459 10995 5466 11025
rect 5506 10995 5528 11025
rect 5528 10995 5540 11025
rect 5580 10995 5597 11025
rect 5597 10995 5614 11025
rect 5654 10995 5666 11025
rect 5666 10995 5688 11025
rect 5728 10995 5735 11025
rect 5735 10995 5762 11025
rect 5802 10995 5804 11025
rect 5804 10995 5836 11025
rect 5876 10995 5907 11025
rect 5907 10995 5910 11025
rect 5950 10995 5976 11025
rect 5976 10995 5984 11025
rect 6024 10995 6045 11025
rect 6045 10995 6058 11025
rect 6098 10995 6114 11025
rect 6114 10995 6132 11025
rect 6172 10995 6183 11025
rect 6183 10995 6206 11025
rect 4772 10990 4806 10994
rect 4844 10990 4878 10994
rect 4916 10991 4950 10995
rect 4989 10991 5023 10995
rect 5062 10991 5096 10995
rect 5136 10991 5170 10995
rect 5210 10991 5244 10995
rect 5284 10991 5318 10995
rect 5358 10991 5392 10995
rect 5432 10991 5466 10995
rect 5506 10991 5540 10995
rect 5580 10991 5614 10995
rect 5654 10991 5688 10995
rect 5728 10991 5762 10995
rect 5802 10991 5836 10995
rect 5876 10991 5910 10995
rect 5950 10991 5984 10995
rect 6024 10991 6058 10995
rect 6098 10991 6132 10995
rect 6172 10991 6206 10995
rect 4772 10925 4776 10951
rect 4776 10925 4806 10951
rect 4844 10925 4878 10951
rect 4916 10926 4946 10952
rect 4946 10926 4950 10952
rect 4772 10917 4806 10925
rect 4844 10917 4878 10925
rect 4916 10918 4950 10926
rect 4772 10856 4776 10878
rect 4776 10856 4806 10878
rect 4844 10856 4878 10878
rect 4916 10857 4946 10879
rect 4946 10857 4950 10879
rect 4772 10844 4806 10856
rect 4844 10844 4878 10856
rect 4916 10845 4950 10857
rect 4772 10787 4776 10805
rect 4776 10787 4806 10805
rect 4844 10787 4878 10805
rect 4916 10788 4946 10806
rect 4946 10788 4950 10806
rect 4772 10771 4806 10787
rect 4844 10771 4878 10787
rect 4916 10772 4950 10788
rect 4772 10718 4776 10732
rect 4776 10718 4806 10732
rect 4844 10718 4878 10732
rect 4916 10719 4946 10733
rect 4946 10719 4950 10733
rect 4772 10698 4806 10718
rect 4844 10698 4878 10718
rect 4916 10699 4950 10719
rect 4772 10649 4776 10659
rect 4776 10649 4806 10659
rect 4844 10649 4878 10659
rect 4916 10650 4946 10660
rect 4946 10650 4950 10660
rect 4772 10625 4806 10649
rect 4844 10625 4878 10649
rect 4916 10626 4950 10650
rect 4772 10580 4776 10586
rect 4776 10580 4806 10586
rect 4844 10580 4878 10586
rect 4916 10581 4946 10587
rect 4946 10581 4950 10587
rect 4772 10552 4806 10580
rect 4844 10552 4878 10580
rect 4916 10553 4950 10581
rect 4772 10511 4776 10513
rect 4776 10511 4806 10513
rect 4844 10511 4878 10513
rect 4916 10512 4946 10514
rect 4946 10512 4950 10514
rect 4772 10479 4806 10511
rect 4844 10479 4878 10511
rect 4916 10480 4950 10512
rect 4772 10407 4806 10440
rect 4844 10407 4878 10440
rect 4916 10408 4950 10441
rect 4772 10406 4776 10407
rect 4776 10406 4806 10407
rect 4844 10406 4878 10407
rect 4916 10407 4946 10408
rect 4946 10407 4950 10408
rect 4772 10338 4806 10367
rect 4844 10338 4878 10367
rect 4916 10339 4950 10368
rect 4772 10333 4776 10338
rect 4776 10333 4806 10338
rect 4844 10333 4878 10338
rect 4916 10334 4946 10339
rect 4946 10334 4950 10339
rect 4772 10269 4806 10294
rect 4844 10269 4878 10294
rect 4916 10270 4950 10295
rect 4772 10260 4776 10269
rect 4776 10260 4806 10269
rect 4844 10260 4878 10269
rect 4916 10261 4946 10270
rect 4946 10261 4950 10270
rect 4772 10200 4806 10221
rect 4844 10200 4878 10221
rect 4916 10201 4950 10222
rect 4772 10187 4776 10200
rect 4776 10187 4806 10200
rect 4844 10187 4878 10200
rect 4916 10188 4946 10201
rect 4946 10188 4950 10201
rect 4772 10131 4806 10148
rect 4844 10131 4878 10148
rect 4916 10132 4950 10149
rect 4772 10114 4776 10131
rect 4776 10114 4806 10131
rect 4844 10114 4878 10131
rect 4916 10115 4946 10132
rect 4946 10115 4950 10132
rect 4772 10062 4806 10075
rect 4844 10062 4878 10075
rect 4916 10063 4950 10076
rect 4772 10041 4776 10062
rect 4776 10041 4806 10062
rect 4844 10041 4878 10062
rect 4916 10042 4946 10063
rect 4946 10042 4950 10063
rect 4772 9993 4806 10002
rect 4844 9993 4878 10002
rect 4916 9994 4950 10003
rect 4772 9968 4776 9993
rect 4776 9968 4806 9993
rect 4844 9968 4878 9993
rect 4916 9969 4946 9994
rect 4946 9969 4950 9994
rect 4772 9924 4806 9929
rect 4844 9924 4878 9929
rect 4916 9925 4950 9930
rect 4772 9895 4776 9924
rect 4776 9895 4806 9924
rect 4844 9895 4878 9924
rect 4916 9896 4946 9925
rect 4946 9896 4950 9925
rect 4916 9856 4950 9857
rect 4772 9855 4806 9856
rect 4844 9855 4878 9856
rect 4772 9822 4776 9855
rect 4776 9822 4806 9855
rect 4844 9822 4878 9855
rect 4916 9823 4946 9856
rect 4946 9823 4950 9856
rect 4772 9752 4776 9783
rect 4776 9752 4806 9783
rect 4844 9752 4878 9783
rect 4916 9753 4946 9784
rect 4946 9753 4950 9784
rect 4772 9749 4806 9752
rect 4844 9749 4878 9752
rect 4916 9750 4950 9753
rect 4772 9683 4776 9710
rect 4776 9683 4806 9710
rect 4844 9683 4878 9710
rect 4916 9684 4946 9711
rect 4946 9684 4950 9711
rect 4772 9676 4806 9683
rect 4844 9676 4878 9683
rect 4916 9677 4950 9684
rect 4772 9614 4776 9637
rect 4776 9614 4806 9637
rect 4844 9614 4878 9637
rect 4916 9615 4946 9638
rect 4946 9615 4950 9638
rect 4772 9603 4806 9614
rect 4844 9603 4878 9614
rect 4916 9604 4950 9615
rect 4772 9545 4776 9564
rect 4776 9545 4806 9564
rect 4844 9545 4878 9564
rect 4916 9546 4946 9565
rect 4946 9546 4950 9565
rect 4772 9530 4806 9545
rect 4844 9530 4878 9545
rect 4916 9531 4950 9546
rect 4772 9476 4776 9491
rect 4776 9476 4806 9491
rect 4844 9476 4878 9491
rect 4916 9477 4946 9492
rect 4946 9477 4950 9492
rect 4772 9457 4806 9476
rect 4844 9457 4878 9476
rect 4916 9458 4950 9477
rect 4772 9407 4776 9418
rect 4776 9407 4806 9418
rect 4844 9407 4878 9418
rect 4916 9408 4946 9419
rect 4946 9408 4950 9419
rect 4772 9384 4806 9407
rect 4844 9384 4878 9407
rect 4916 9385 4950 9408
rect 4772 9338 4776 9345
rect 4776 9338 4806 9345
rect 4844 9338 4878 9345
rect 4916 9339 4946 9346
rect 4946 9339 4950 9346
rect 4772 9311 4806 9338
rect 4844 9311 4878 9338
rect 4916 9312 4950 9339
rect 4772 9269 4776 9272
rect 4776 9269 4806 9272
rect 4844 9269 4878 9272
rect 4916 9270 4946 9273
rect 4946 9270 4950 9273
rect 4772 9238 4806 9269
rect 4844 9238 4878 9269
rect 4916 9239 4950 9270
rect 4772 9165 4806 9199
rect 4844 9165 4878 9199
rect 4916 9166 4950 9200
rect 4772 9096 4806 9126
rect 4844 9096 4878 9126
rect 4916 9097 4950 9127
rect 4772 9092 4776 9096
rect 4776 9092 4806 9096
rect 4844 9092 4878 9096
rect 4916 9093 4946 9097
rect 4946 9093 4950 9097
rect 4772 9027 4806 9053
rect 4844 9027 4878 9053
rect 4916 9028 4950 9054
rect 4772 9019 4776 9027
rect 4776 9019 4806 9027
rect 4844 9019 4878 9027
rect 4916 9020 4946 9028
rect 4946 9020 4950 9028
rect 4772 8958 4806 8980
rect 4844 8958 4878 8980
rect 4916 8959 4950 8981
rect 4772 8946 4776 8958
rect 4776 8946 4806 8958
rect 4844 8946 4878 8958
rect 4916 8947 4946 8959
rect 4946 8947 4950 8959
rect 4772 8889 4806 8907
rect 4844 8889 4878 8907
rect 4916 8890 4950 8908
rect 4772 8873 4776 8889
rect 4776 8873 4806 8889
rect 4844 8873 4878 8889
rect 4916 8874 4946 8890
rect 4946 8874 4950 8890
rect 4772 8820 4878 8834
rect 4916 8821 4950 8835
rect 4772 8786 4776 8820
rect 4776 8786 4810 8820
rect 4810 8786 4844 8820
rect 4844 8786 4878 8820
rect 4916 8801 4946 8821
rect 4946 8801 4950 8821
rect 4772 8762 4878 8786
rect 4772 8752 4950 8762
rect 4772 8751 4912 8752
rect 4772 8717 4776 8751
rect 4776 8717 4810 8751
rect 4810 8717 4844 8751
rect 4844 8717 4878 8751
rect 4878 8718 4912 8751
rect 4912 8718 4946 8752
rect 4946 8718 4950 8752
rect 4878 8717 4950 8718
rect 4772 8683 4950 8717
rect 4772 8682 4912 8683
rect 4772 8648 4776 8682
rect 4776 8648 4810 8682
rect 4810 8648 4844 8682
rect 4844 8648 4878 8682
rect 4878 8649 4912 8682
rect 4912 8649 4946 8683
rect 4946 8649 4950 8683
rect 4878 8648 4950 8649
rect 4772 8614 4950 8648
rect 4772 8613 4912 8614
rect 4772 8579 4776 8613
rect 4776 8579 4810 8613
rect 4810 8579 4844 8613
rect 4844 8579 4878 8613
rect 4878 8580 4912 8613
rect 4912 8580 4946 8614
rect 4946 8580 4950 8614
rect 4878 8579 4950 8580
rect 4772 8545 4950 8579
rect 4772 8544 4912 8545
rect 4772 8510 4776 8544
rect 4776 8510 4810 8544
rect 4810 8510 4844 8544
rect 4844 8510 4878 8544
rect 4878 8511 4912 8544
rect 4912 8511 4946 8545
rect 4946 8511 4950 8545
rect 4878 8510 4950 8511
rect 4772 8476 4950 8510
rect 4772 8475 4912 8476
rect 4772 8441 4776 8475
rect 4776 8441 4810 8475
rect 4810 8441 4844 8475
rect 4844 8441 4878 8475
rect 4878 8442 4912 8475
rect 4912 8442 4946 8476
rect 4946 8442 4950 8476
rect 4878 8441 4950 8442
rect 4772 8407 4950 8441
rect 4772 8406 4912 8407
rect 4772 8372 4776 8406
rect 4776 8372 4810 8406
rect 4810 8372 4844 8406
rect 4844 8372 4878 8406
rect 4878 8373 4912 8406
rect 4912 8373 4946 8407
rect 4946 8373 4950 8407
rect 4878 8372 4950 8373
rect 4772 8338 4950 8372
rect 4772 8337 4912 8338
rect 4772 8303 4776 8337
rect 4776 8303 4810 8337
rect 4810 8303 4844 8337
rect 4844 8303 4878 8337
rect 4878 8304 4912 8337
rect 4912 8304 4946 8338
rect 4946 8304 4950 8338
rect 4878 8303 4950 8304
rect 4772 8269 4950 8303
rect 4772 8268 4912 8269
rect 4772 8234 4776 8268
rect 4776 8234 4810 8268
rect 4810 8234 4844 8268
rect 4844 8234 4878 8268
rect 4878 8235 4912 8268
rect 4912 8235 4946 8269
rect 4946 8235 4950 8269
rect 4878 8234 4950 8235
rect 4772 8200 4950 8234
rect 4772 8199 4912 8200
rect 4772 8165 4776 8199
rect 4776 8165 4810 8199
rect 4810 8165 4844 8199
rect 4844 8165 4878 8199
rect 4878 8166 4912 8199
rect 4912 8166 4946 8200
rect 4946 8166 4950 8200
rect 4878 8165 4950 8166
rect 4772 8131 4950 8165
rect 4772 8130 4912 8131
rect 4772 8096 4776 8130
rect 4776 8096 4810 8130
rect 4810 8096 4844 8130
rect 4844 8096 4878 8130
rect 4878 8097 4912 8130
rect 4912 8097 4946 8131
rect 4946 8097 4950 8131
rect 4878 8096 4950 8097
rect 4772 8062 4950 8096
rect 4772 8061 4912 8062
rect 4772 8027 4776 8061
rect 4776 8027 4810 8061
rect 4810 8027 4844 8061
rect 4844 8027 4878 8061
rect 4878 8028 4912 8061
rect 4912 8028 4946 8062
rect 4946 8028 4950 8062
rect 4878 8027 4950 8028
rect 4772 7993 4950 8027
rect 4772 7992 4912 7993
rect 4772 7958 4776 7992
rect 4776 7958 4810 7992
rect 4810 7958 4844 7992
rect 4844 7958 4878 7992
rect 4878 7959 4912 7992
rect 4912 7959 4946 7993
rect 4946 7959 4950 7993
rect 4878 7958 4950 7959
rect 4772 7924 4950 7958
rect 4772 7923 4912 7924
rect 4772 7889 4776 7923
rect 4776 7889 4810 7923
rect 4810 7889 4844 7923
rect 4844 7889 4878 7923
rect 4878 7890 4912 7923
rect 4912 7890 4946 7924
rect 4946 7890 4950 7924
rect 4878 7889 4950 7890
rect 4772 7855 4950 7889
rect 4772 7854 4912 7855
rect 4772 7820 4776 7854
rect 4776 7820 4810 7854
rect 4810 7820 4844 7854
rect 4844 7820 4878 7854
rect 4878 7821 4912 7854
rect 4912 7821 4946 7855
rect 4946 7821 4950 7855
rect 4878 7820 4950 7821
rect 4772 7786 4950 7820
rect 4772 7785 4912 7786
rect 4772 7751 4776 7785
rect 4776 7751 4810 7785
rect 4810 7751 4844 7785
rect 4844 7751 4878 7785
rect 4878 7752 4912 7785
rect 4912 7752 4946 7786
rect 4946 7752 4950 7786
rect 4878 7751 4950 7752
rect 4772 7717 4950 7751
rect 4772 7716 4912 7717
rect 4772 7682 4776 7716
rect 4776 7682 4810 7716
rect 4810 7682 4844 7716
rect 4844 7682 4878 7716
rect 4878 7683 4912 7716
rect 4912 7683 4946 7717
rect 4946 7683 4950 7717
rect 4878 7682 4950 7683
rect 4772 7648 4950 7682
rect 4772 7647 4912 7648
rect 4772 7613 4776 7647
rect 4776 7613 4810 7647
rect 4810 7613 4844 7647
rect 4844 7613 4878 7647
rect 4878 7614 4912 7647
rect 4912 7614 4946 7648
rect 4946 7614 4950 7648
rect 4878 7613 4950 7614
rect 4772 7579 4950 7613
rect 4772 7578 4912 7579
rect 4772 7544 4776 7578
rect 4776 7544 4810 7578
rect 4810 7544 4844 7578
rect 4844 7544 4878 7578
rect 4878 7545 4912 7578
rect 4912 7545 4946 7579
rect 4946 7545 4950 7579
rect 4878 7544 4950 7545
rect 4772 7510 4950 7544
rect 4772 7509 4912 7510
rect 4772 7475 4776 7509
rect 4776 7475 4810 7509
rect 4810 7475 4844 7509
rect 4844 7475 4878 7509
rect 4878 7476 4912 7509
rect 4912 7476 4946 7510
rect 4946 7476 4950 7510
rect 4878 7475 4950 7476
rect 4772 7441 4950 7475
rect 4772 7440 4912 7441
rect 4772 7406 4776 7440
rect 4776 7406 4810 7440
rect 4810 7406 4844 7440
rect 4844 7406 4878 7440
rect 4878 7407 4912 7440
rect 4912 7407 4946 7441
rect 4946 7407 4950 7441
rect 4878 7406 4950 7407
rect 4772 7372 4950 7406
rect 4772 7371 4912 7372
rect 4772 7337 4776 7371
rect 4776 7337 4810 7371
rect 4810 7337 4844 7371
rect 4844 7337 4878 7371
rect 4878 7338 4912 7371
rect 4912 7338 4946 7372
rect 4946 7338 4950 7372
rect 4878 7337 4950 7338
rect 4772 7303 4950 7337
rect 4772 7302 4912 7303
rect 4772 7268 4776 7302
rect 4776 7268 4810 7302
rect 4810 7268 4844 7302
rect 4844 7268 4878 7302
rect 4878 7269 4912 7302
rect 4912 7269 4946 7303
rect 4946 7269 4950 7303
rect 4878 7268 4950 7269
rect 4772 7234 4950 7268
rect 4772 7233 4912 7234
rect 4772 7199 4776 7233
rect 4776 7199 4810 7233
rect 4810 7199 4844 7233
rect 4844 7199 4878 7233
rect 4878 7200 4912 7233
rect 4912 7200 4946 7234
rect 4946 7200 4950 7234
rect 4878 7199 4950 7200
rect 4772 7165 4950 7199
rect 4772 7164 4912 7165
rect 4772 7130 4776 7164
rect 4776 7130 4810 7164
rect 4810 7130 4844 7164
rect 4844 7130 4878 7164
rect 4878 7131 4912 7164
rect 4912 7131 4946 7165
rect 4946 7131 4950 7165
rect 4878 7130 4950 7131
rect 4772 7096 4950 7130
rect 4772 7095 4912 7096
rect 4772 7061 4776 7095
rect 4776 7061 4810 7095
rect 4810 7061 4844 7095
rect 4844 7061 4878 7095
rect 4878 7062 4912 7095
rect 4912 7062 4946 7096
rect 4946 7062 4950 7096
rect 4878 7061 4950 7062
rect 4772 7027 4950 7061
rect 4772 7026 4912 7027
rect 4772 6992 4776 7026
rect 4776 6992 4810 7026
rect 4810 6992 4844 7026
rect 4844 6992 4878 7026
rect 4878 6993 4912 7026
rect 4912 6993 4946 7027
rect 4946 6993 4950 7027
rect 4878 6992 4950 6993
rect 4772 6958 4950 6992
rect 4772 6957 4912 6958
rect 4772 6923 4776 6957
rect 4776 6923 4810 6957
rect 4810 6923 4844 6957
rect 4844 6923 4878 6957
rect 4878 6924 4912 6957
rect 4912 6924 4946 6958
rect 4946 6924 4950 6958
rect 4878 6923 4950 6924
rect 4772 6889 4950 6923
rect 4772 6888 4912 6889
rect 4772 6854 4776 6888
rect 4776 6854 4810 6888
rect 4810 6854 4844 6888
rect 4844 6854 4878 6888
rect 4878 6855 4912 6888
rect 4912 6855 4946 6889
rect 4946 6855 4950 6889
rect 4878 6854 4950 6855
rect 4772 6820 4950 6854
rect 4772 6819 4912 6820
rect 4772 6785 4776 6819
rect 4776 6785 4810 6819
rect 4810 6785 4844 6819
rect 4844 6785 4878 6819
rect 4878 6786 4912 6819
rect 4912 6786 4946 6820
rect 4946 6786 4950 6820
rect 4878 6785 4950 6786
rect 4772 6751 4950 6785
rect 4772 6750 4912 6751
rect 4772 6716 4776 6750
rect 4776 6716 4810 6750
rect 4810 6716 4844 6750
rect 4844 6716 4878 6750
rect 4878 6717 4912 6750
rect 4912 6717 4946 6751
rect 4946 6717 4950 6751
rect 4878 6716 4950 6717
rect 4772 6682 4950 6716
rect 4772 6681 4912 6682
rect 4772 6647 4776 6681
rect 4776 6647 4810 6681
rect 4810 6647 4844 6681
rect 4844 6647 4878 6681
rect 4878 6648 4912 6681
rect 4912 6648 4946 6682
rect 4946 6648 4950 6682
rect 4878 6647 4950 6648
rect 4772 6613 4950 6647
rect 4772 6612 4912 6613
rect 4772 6578 4776 6612
rect 4776 6578 4810 6612
rect 4810 6578 4844 6612
rect 4844 6578 4878 6612
rect 4878 6579 4912 6612
rect 4912 6579 4946 6613
rect 4946 6579 4950 6613
rect 4878 6578 4950 6579
rect 4772 6544 4950 6578
rect 4772 6543 4912 6544
rect 4772 4265 4776 6543
rect 4776 6475 4878 6543
rect 4878 6510 4912 6543
rect 4912 6510 4946 6544
rect 4946 6510 4950 6544
rect 4878 6475 4950 6510
rect 4776 4336 4946 6475
rect 4946 4336 4950 6475
rect 5174 10843 5208 10845
rect 5174 10811 5208 10843
rect 5252 10811 5286 10845
rect 5330 10843 5364 10845
rect 5408 10843 5442 10845
rect 5486 10843 5520 10845
rect 5564 10843 5598 10845
rect 5642 10843 5676 10845
rect 5720 10843 5754 10845
rect 5330 10811 5364 10843
rect 5408 10811 5442 10843
rect 5486 10811 5520 10843
rect 5564 10811 5598 10843
rect 5642 10811 5676 10843
rect 5720 10811 5754 10843
rect 5096 10739 5098 10773
rect 5098 10739 5130 10773
rect 5168 10739 5200 10773
rect 5200 10739 5202 10773
rect 5252 10739 5286 10773
rect 5330 10741 5364 10773
rect 5408 10741 5442 10773
rect 5486 10741 5520 10773
rect 5564 10741 5598 10773
rect 5642 10741 5676 10773
rect 5720 10741 5756 10773
rect 5756 10762 5826 10773
rect 5756 10741 5790 10762
rect 5330 10739 5364 10741
rect 5408 10739 5442 10741
rect 5486 10739 5520 10741
rect 5564 10739 5598 10741
rect 5642 10739 5676 10741
rect 5096 10666 5098 10700
rect 5098 10666 5130 10700
rect 5168 10666 5200 10700
rect 5200 10666 5202 10700
rect 5096 10593 5098 10627
rect 5098 10593 5130 10627
rect 5168 10593 5200 10627
rect 5200 10593 5202 10627
rect 5720 10728 5790 10741
rect 5790 10728 5824 10762
rect 5824 10728 5826 10762
rect 5720 10694 5826 10728
rect 5720 10667 5722 10694
rect 5722 10667 5824 10694
rect 5824 10667 5826 10694
rect 5720 10594 5722 10628
rect 5722 10594 5754 10628
rect 5792 10594 5824 10628
rect 5824 10594 5826 10628
rect 5096 10520 5098 10554
rect 5098 10520 5130 10554
rect 5168 10520 5200 10554
rect 5200 10520 5202 10554
rect 5366 10548 5400 10571
rect 5096 10447 5098 10481
rect 5098 10447 5130 10481
rect 5168 10447 5200 10481
rect 5200 10447 5202 10481
rect 5366 10537 5400 10548
rect 5522 10548 5556 10571
rect 5366 10465 5400 10499
rect 5522 10537 5556 10548
rect 5522 10465 5556 10499
rect 5720 10521 5722 10555
rect 5722 10521 5754 10555
rect 5792 10521 5824 10555
rect 5824 10521 5826 10555
rect 5096 10374 5098 10408
rect 5098 10374 5130 10408
rect 5168 10374 5200 10408
rect 5200 10374 5202 10408
rect 5096 10301 5098 10335
rect 5098 10301 5130 10335
rect 5168 10301 5200 10335
rect 5200 10301 5202 10335
rect 5096 10228 5098 10262
rect 5098 10228 5130 10262
rect 5168 10228 5200 10262
rect 5200 10228 5202 10262
rect 5096 10155 5098 10189
rect 5098 10155 5130 10189
rect 5168 10155 5200 10189
rect 5200 10155 5202 10189
rect 5096 4961 5098 10116
rect 5098 4961 5200 10116
rect 5200 4961 5202 10116
rect 5096 4927 5202 4961
rect 5096 4689 5098 4927
rect 5098 4689 5200 4927
rect 5200 4689 5202 4927
rect 5096 4655 5202 4689
rect 5096 4621 5098 4655
rect 5098 4621 5132 4655
rect 5132 4642 5202 4655
rect 5720 10448 5722 10482
rect 5722 10448 5754 10482
rect 5792 10448 5824 10482
rect 5824 10448 5826 10482
rect 5720 10375 5722 10409
rect 5722 10375 5754 10409
rect 5792 10375 5824 10409
rect 5824 10375 5826 10409
rect 5720 10302 5722 10336
rect 5722 10302 5754 10336
rect 5792 10302 5824 10336
rect 5824 10302 5826 10336
rect 5720 10229 5722 10263
rect 5722 10229 5754 10263
rect 5792 10229 5824 10263
rect 5824 10229 5826 10263
rect 5720 10156 5722 10190
rect 5722 10156 5754 10190
rect 5792 10156 5824 10190
rect 5824 10156 5826 10190
rect 5720 10083 5722 10117
rect 5722 10083 5754 10117
rect 5792 10083 5824 10117
rect 5824 10083 5826 10117
rect 5720 10010 5722 10044
rect 5722 10010 5754 10044
rect 5792 10010 5824 10044
rect 5824 10010 5826 10044
rect 5720 9937 5722 9971
rect 5722 9937 5754 9971
rect 5792 9937 5824 9971
rect 5824 9937 5826 9971
rect 5366 9852 5400 9886
rect 5366 9780 5400 9814
rect 5522 9852 5556 9886
rect 5720 9864 5722 9898
rect 5722 9864 5754 9898
rect 5792 9864 5824 9898
rect 5824 9864 5826 9898
rect 5522 9780 5556 9814
rect 5720 9791 5722 9825
rect 5722 9791 5754 9825
rect 5792 9791 5824 9825
rect 5824 9791 5826 9825
rect 5720 9718 5722 9752
rect 5722 9718 5754 9752
rect 5792 9718 5824 9752
rect 5824 9718 5826 9752
rect 5720 9645 5722 9679
rect 5722 9645 5754 9679
rect 5792 9645 5824 9679
rect 5824 9645 5826 9679
rect 5720 9572 5722 9606
rect 5722 9572 5754 9606
rect 5792 9572 5824 9606
rect 5824 9572 5826 9606
rect 5720 9499 5722 9533
rect 5722 9499 5754 9533
rect 5792 9499 5824 9533
rect 5824 9499 5826 9533
rect 5720 9426 5722 9460
rect 5722 9426 5754 9460
rect 5792 9426 5824 9460
rect 5824 9426 5826 9460
rect 5720 9353 5722 9387
rect 5722 9353 5754 9387
rect 5792 9353 5824 9387
rect 5824 9353 5826 9387
rect 5720 9280 5722 9314
rect 5722 9280 5754 9314
rect 5792 9280 5824 9314
rect 5824 9280 5826 9314
rect 5720 9182 5722 9216
rect 5722 9182 5754 9216
rect 5792 9182 5824 9216
rect 5824 9182 5826 9216
rect 5366 9120 5400 9154
rect 5366 9048 5400 9082
rect 5522 9120 5556 9154
rect 5522 9048 5556 9082
rect 5720 9109 5722 9143
rect 5722 9109 5754 9143
rect 5792 9109 5824 9143
rect 5824 9109 5826 9143
rect 5720 9036 5722 9070
rect 5722 9036 5754 9070
rect 5792 9036 5824 9070
rect 5824 9036 5826 9070
rect 5720 8963 5722 8997
rect 5722 8963 5754 8997
rect 5792 8963 5824 8997
rect 5824 8963 5826 8997
rect 5720 8890 5722 8924
rect 5722 8890 5754 8924
rect 5792 8890 5824 8924
rect 5824 8890 5826 8924
rect 5720 8817 5722 8851
rect 5722 8817 5754 8851
rect 5792 8817 5824 8851
rect 5824 8817 5826 8851
rect 5720 8744 5722 8778
rect 5722 8744 5754 8778
rect 5792 8744 5824 8778
rect 5824 8744 5826 8778
rect 5720 8671 5722 8705
rect 5722 8671 5754 8705
rect 5792 8671 5824 8705
rect 5824 8671 5826 8705
rect 5720 8598 5722 8632
rect 5722 8598 5754 8632
rect 5792 8598 5824 8632
rect 5824 8598 5826 8632
rect 5720 8525 5722 8559
rect 5722 8525 5754 8559
rect 5792 8525 5824 8559
rect 5824 8525 5826 8559
rect 5720 8452 5722 8486
rect 5722 8452 5754 8486
rect 5792 8452 5824 8486
rect 5824 8452 5826 8486
rect 5366 8388 5400 8422
rect 5366 8316 5400 8350
rect 5522 8388 5556 8422
rect 5522 8316 5556 8350
rect 5720 8379 5722 8413
rect 5722 8379 5754 8413
rect 5792 8379 5824 8413
rect 5824 8379 5826 8413
rect 5720 8306 5722 8340
rect 5722 8306 5754 8340
rect 5792 8306 5824 8340
rect 5824 8306 5826 8340
rect 5720 8233 5722 8267
rect 5722 8233 5754 8267
rect 5792 8233 5824 8267
rect 5824 8233 5826 8267
rect 5720 8160 5722 8194
rect 5722 8160 5754 8194
rect 5792 8160 5824 8194
rect 5824 8160 5826 8194
rect 5720 8087 5722 8121
rect 5722 8087 5754 8121
rect 5792 8087 5824 8121
rect 5824 8087 5826 8121
rect 5720 8014 5722 8048
rect 5722 8014 5754 8048
rect 5792 8014 5824 8048
rect 5824 8014 5826 8048
rect 5720 7941 5722 7975
rect 5722 7941 5754 7975
rect 5792 7941 5824 7975
rect 5824 7941 5826 7975
rect 5720 7868 5722 7902
rect 5722 7868 5754 7902
rect 5792 7868 5824 7902
rect 5824 7868 5826 7902
rect 5720 7795 5722 7829
rect 5722 7795 5754 7829
rect 5792 7795 5824 7829
rect 5824 7795 5826 7829
rect 5720 7722 5722 7756
rect 5722 7722 5754 7756
rect 5792 7722 5824 7756
rect 5824 7722 5826 7756
rect 5366 7656 5400 7690
rect 5366 7584 5400 7618
rect 5522 7656 5556 7690
rect 5522 7584 5556 7618
rect 5720 7649 5722 7683
rect 5722 7649 5754 7683
rect 5792 7649 5824 7683
rect 5824 7649 5826 7683
rect 5720 7576 5722 7610
rect 5722 7576 5754 7610
rect 5792 7576 5824 7610
rect 5824 7576 5826 7610
rect 5720 7503 5722 7537
rect 5722 7503 5754 7537
rect 5792 7503 5824 7537
rect 5824 7503 5826 7537
rect 5720 7430 5722 7464
rect 5722 7430 5754 7464
rect 5792 7430 5824 7464
rect 5824 7430 5826 7464
rect 5720 7357 5722 7391
rect 5722 7357 5754 7391
rect 5792 7357 5824 7391
rect 5824 7357 5826 7391
rect 5720 7284 5722 7318
rect 5722 7284 5754 7318
rect 5792 7284 5824 7318
rect 5824 7284 5826 7318
rect 5720 7211 5722 7245
rect 5722 7211 5754 7245
rect 5792 7211 5824 7245
rect 5824 7211 5826 7245
rect 5720 7138 5722 7172
rect 5722 7138 5754 7172
rect 5792 7138 5824 7172
rect 5824 7138 5826 7172
rect 5720 7065 5722 7099
rect 5722 7065 5754 7099
rect 5792 7065 5824 7099
rect 5824 7065 5826 7099
rect 5720 6992 5722 7026
rect 5722 6992 5754 7026
rect 5792 6992 5824 7026
rect 5824 6992 5826 7026
rect 5366 6924 5400 6958
rect 5366 6852 5400 6886
rect 5522 6924 5556 6958
rect 5522 6852 5556 6886
rect 5720 6919 5722 6953
rect 5722 6919 5754 6953
rect 5792 6919 5824 6953
rect 5824 6919 5826 6953
rect 5720 6846 5722 6880
rect 5722 6846 5754 6880
rect 5792 6846 5824 6880
rect 5824 6846 5826 6880
rect 5720 6773 5722 6807
rect 5722 6773 5754 6807
rect 5792 6773 5824 6807
rect 5824 6773 5826 6807
rect 5720 6700 5722 6734
rect 5722 6700 5754 6734
rect 5792 6700 5824 6734
rect 5824 6700 5826 6734
rect 5366 6192 5400 6226
rect 5366 6120 5400 6154
rect 5522 6192 5556 6226
rect 5522 6120 5556 6154
rect 5720 4683 5722 6661
rect 5722 4956 5824 6661
rect 5722 4683 5824 4956
rect 5824 4683 5826 6661
rect 5244 4642 5278 4644
rect 5320 4642 5354 4644
rect 5395 4642 5429 4644
rect 5470 4642 5504 4644
rect 5545 4642 5579 4644
rect 5620 4642 5654 4644
rect 5132 4621 5166 4642
rect 5096 4610 5166 4621
rect 5166 4610 5202 4642
rect 5244 4610 5278 4642
rect 5320 4610 5354 4642
rect 5395 4610 5429 4642
rect 5470 4610 5504 4642
rect 5545 4610 5579 4642
rect 5620 4610 5654 4642
rect 5695 4610 5722 4644
rect 5722 4610 5729 4644
rect 5168 4540 5202 4572
rect 5246 4540 5280 4572
rect 5324 4540 5358 4572
rect 5402 4540 5436 4572
rect 5480 4540 5514 4572
rect 5558 4540 5592 4572
rect 5636 4540 5670 4572
rect 5714 4540 5744 4572
rect 5744 4540 5748 4572
rect 5792 4561 5826 4595
rect 5168 4538 5202 4540
rect 5246 4538 5280 4540
rect 5324 4538 5358 4540
rect 5402 4538 5436 4540
rect 5480 4538 5514 4540
rect 5558 4538 5592 4540
rect 5636 4538 5670 4540
rect 5714 4538 5748 4540
rect 4990 4367 5024 4370
rect 5064 4367 5098 4370
rect 5138 4367 5172 4370
rect 5212 4367 5246 4370
rect 5286 4367 5320 4370
rect 4990 4336 5015 4367
rect 5015 4336 5024 4367
rect 5064 4336 5084 4367
rect 5084 4336 5098 4367
rect 5138 4336 5153 4367
rect 5153 4336 5172 4367
rect 5212 4336 5222 4367
rect 5222 4336 5246 4367
rect 5286 4336 5291 4367
rect 5291 4336 5320 4367
rect 4776 4265 4878 4336
rect 5360 4336 5394 4370
rect 5434 4367 5468 4370
rect 5508 4367 5542 4370
rect 5582 4367 5616 4370
rect 5656 4367 5690 4370
rect 5730 4367 5764 4370
rect 5804 4367 5838 4370
rect 5878 4367 5912 4370
rect 5952 4367 5986 4370
rect 6026 4367 6060 4370
rect 6099 4367 6133 4370
rect 6172 4367 6206 4370
rect 5434 4336 5464 4367
rect 5464 4336 5468 4367
rect 5508 4336 5533 4367
rect 5533 4336 5542 4367
rect 5582 4336 5602 4367
rect 5602 4336 5616 4367
rect 5656 4336 5671 4367
rect 5671 4336 5690 4367
rect 5730 4336 5740 4367
rect 5740 4336 5764 4367
rect 5804 4336 5809 4367
rect 5809 4336 5838 4367
rect 5878 4336 5912 4367
rect 5952 4336 5986 4367
rect 6026 4336 6060 4367
rect 6099 4336 6133 4367
rect 6172 4336 6183 4367
rect 6183 4336 6206 4367
rect 4918 4265 4947 4298
rect 4947 4265 4952 4298
rect 4992 4265 5016 4298
rect 5016 4265 5026 4298
rect 5066 4265 5085 4298
rect 5085 4265 5100 4298
rect 5140 4265 5154 4298
rect 5154 4265 5174 4298
rect 5214 4265 5223 4298
rect 5223 4265 5248 4298
rect 5288 4265 5292 4298
rect 5292 4265 5322 4298
rect 4772 4264 4878 4265
rect 4918 4264 4952 4265
rect 4992 4264 5026 4265
rect 5066 4264 5100 4265
rect 5140 4264 5174 4265
rect 5214 4264 5248 4265
rect 5288 4264 5322 4265
rect 5362 4264 5396 4298
rect 5436 4265 5465 4298
rect 5465 4265 5470 4298
rect 5510 4265 5534 4298
rect 5534 4265 5544 4298
rect 5584 4265 5603 4298
rect 5603 4265 5618 4298
rect 5658 4265 5672 4298
rect 5672 4265 5692 4298
rect 5436 4264 5470 4265
rect 5510 4264 5544 4265
rect 5584 4264 5618 4265
rect 5658 4264 5692 4265
rect 5732 4264 5741 4298
rect 5741 4264 5766 4298
rect 5806 4264 5840 4298
rect 5880 4264 5914 4298
rect 5953 4264 5987 4298
rect 6026 4264 6060 4298
rect 6099 4264 6133 4298
rect 6172 4264 6183 4298
rect 6183 4264 6206 4298
rect 4844 4197 4878 4226
rect 4918 4197 4947 4226
rect 4947 4197 4952 4226
rect 4992 4197 5016 4226
rect 5016 4197 5026 4226
rect 5066 4197 5085 4226
rect 5085 4197 5100 4226
rect 5140 4197 5154 4226
rect 5154 4197 5174 4226
rect 5214 4197 5223 4226
rect 5223 4197 5248 4226
rect 5288 4197 5292 4226
rect 5292 4197 5322 4226
rect 4844 4192 4878 4197
rect 4918 4192 4952 4197
rect 4992 4192 5026 4197
rect 5066 4192 5100 4197
rect 5140 4192 5174 4197
rect 5214 4192 5248 4197
rect 5288 4192 5322 4197
rect 5362 4192 5396 4226
rect 5436 4197 5465 4226
rect 5465 4197 5470 4226
rect 5510 4197 5534 4226
rect 5534 4197 5544 4226
rect 5584 4197 5603 4226
rect 5603 4197 5618 4226
rect 5658 4197 5672 4226
rect 5672 4197 5692 4226
rect 5732 4197 5741 4226
rect 5741 4197 5766 4226
rect 5806 4197 5840 4226
rect 5880 4197 5914 4226
rect 5953 4197 5987 4226
rect 6026 4197 6060 4226
rect 6099 4197 6133 4226
rect 6172 4197 6183 4226
rect 6183 4197 6206 4226
rect 5436 4192 5470 4197
rect 5510 4192 5544 4197
rect 5584 4192 5618 4197
rect 5658 4192 5692 4197
rect 5732 4192 5766 4197
rect 5806 4192 5840 4197
rect 5880 4192 5914 4197
rect 5953 4192 5987 4197
rect 6026 4192 6060 4197
rect 6099 4192 6133 4197
rect 6172 4192 6206 4197
rect 5301 333 5305 367
rect 5305 333 5335 367
rect 5382 333 5400 367
rect 5400 333 5416 367
rect 5462 333 5495 367
rect 5495 333 5496 367
rect 5542 333 5576 367
rect 5622 333 5656 367
rect 5702 333 5736 367
rect 5782 333 5816 367
rect 5862 333 5877 367
rect 5877 333 5896 367
rect 5942 333 5972 367
rect 5972 333 5976 367
rect 5244 198 5278 232
rect 5244 125 5278 159
rect 5244 51 5278 85
rect 5535 198 5569 232
rect 5535 125 5569 159
rect 5535 51 5569 85
rect 5687 93 5721 127
rect 5400 -43 5434 -9
rect 5687 -16 5721 18
rect 5999 93 6033 127
rect 5999 -16 6033 18
rect 5400 -115 5434 -81
rect 5843 -204 5877 -170
rect 5843 -276 5877 -242
rect 5301 -466 5305 -432
rect 5305 -466 5335 -432
rect 5382 -466 5400 -432
rect 5400 -466 5416 -432
rect 5462 -466 5495 -432
rect 5495 -466 5496 -432
rect 5542 -466 5576 -432
rect 5622 -466 5656 -432
rect 5702 -466 5736 -432
rect 5782 -466 5816 -432
rect 5862 -466 5877 -432
rect 5877 -466 5896 -432
rect 5942 -466 5972 -432
rect 5972 -466 5976 -432
rect 5244 -563 5278 -529
rect 5244 -636 5278 -602
rect 5244 -710 5278 -676
rect 5556 -563 5590 -529
rect 5556 -636 5590 -602
rect 5556 -710 5590 -676
rect 5687 -563 5721 -529
rect 5687 -636 5721 -602
rect 5687 -710 5721 -676
rect 5999 -563 6033 -529
rect 5999 -636 6033 -602
rect 5999 -710 6033 -676
rect 5400 -825 5434 -791
rect 5400 -897 5434 -863
rect 5843 -911 5877 -877
rect 5843 -983 5877 -949
rect 5301 -1272 5305 -1238
rect 5305 -1272 5335 -1238
rect 5382 -1272 5400 -1238
rect 5400 -1272 5416 -1238
rect 5462 -1272 5495 -1238
rect 5495 -1272 5496 -1238
rect 5542 -1272 5576 -1238
rect 5622 -1272 5656 -1238
rect 5702 -1272 5736 -1238
rect 5782 -1272 5816 -1238
rect 5862 -1272 5877 -1238
rect 5877 -1272 5896 -1238
rect 5942 -1272 5972 -1238
rect 5972 -1272 5976 -1238
rect 5244 -1357 5278 -1323
rect 5244 -1430 5278 -1396
rect 5244 -1504 5278 -1470
rect 5556 -1357 5590 -1323
rect 5556 -1430 5590 -1396
rect 5556 -1504 5590 -1470
rect 5687 -1357 5721 -1323
rect 5687 -1430 5721 -1396
rect 5687 -1504 5721 -1470
rect 5999 -1357 6033 -1323
rect 5999 -1430 6033 -1396
rect 5999 -1504 6033 -1470
rect 5400 -1621 5434 -1587
rect 5400 -1693 5434 -1659
rect 5843 -1707 5877 -1673
rect 5843 -1779 5877 -1745
rect 5301 -2068 5305 -2034
rect 5305 -2068 5335 -2034
rect 5400 -2068 5434 -2034
rect 5499 -2068 5529 -2034
rect 5529 -2068 5533 -2034
rect 5244 -2165 5278 -2131
rect 5244 -2238 5278 -2204
rect 5244 -2312 5278 -2278
rect 5556 -2165 5590 -2131
rect 5556 -2238 5590 -2204
rect 5556 -2312 5590 -2278
rect 5400 -2402 5434 -2368
rect 5400 -2474 5434 -2440
<< metal1 >>
rect 4766 11169 6251 11175
rect 4766 11135 4845 11169
rect 4879 11135 4918 11169
rect 4952 11135 4991 11169
rect 5025 11135 5064 11169
rect 5098 11135 5137 11169
rect 5171 11135 5210 11169
rect 5244 11135 5284 11169
rect 5318 11135 5358 11169
rect 5392 11135 5432 11169
rect 5466 11135 5506 11169
rect 5540 11135 5580 11169
rect 5614 11135 5654 11169
rect 5688 11135 5728 11169
rect 5762 11135 5802 11169
rect 5836 11135 5876 11169
rect 5910 11135 5950 11169
rect 5984 11135 6024 11169
rect 6058 11135 6098 11169
rect 6132 11135 6172 11169
rect 6206 11135 6251 11169
rect 4766 11097 6251 11135
rect 4766 11063 4772 11097
rect 4806 11063 4844 11097
rect 4878 11063 4918 11097
rect 4952 11063 4991 11097
rect 5025 11063 5064 11097
rect 5098 11063 5137 11097
rect 5171 11063 5210 11097
rect 5244 11063 5284 11097
rect 5318 11063 5358 11097
rect 5392 11063 5432 11097
rect 5466 11063 5506 11097
rect 5540 11063 5580 11097
rect 5614 11063 5654 11097
rect 5688 11063 5728 11097
rect 5762 11063 5802 11097
rect 5836 11063 5876 11097
rect 5910 11063 5950 11097
rect 5984 11063 6024 11097
rect 6058 11063 6098 11097
rect 6132 11063 6172 11097
rect 6206 11063 6251 11097
rect 4766 11025 6251 11063
rect 4766 11024 4916 11025
rect 4766 10990 4772 11024
rect 4806 10990 4844 11024
rect 4878 10991 4916 11024
rect 4950 10991 4989 11025
rect 5023 10991 5062 11025
rect 5096 10991 5136 11025
rect 5170 10991 5210 11025
rect 5244 10991 5284 11025
rect 5318 10991 5358 11025
rect 5392 10991 5432 11025
rect 5466 10991 5506 11025
rect 5540 10991 5580 11025
rect 5614 10991 5654 11025
rect 5688 10991 5728 11025
rect 5762 10991 5802 11025
rect 5836 10991 5876 11025
rect 5910 10991 5950 11025
rect 5984 10991 6024 11025
rect 6058 10991 6098 11025
rect 6132 10991 6172 11025
rect 6206 10991 6251 11025
rect 4878 10990 6251 10991
rect 4766 10985 6251 10990
rect 4766 10952 4956 10985
rect 4766 10951 4916 10952
rect 4766 10917 4772 10951
rect 4806 10917 4844 10951
rect 4878 10918 4916 10951
rect 4950 10918 4956 10952
rect 4878 10917 4956 10918
rect 4766 10879 4956 10917
rect 4766 10878 4916 10879
rect 4766 10844 4772 10878
rect 4806 10844 4844 10878
rect 4878 10845 4916 10878
rect 4950 10845 4956 10879
rect 4878 10844 4956 10845
rect 4766 10806 4956 10844
rect 4766 10805 4916 10806
rect 4766 10771 4772 10805
rect 4806 10771 4844 10805
rect 4878 10772 4916 10805
rect 4950 10772 4956 10806
rect 4878 10771 4956 10772
rect 4766 10733 4956 10771
rect 4766 10732 4916 10733
rect 4766 10698 4772 10732
rect 4806 10698 4844 10732
rect 4878 10699 4916 10732
rect 4950 10699 4956 10733
rect 4878 10698 4956 10699
rect 4766 10660 4956 10698
rect 4766 10659 4916 10660
rect 4766 10625 4772 10659
rect 4806 10625 4844 10659
rect 4878 10626 4916 10659
rect 4950 10626 4956 10660
rect 4878 10625 4956 10626
rect 4766 10587 4956 10625
rect 4766 10586 4916 10587
rect 4766 10552 4772 10586
rect 4806 10552 4844 10586
rect 4878 10553 4916 10586
rect 4950 10553 4956 10587
rect 4878 10552 4956 10553
rect 4766 10514 4956 10552
rect 4766 10513 4916 10514
rect 4766 10479 4772 10513
rect 4806 10479 4844 10513
rect 4878 10480 4916 10513
rect 4950 10480 4956 10514
rect 4878 10479 4956 10480
rect 4766 10441 4956 10479
rect 4766 10440 4916 10441
rect 4766 10406 4772 10440
rect 4806 10406 4844 10440
rect 4878 10407 4916 10440
rect 4950 10407 4956 10441
rect 4878 10406 4956 10407
rect 4766 10368 4956 10406
rect 4766 10367 4916 10368
rect 4766 10333 4772 10367
rect 4806 10333 4844 10367
rect 4878 10334 4916 10367
rect 4950 10334 4956 10368
rect 4878 10333 4956 10334
rect 4766 10295 4956 10333
rect 4766 10294 4916 10295
rect 4766 10260 4772 10294
rect 4806 10260 4844 10294
rect 4878 10261 4916 10294
rect 4950 10261 4956 10295
rect 4878 10260 4956 10261
rect 4766 10222 4956 10260
rect 4766 10221 4916 10222
rect 4766 10187 4772 10221
rect 4806 10187 4844 10221
rect 4878 10188 4916 10221
rect 4950 10188 4956 10222
rect 4878 10187 4956 10188
rect 4766 10149 4956 10187
rect 4766 10148 4916 10149
rect 4766 10114 4772 10148
rect 4806 10114 4844 10148
rect 4878 10115 4916 10148
rect 4950 10115 4956 10149
rect 4878 10114 4956 10115
rect 4766 10076 4956 10114
rect 4766 10075 4916 10076
rect 4766 10041 4772 10075
rect 4806 10041 4844 10075
rect 4878 10042 4916 10075
rect 4950 10042 4956 10076
rect 4878 10041 4956 10042
rect 4766 10003 4956 10041
rect 4766 10002 4916 10003
rect 4766 9968 4772 10002
rect 4806 9968 4844 10002
rect 4878 9969 4916 10002
rect 4950 9969 4956 10003
rect 4878 9968 4956 9969
rect 4766 9930 4956 9968
rect 4766 9929 4916 9930
rect 4766 9895 4772 9929
rect 4806 9895 4844 9929
rect 4878 9896 4916 9929
rect 4950 9896 4956 9930
rect 4878 9895 4956 9896
rect 4766 9857 4956 9895
rect 4766 9856 4916 9857
rect 4766 9822 4772 9856
rect 4806 9822 4844 9856
rect 4878 9823 4916 9856
rect 4950 9823 4956 9857
rect 4878 9822 4956 9823
rect 4766 9784 4956 9822
rect 4766 9783 4916 9784
rect 4766 9749 4772 9783
rect 4806 9749 4844 9783
rect 4878 9750 4916 9783
rect 4950 9750 4956 9784
rect 4878 9749 4956 9750
rect 4766 9711 4956 9749
rect 4766 9710 4916 9711
rect 4766 9676 4772 9710
rect 4806 9676 4844 9710
rect 4878 9677 4916 9710
rect 4950 9677 4956 9711
rect 4878 9676 4956 9677
rect 4766 9638 4956 9676
rect 4766 9637 4916 9638
rect 4766 9603 4772 9637
rect 4806 9603 4844 9637
rect 4878 9604 4916 9637
rect 4950 9604 4956 9638
rect 4878 9603 4956 9604
rect 4766 9565 4956 9603
rect 4766 9564 4916 9565
rect 4766 9530 4772 9564
rect 4806 9530 4844 9564
rect 4878 9531 4916 9564
rect 4950 9531 4956 9565
rect 4878 9530 4956 9531
rect 4766 9492 4956 9530
rect 4766 9491 4916 9492
rect 4766 9457 4772 9491
rect 4806 9457 4844 9491
rect 4878 9458 4916 9491
rect 4950 9458 4956 9492
rect 4878 9457 4956 9458
rect 4766 9419 4956 9457
rect 4766 9418 4916 9419
rect 4766 9384 4772 9418
rect 4806 9384 4844 9418
rect 4878 9385 4916 9418
rect 4950 9385 4956 9419
rect 4878 9384 4956 9385
rect 4766 9346 4956 9384
rect 4766 9345 4916 9346
rect 4766 9311 4772 9345
rect 4806 9311 4844 9345
rect 4878 9312 4916 9345
rect 4950 9312 4956 9346
rect 4878 9311 4956 9312
rect 4766 9273 4956 9311
rect 4766 9272 4916 9273
rect 4766 9238 4772 9272
rect 4806 9238 4844 9272
rect 4878 9239 4916 9272
rect 4950 9239 4956 9273
rect 4878 9238 4956 9239
rect 4766 9200 4956 9238
rect 4766 9199 4916 9200
rect 4766 9165 4772 9199
rect 4806 9165 4844 9199
rect 4878 9166 4916 9199
rect 4950 9166 4956 9200
rect 4878 9165 4956 9166
rect 4766 9127 4956 9165
rect 4766 9126 4916 9127
rect 4766 9092 4772 9126
rect 4806 9092 4844 9126
rect 4878 9093 4916 9126
rect 4950 9093 4956 9127
rect 4878 9092 4956 9093
rect 4766 9054 4956 9092
rect 4766 9053 4916 9054
rect 4766 9019 4772 9053
rect 4806 9019 4844 9053
rect 4878 9020 4916 9053
rect 4950 9020 4956 9054
rect 4878 9019 4956 9020
rect 4766 8981 4956 9019
rect 4766 8980 4916 8981
rect 4766 8946 4772 8980
rect 4806 8946 4844 8980
rect 4878 8947 4916 8980
rect 4950 8947 4956 8981
rect 4878 8946 4956 8947
rect 4766 8908 4956 8946
rect 4766 8907 4916 8908
rect 4766 8873 4772 8907
rect 4806 8873 4844 8907
rect 4878 8874 4916 8907
rect 4950 8874 4956 8908
rect 4878 8873 4956 8874
rect 4766 8835 4956 8873
rect 4766 8834 4916 8835
rect 4766 4264 4772 8834
rect 4878 8801 4916 8834
rect 4950 8801 4956 8835
rect 4878 8762 4956 8801
rect 4950 4376 4956 8762
rect 5090 10845 5832 10851
rect 5090 10811 5174 10845
rect 5208 10811 5252 10845
rect 5286 10817 5330 10845
rect 5364 10817 5408 10845
rect 5442 10817 5486 10845
rect 5364 10811 5374 10817
rect 5442 10811 5467 10817
rect 5520 10811 5564 10845
rect 5598 10811 5642 10845
rect 5676 10811 5720 10845
rect 5754 10811 5832 10845
rect 5090 10773 5281 10811
rect 5333 10773 5374 10811
rect 5426 10773 5467 10811
rect 5519 10773 5832 10811
rect 5090 10739 5096 10773
rect 5130 10739 5168 10773
rect 5202 10739 5252 10773
rect 5364 10765 5374 10773
rect 5442 10765 5467 10773
rect 5286 10739 5330 10765
rect 5364 10739 5408 10765
rect 5442 10739 5486 10765
rect 5520 10739 5564 10773
rect 5598 10739 5642 10773
rect 5676 10739 5720 10773
rect 5090 10733 5720 10739
rect 5090 10700 5208 10733
rect 5090 10666 5096 10700
rect 5130 10666 5168 10700
rect 5202 10666 5208 10700
rect 5090 10627 5208 10666
rect 5090 10593 5096 10627
rect 5130 10593 5168 10627
rect 5202 10593 5208 10627
rect 5714 10667 5720 10733
rect 5826 10667 5832 10773
rect 5714 10628 5832 10667
rect 5714 10594 5720 10628
rect 5754 10594 5792 10628
rect 5826 10594 5832 10628
rect 5090 10554 5208 10593
rect 5090 10520 5096 10554
rect 5130 10520 5168 10554
rect 5202 10520 5208 10554
rect 5090 10481 5208 10520
rect 5090 10447 5096 10481
rect 5130 10447 5168 10481
rect 5202 10447 5208 10481
tri 5357 10591 5360 10594 se
rect 5360 10591 5406 10594
tri 5406 10591 5409 10594 sw
rect 5357 10585 5409 10591
rect 5357 10521 5409 10533
rect 5357 10465 5366 10469
rect 5400 10465 5409 10469
rect 5357 10456 5409 10465
tri 5357 10453 5360 10456 ne
rect 5090 10408 5208 10447
rect 5090 10374 5096 10408
rect 5130 10374 5168 10408
rect 5202 10374 5208 10408
rect 5090 10335 5208 10374
rect 5090 10301 5096 10335
rect 5130 10301 5168 10335
rect 5202 10301 5208 10335
rect 5090 10262 5208 10301
rect 5090 10228 5096 10262
rect 5130 10228 5168 10262
rect 5202 10228 5208 10262
rect 5090 10189 5208 10228
rect 5090 10155 5096 10189
rect 5130 10155 5168 10189
rect 5202 10155 5208 10189
rect 5090 10116 5208 10155
rect 5090 4610 5096 10116
rect 5202 4683 5208 10116
tri 5279 10091 5282 10094 se
rect 5282 10091 5328 10094
tri 5328 10091 5331 10094 sw
rect 5279 10085 5331 10091
rect 5279 10021 5331 10033
rect 5279 9957 5331 9969
rect 5279 9883 5331 9905
rect 5360 9886 5406 10456
tri 5406 10453 5409 10456 nw
tri 5513 10591 5516 10594 se
rect 5516 10591 5562 10594
tri 5562 10591 5565 10594 sw
rect 5513 10585 5565 10591
rect 5513 10521 5565 10533
rect 5513 10465 5522 10469
rect 5556 10465 5565 10469
rect 5513 10456 5565 10465
tri 5513 10453 5516 10456 ne
rect 5435 10423 5487 10445
rect 5435 10359 5487 10371
rect 5435 10295 5487 10307
rect 5435 10237 5487 10243
tri 5435 10234 5438 10237 ne
rect 5438 10234 5484 10237
tri 5484 10234 5487 10237 nw
rect 5360 9852 5366 9886
rect 5400 9852 5406 9886
rect 5360 9814 5406 9852
rect 5279 9761 5331 9783
rect 5279 9697 5331 9709
rect 5279 9633 5331 9645
rect 5279 9575 5331 9581
tri 5279 9572 5282 9575 ne
rect 5282 9572 5328 9575
tri 5328 9572 5331 9575 nw
rect 5360 9780 5366 9814
rect 5400 9780 5406 9814
rect 5360 9154 5406 9780
rect 5516 9886 5562 10456
tri 5562 10453 5565 10456 nw
rect 5714 10555 5832 10594
rect 5714 10521 5720 10555
rect 5754 10521 5792 10555
rect 5826 10521 5832 10555
rect 5714 10482 5832 10521
rect 5714 10448 5720 10482
rect 5754 10448 5792 10482
rect 5826 10448 5832 10482
rect 5714 10409 5832 10448
rect 5714 10375 5720 10409
rect 5754 10375 5792 10409
rect 5826 10375 5832 10409
rect 5714 10336 5832 10375
rect 5714 10302 5720 10336
rect 5754 10302 5792 10336
rect 5826 10302 5832 10336
rect 5714 10263 5832 10302
rect 5714 10229 5720 10263
rect 5754 10229 5792 10263
rect 5826 10229 5832 10263
rect 5714 10190 5832 10229
rect 5714 10156 5720 10190
rect 5754 10156 5792 10190
rect 5826 10156 5832 10190
rect 5714 10117 5832 10156
rect 5516 9852 5522 9886
rect 5556 9852 5562 9886
tri 5591 10091 5594 10094 se
rect 5594 10091 5640 10094
tri 5640 10091 5643 10094 sw
rect 5591 10085 5643 10091
rect 5591 10021 5643 10033
rect 5591 9957 5643 9969
rect 5591 9883 5643 9905
rect 5714 10083 5720 10117
rect 5754 10083 5792 10117
rect 5826 10083 5832 10117
rect 5714 10044 5832 10083
rect 5714 10010 5720 10044
rect 5754 10010 5792 10044
rect 5826 10010 5832 10044
rect 5714 9971 5832 10010
rect 5714 9937 5720 9971
rect 5754 9937 5792 9971
rect 5826 9937 5832 9971
rect 5714 9898 5832 9937
rect 5516 9814 5562 9852
rect 5516 9780 5522 9814
rect 5556 9780 5562 9814
rect 5714 9864 5720 9898
rect 5754 9864 5792 9898
rect 5826 9864 5832 9898
rect 5714 9825 5832 9864
rect 5714 9791 5720 9825
rect 5754 9791 5792 9825
rect 5826 9791 5832 9825
tri 5435 9429 5438 9432 se
rect 5438 9429 5484 9432
tri 5484 9429 5487 9432 sw
rect 5435 9423 5487 9429
rect 5435 9359 5487 9371
rect 5435 9295 5487 9307
rect 5435 9221 5487 9243
rect 5360 9120 5366 9154
rect 5400 9120 5406 9154
rect 5360 9082 5406 9120
rect 5360 9048 5366 9082
rect 5400 9048 5406 9082
tri 5279 8627 5282 8630 se
rect 5282 8627 5328 8630
tri 5328 8627 5331 8630 sw
rect 5279 8621 5331 8627
rect 5279 8557 5331 8569
rect 5279 8493 5331 8505
rect 5279 8419 5331 8441
rect 5360 8422 5406 9048
rect 5516 9154 5562 9780
rect 5591 9761 5643 9783
rect 5591 9697 5643 9709
rect 5591 9633 5643 9645
rect 5591 9575 5643 9581
tri 5591 9572 5594 9575 ne
rect 5594 9572 5640 9575
tri 5640 9572 5643 9575 nw
rect 5714 9752 5832 9791
rect 5714 9718 5720 9752
rect 5754 9718 5792 9752
rect 5826 9718 5832 9752
rect 5714 9679 5832 9718
rect 5714 9645 5720 9679
rect 5754 9645 5792 9679
rect 5826 9645 5832 9679
rect 5714 9606 5832 9645
rect 5714 9572 5720 9606
rect 5754 9572 5792 9606
rect 5826 9572 5832 9606
rect 5516 9120 5522 9154
rect 5556 9120 5562 9154
rect 5516 9082 5562 9120
rect 5516 9048 5522 9082
rect 5556 9048 5562 9082
rect 5435 8959 5487 8981
rect 5435 8895 5487 8907
rect 5435 8831 5487 8843
rect 5435 8773 5487 8779
tri 5435 8770 5438 8773 ne
rect 5438 8770 5484 8773
tri 5484 8770 5487 8773 nw
rect 5360 8388 5366 8422
rect 5400 8388 5406 8422
rect 5360 8350 5406 8388
rect 5279 8297 5331 8319
rect 5279 8233 5331 8245
rect 5279 8169 5331 8181
rect 5279 8111 5331 8117
tri 5279 8108 5282 8111 ne
rect 5282 8108 5328 8111
tri 5328 8108 5331 8111 nw
rect 5360 8316 5366 8350
rect 5400 8316 5406 8350
rect 5360 7690 5406 8316
rect 5516 8422 5562 9048
rect 5714 9533 5832 9572
rect 5714 9499 5720 9533
rect 5754 9499 5792 9533
rect 5826 9499 5832 9533
rect 5714 9460 5832 9499
rect 5714 9426 5720 9460
rect 5754 9426 5792 9460
rect 5826 9426 5832 9460
rect 5714 9387 5832 9426
rect 5714 9353 5720 9387
rect 5754 9353 5792 9387
rect 5826 9353 5832 9387
rect 5714 9314 5832 9353
rect 5714 9280 5720 9314
rect 5754 9280 5792 9314
rect 5826 9280 5832 9314
rect 5714 9216 5832 9280
rect 5714 9182 5720 9216
rect 5754 9182 5792 9216
rect 5826 9182 5832 9216
rect 5714 9143 5832 9182
rect 5714 9109 5720 9143
rect 5754 9109 5792 9143
rect 5826 9109 5832 9143
rect 5714 9070 5832 9109
rect 5714 9036 5720 9070
rect 5754 9036 5792 9070
rect 5826 9036 5832 9070
rect 5714 8997 5832 9036
rect 5714 8963 5720 8997
rect 5754 8963 5792 8997
rect 5826 8963 5832 8997
rect 5714 8924 5832 8963
rect 5714 8890 5720 8924
rect 5754 8890 5792 8924
rect 5826 8890 5832 8924
rect 5714 8851 5832 8890
rect 5714 8817 5720 8851
rect 5754 8817 5792 8851
rect 5826 8817 5832 8851
rect 5714 8778 5832 8817
rect 5714 8744 5720 8778
rect 5754 8744 5792 8778
rect 5826 8744 5832 8778
rect 5714 8705 5832 8744
rect 5714 8671 5720 8705
rect 5754 8671 5792 8705
rect 5826 8671 5832 8705
rect 5714 8632 5832 8671
rect 5516 8388 5522 8422
rect 5556 8388 5562 8422
tri 5591 8627 5594 8630 se
rect 5594 8627 5640 8630
tri 5640 8627 5643 8630 sw
rect 5591 8621 5643 8627
rect 5591 8557 5643 8569
rect 5591 8493 5643 8505
rect 5591 8419 5643 8441
rect 5714 8598 5720 8632
rect 5754 8598 5792 8632
rect 5826 8598 5832 8632
rect 5714 8559 5832 8598
rect 5714 8525 5720 8559
rect 5754 8525 5792 8559
rect 5826 8525 5832 8559
rect 5714 8486 5832 8525
rect 5714 8452 5720 8486
rect 5754 8452 5792 8486
rect 5826 8452 5832 8486
rect 5516 8350 5562 8388
rect 5516 8316 5522 8350
rect 5556 8316 5562 8350
rect 5714 8413 5832 8452
rect 5714 8379 5720 8413
rect 5754 8379 5792 8413
rect 5826 8379 5832 8413
rect 5714 8340 5832 8379
tri 5435 7965 5438 7968 se
rect 5438 7965 5484 7968
tri 5484 7965 5487 7968 sw
rect 5435 7959 5487 7965
rect 5435 7895 5487 7907
rect 5435 7831 5487 7843
rect 5435 7757 5487 7779
rect 5360 7656 5366 7690
rect 5400 7656 5406 7690
rect 5360 7618 5406 7656
rect 5360 7584 5366 7618
rect 5400 7584 5406 7618
tri 5279 7163 5282 7166 se
rect 5282 7163 5328 7166
tri 5328 7163 5331 7166 sw
rect 5279 7157 5331 7163
rect 5279 7093 5331 7105
rect 5279 7029 5331 7041
rect 5279 6955 5331 6977
rect 5360 6958 5406 7584
rect 5516 7690 5562 8316
rect 5591 8297 5643 8319
rect 5591 8233 5643 8245
rect 5591 8169 5643 8181
rect 5591 8111 5643 8117
tri 5591 8108 5594 8111 ne
rect 5594 8108 5640 8111
tri 5640 8108 5643 8111 nw
rect 5714 8306 5720 8340
rect 5754 8306 5792 8340
rect 5826 8306 5832 8340
rect 5714 8267 5832 8306
rect 5714 8233 5720 8267
rect 5754 8233 5792 8267
rect 5826 8233 5832 8267
rect 5714 8194 5832 8233
rect 5714 8160 5720 8194
rect 5754 8160 5792 8194
rect 5826 8160 5832 8194
rect 5714 8121 5832 8160
rect 5516 7656 5522 7690
rect 5556 7656 5562 7690
rect 5516 7618 5562 7656
rect 5516 7584 5522 7618
rect 5556 7584 5562 7618
rect 5435 7495 5487 7517
rect 5435 7431 5487 7443
rect 5435 7367 5487 7379
rect 5435 7309 5487 7315
tri 5435 7306 5438 7309 ne
rect 5438 7306 5484 7309
tri 5484 7306 5487 7309 nw
rect 5360 6924 5366 6958
rect 5400 6924 5406 6958
rect 5360 6886 5406 6924
rect 5279 6833 5331 6855
rect 5279 6769 5331 6781
rect 5279 6705 5331 6717
rect 5279 6647 5331 6653
tri 5279 6644 5282 6647 ne
rect 5282 6644 5328 6647
tri 5328 6644 5331 6647 nw
rect 5360 6852 5366 6886
rect 5400 6852 5406 6886
rect 5360 6226 5406 6852
rect 5516 6958 5562 7584
rect 5714 8087 5720 8121
rect 5754 8087 5792 8121
rect 5826 8087 5832 8121
rect 5714 8048 5832 8087
rect 5714 8014 5720 8048
rect 5754 8014 5792 8048
rect 5826 8014 5832 8048
rect 5714 7975 5832 8014
rect 5714 7941 5720 7975
rect 5754 7941 5792 7975
rect 5826 7941 5832 7975
rect 5714 7902 5832 7941
rect 5714 7868 5720 7902
rect 5754 7868 5792 7902
rect 5826 7868 5832 7902
rect 5714 7829 5832 7868
rect 5714 7795 5720 7829
rect 5754 7795 5792 7829
rect 5826 7795 5832 7829
rect 5714 7756 5832 7795
rect 5714 7722 5720 7756
rect 5754 7722 5792 7756
rect 5826 7722 5832 7756
rect 5714 7683 5832 7722
rect 5714 7649 5720 7683
rect 5754 7649 5792 7683
rect 5826 7649 5832 7683
rect 5714 7610 5832 7649
rect 5714 7576 5720 7610
rect 5754 7576 5792 7610
rect 5826 7576 5832 7610
rect 5714 7537 5832 7576
rect 5714 7503 5720 7537
rect 5754 7503 5792 7537
rect 5826 7503 5832 7537
rect 5714 7464 5832 7503
rect 5714 7430 5720 7464
rect 5754 7430 5792 7464
rect 5826 7430 5832 7464
rect 5714 7391 5832 7430
rect 5714 7357 5720 7391
rect 5754 7357 5792 7391
rect 5826 7357 5832 7391
rect 5714 7318 5832 7357
rect 5714 7284 5720 7318
rect 5754 7284 5792 7318
rect 5826 7284 5832 7318
rect 5714 7245 5832 7284
rect 5714 7211 5720 7245
rect 5754 7211 5792 7245
rect 5826 7211 5832 7245
rect 5714 7172 5832 7211
rect 5516 6924 5522 6958
rect 5556 6924 5562 6958
tri 5591 7163 5594 7166 se
rect 5594 7163 5640 7166
tri 5640 7163 5643 7166 sw
rect 5591 7157 5643 7163
rect 5591 7093 5643 7105
rect 5591 7029 5643 7041
rect 5591 6955 5643 6977
rect 5714 7138 5720 7172
rect 5754 7138 5792 7172
rect 5826 7138 5832 7172
rect 5714 7099 5832 7138
rect 5714 7065 5720 7099
rect 5754 7065 5792 7099
rect 5826 7065 5832 7099
rect 5714 7026 5832 7065
rect 5714 6992 5720 7026
rect 5754 6992 5792 7026
rect 5826 6992 5832 7026
rect 5516 6886 5562 6924
rect 5516 6852 5522 6886
rect 5556 6852 5562 6886
rect 5714 6953 5832 6992
rect 5714 6919 5720 6953
rect 5754 6919 5792 6953
rect 5826 6919 5832 6953
rect 5714 6880 5832 6919
tri 5435 6501 5438 6504 se
rect 5438 6501 5484 6504
tri 5484 6501 5487 6504 sw
rect 5435 6495 5487 6501
rect 5435 6431 5487 6443
rect 5435 6367 5487 6379
rect 5435 6293 5487 6315
rect 5360 6192 5366 6226
rect 5400 6192 5406 6226
rect 5360 6154 5406 6192
rect 5360 6120 5366 6154
rect 5400 6120 5406 6154
rect 5360 6108 5406 6120
rect 5516 6226 5562 6852
rect 5591 6833 5643 6855
rect 5591 6769 5643 6781
rect 5591 6705 5643 6717
rect 5591 6647 5643 6653
tri 5591 6644 5594 6647 ne
rect 5594 6644 5640 6647
tri 5640 6644 5643 6647 nw
rect 5714 6846 5720 6880
rect 5754 6846 5792 6880
rect 5826 6846 5832 6880
rect 5714 6807 5832 6846
rect 5714 6773 5720 6807
rect 5754 6773 5792 6807
rect 5826 6773 5832 6807
rect 5714 6734 5832 6773
rect 5714 6700 5720 6734
rect 5754 6700 5792 6734
rect 5826 6700 5832 6734
rect 5714 6661 5832 6700
rect 5516 6192 5522 6226
rect 5556 6192 5562 6226
rect 5516 6154 5562 6192
rect 5516 6120 5522 6154
rect 5556 6120 5562 6154
rect 5516 6108 5562 6120
rect 5435 6031 5487 6053
rect 5435 5967 5487 5979
rect 5435 5903 5487 5915
rect 5435 5845 5487 5851
tri 5435 5842 5438 5845 ne
rect 5438 5842 5484 5845
tri 5484 5842 5487 5845 nw
tri 5279 5699 5282 5702 se
rect 5282 5699 5328 5702
tri 5328 5699 5331 5702 sw
tri 5591 5699 5594 5702 se
rect 5594 5699 5640 5702
tri 5640 5699 5643 5702 sw
rect 5279 5693 5331 5699
rect 5279 5629 5331 5641
rect 5279 5565 5331 5577
rect 5279 5491 5331 5513
rect 5525 5693 5643 5699
rect 5577 5641 5643 5693
rect 5525 5629 5643 5641
rect 5577 5577 5643 5629
rect 5525 5565 5643 5577
rect 5577 5513 5643 5565
rect 5525 5507 5643 5513
tri 5575 5491 5591 5507 ne
rect 5591 5491 5643 5507
tri 5208 4683 5245 4720 sw
tri 5677 4683 5714 4720 se
rect 5714 4683 5720 6661
rect 5826 4683 5832 6661
rect 5202 4650 5245 4683
tri 5245 4650 5278 4683 sw
tri 5644 4650 5677 4683 se
rect 5677 4650 5832 4683
rect 5202 4644 5832 4650
rect 5202 4610 5244 4644
rect 5278 4610 5320 4644
rect 5354 4610 5395 4644
rect 5429 4610 5470 4644
rect 5504 4610 5545 4644
rect 5579 4610 5620 4644
rect 5654 4610 5695 4644
rect 5729 4610 5832 4644
rect 5090 4595 5832 4610
rect 5090 4572 5792 4595
rect 5090 4538 5168 4572
rect 5202 4538 5246 4572
rect 5280 4538 5324 4572
rect 5358 4538 5402 4572
rect 5436 4538 5480 4572
rect 5514 4538 5558 4572
rect 5592 4538 5636 4572
rect 5670 4538 5714 4572
rect 5748 4561 5792 4572
rect 5826 4561 5832 4595
rect 5748 4538 5832 4561
rect 5090 4532 5832 4538
tri 6165 4376 6243 4454 se
rect 4950 4370 6251 4376
rect 4950 4336 4990 4370
rect 5024 4336 5064 4370
rect 5098 4336 5138 4370
rect 5172 4336 5212 4370
rect 5246 4336 5286 4370
rect 5320 4336 5360 4370
rect 5394 4336 5434 4370
rect 5468 4336 5508 4370
rect 5542 4336 5582 4370
rect 5616 4336 5656 4370
rect 5690 4336 5730 4370
rect 5764 4336 5804 4370
rect 5838 4336 5878 4370
rect 5912 4336 5952 4370
rect 5986 4336 6026 4370
rect 6060 4336 6099 4370
rect 6133 4336 6172 4370
rect 6206 4336 6251 4370
rect 4878 4298 6251 4336
rect 4878 4264 4918 4298
rect 4952 4264 4992 4298
rect 5026 4264 5066 4298
rect 5100 4264 5140 4298
rect 5174 4264 5214 4298
rect 5248 4264 5288 4298
rect 5322 4264 5362 4298
rect 5396 4264 5436 4298
rect 5470 4264 5510 4298
rect 5544 4264 5584 4298
rect 5618 4264 5658 4298
rect 5692 4264 5732 4298
rect 5766 4264 5806 4298
rect 5840 4264 5880 4298
rect 5914 4264 5953 4298
rect 5987 4264 6026 4298
rect 6060 4264 6099 4298
rect 6133 4264 6172 4298
rect 6206 4264 6251 4298
rect 4766 4226 6251 4264
rect 4766 4192 4844 4226
rect 4878 4192 4918 4226
rect 4952 4192 4992 4226
rect 5026 4192 5066 4226
rect 5100 4192 5140 4226
rect 5174 4192 5214 4226
rect 5248 4192 5288 4226
rect 5322 4192 5362 4226
rect 5396 4192 5436 4226
rect 5470 4192 5510 4226
rect 5544 4192 5584 4226
rect 5618 4192 5658 4226
rect 5692 4192 5732 4226
rect 5766 4192 5806 4226
rect 5840 4192 5880 4226
rect 5914 4192 5953 4226
rect 5987 4192 6026 4226
rect 6060 4192 6099 4226
rect 6133 4192 6172 4226
rect 6206 4192 6251 4226
rect 4766 4186 6251 4192
tri 6165 4108 6243 4186 ne
rect 6204 3227 6327 3233
rect 6204 3175 6211 3227
rect 6263 3175 6275 3227
tri 6327 3206 6354 3233 sw
rect 6327 3175 21455 3206
rect 6204 3152 21455 3175
rect 6204 3100 6211 3152
rect 6263 3100 6275 3152
rect 6327 3100 21455 3152
rect 6204 3094 21455 3100
tri 21269 3026 21337 3094 ne
rect 5928 2871 5980 2877
rect 5928 2796 5980 2819
tri 5913 2760 5928 2775 se
tri 5249 2688 5321 2760 se
rect 5321 2744 5928 2760
rect 5321 2738 5980 2744
rect 6020 2818 6072 2824
rect 6020 2743 6072 2766
rect 5321 2708 5949 2738
tri 5949 2708 5979 2738 nw
rect 5321 2688 5332 2708
tri 5332 2688 5352 2708 nw
rect 5249 2683 5327 2688
tri 5327 2683 5332 2688 nw
rect 5249 2668 5312 2683
tri 5312 2668 5327 2683 nw
tri 6005 2668 6020 2683 se
rect 6020 2668 6072 2691
rect 5249 2480 5301 2668
tri 5301 2657 5312 2668 nw
tri 5402 2657 5413 2668 se
rect 5413 2657 6072 2668
rect 5249 2405 5301 2428
rect 5249 2347 5301 2353
tri 5341 2596 5402 2657 se
rect 5402 2647 6072 2657
rect 5402 2616 6041 2647
tri 6041 2616 6072 2647 nw
rect 6112 2818 6164 2824
rect 6112 2743 6164 2766
rect 5402 2596 5424 2616
tri 5424 2596 5444 2616 nw
rect 5341 2595 5423 2596
tri 5423 2595 5424 2596 nw
rect 5341 2580 5408 2595
tri 5408 2580 5423 2595 nw
tri 6097 2580 6112 2595 se
rect 6112 2580 6164 2691
rect 5341 2480 5393 2580
tri 5393 2565 5408 2580 nw
tri 5490 2565 5505 2580 se
rect 5505 2565 6164 2580
rect 5341 2405 5393 2428
rect 5341 2347 5393 2353
tri 5433 2508 5490 2565 se
rect 5490 2557 6164 2565
rect 5490 2528 6135 2557
tri 6135 2528 6164 2557 nw
rect 5490 2508 5516 2528
tri 5516 2508 5536 2528 nw
rect 5433 2478 5485 2508
tri 5485 2477 5516 2508 nw
rect 5433 2403 5485 2426
rect 5433 2345 5485 2351
rect 5525 2211 5577 2217
rect 5525 2147 5577 2159
rect 21337 2154 21455 3094
rect 25918 2210 25970 2219
tri 25970 2210 25979 2219 sw
rect 20805 2133 20811 2141
rect 5577 2095 20811 2133
rect 5525 2089 20811 2095
rect 20863 2089 20875 2141
rect 20927 2089 20933 2141
rect 21337 2038 21338 2154
rect 21454 2038 21455 2154
rect 21337 2027 21455 2038
tri 25670 2142 25678 2150 se
rect 25678 2142 25730 2207
rect 25670 2136 25730 2142
rect 25722 2135 25730 2136
tri 25722 2127 25730 2135 nw
rect 25758 2142 25810 2207
rect 25838 2182 25890 2207
rect 25918 2204 25979 2210
tri 25918 2195 25927 2204 ne
rect 25927 2201 25979 2204
tri 25890 2182 25899 2191 sw
rect 25838 2176 25899 2182
tri 25838 2167 25847 2176 ne
rect 25847 2175 25899 2176
tri 25810 2142 25818 2150 sw
rect 25758 2136 25818 2142
rect 25758 2135 25766 2136
tri 25758 2127 25766 2135 ne
rect 25670 2072 25722 2084
rect 25670 2014 25722 2020
rect 25766 2072 25818 2084
rect 25847 2111 25899 2123
rect 25927 2137 25979 2149
rect 25927 2079 25979 2085
tri 26856 2160 26876 2180 se
rect 26876 2160 26973 2180
rect 25847 2053 25899 2059
rect 26856 2063 26973 2160
rect 26856 2053 26963 2063
tri 26963 2053 26973 2063 nw
rect 25766 2014 25818 2020
tri 26799 1934 26856 1991 se
rect 26856 1934 26933 2053
tri 26933 2023 26963 2053 nw
rect 25511 1818 25517 1934
rect 25633 1818 26209 1934
rect 26326 1861 26933 1934
rect 26326 1818 26890 1861
tri 26890 1818 26933 1861 nw
rect 20805 1516 20811 1568
rect 20863 1516 20875 1568
rect 20927 1561 20933 1568
rect 26003 1561 26009 1569
rect 20927 1517 26009 1561
rect 26061 1517 26073 1569
rect 26125 1517 26131 1569
rect 20927 1516 20933 1517
rect 5618 1485 5624 1493
rect 5617 1441 5624 1485
rect 5676 1441 5688 1493
rect 5740 1485 5746 1493
rect 26179 1485 26185 1493
rect 5740 1441 26185 1485
rect 26237 1441 26249 1493
rect 26301 1441 26307 1493
rect 25886 1180 25892 1188
rect 5709 1174 25892 1180
rect 5761 1136 25892 1174
rect 25944 1136 25956 1188
rect 26008 1136 26014 1188
rect 5709 1110 5761 1122
rect 5709 1052 5761 1058
rect 5801 1054 5807 1106
rect 5859 1054 5871 1106
rect 5923 1104 5929 1106
rect 26056 1104 26062 1112
rect 5923 1060 26062 1104
rect 26114 1060 26126 1112
rect 26178 1060 26184 1112
rect 5923 1054 5929 1060
rect 5289 367 6008 373
rect 5289 333 5301 367
rect 5335 333 5382 367
rect 5416 333 5462 367
rect 5496 333 5542 367
rect 5576 333 5622 367
rect 5656 333 5702 367
rect 5736 333 5782 367
rect 5816 333 5862 367
rect 5896 333 5942 367
rect 5976 333 6008 367
rect 5289 327 6008 333
tri 6008 327 6054 373 sw
tri 5988 317 5998 327 ne
rect 5998 317 6054 327
tri 6054 317 6064 327 sw
tri 5998 279 6036 317 ne
rect 6036 279 6252 317
rect 6246 265 6252 279
rect 6304 265 6316 317
rect 6368 265 6374 317
rect 5238 238 5577 244
rect 5238 232 5525 238
rect 5238 198 5244 232
rect 5278 198 5525 232
rect 5238 186 5525 198
rect 5238 168 5577 186
rect 5238 159 5525 168
rect 5238 125 5244 159
rect 5278 125 5525 159
rect 5238 116 5525 125
rect 5238 97 5577 116
rect 5238 85 5525 97
rect 5238 51 5244 85
rect 5278 51 5525 85
rect 5238 45 5525 51
rect 5238 39 5577 45
rect 5617 133 6039 139
rect 5669 127 6039 133
rect 5669 93 5687 127
rect 5721 93 5999 127
rect 6033 93 6039 127
rect 5669 81 6039 93
rect 5617 30 6039 81
rect 5149 23 5201 29
rect 5149 -41 5201 -29
rect 5149 -99 5201 -93
rect 5394 -9 5440 3
rect 5394 -43 5400 -9
rect 5434 -43 5440 -9
rect 5669 18 6039 30
rect 5669 -16 5687 18
rect 5721 -16 5999 18
rect 6033 -16 6039 18
rect 5669 -22 6039 -16
rect 5617 -28 6039 -22
rect 5394 -81 5440 -43
rect 5394 -115 5400 -81
rect 5434 -115 5440 -81
rect 5394 -127 5440 -115
rect 5148 -164 5200 -158
rect 5148 -228 5200 -216
rect 5148 -286 5200 -280
rect 5837 -170 5883 -158
rect 5837 -204 5843 -170
rect 5877 -204 5883 -170
rect 5837 -242 5883 -204
rect 5837 -276 5843 -242
rect 5877 -276 5883 -242
rect 5837 -288 5883 -276
rect 5289 -432 6086 -426
rect 5289 -466 5301 -432
rect 5335 -466 5382 -432
rect 5416 -466 5462 -432
rect 5496 -466 5542 -432
rect 5576 -466 5622 -432
rect 5656 -466 5702 -432
rect 5736 -466 5782 -432
rect 5816 -466 5862 -432
rect 5896 -466 5942 -432
rect 5976 -466 6086 -432
rect 5289 -469 6086 -466
tri 6086 -469 6129 -426 sw
rect 5289 -472 6471 -469
tri 6050 -507 6085 -472 ne
rect 6085 -475 6471 -472
rect 6085 -507 6419 -475
rect 5238 -523 5596 -517
rect 5238 -529 5525 -523
rect 5577 -529 5596 -523
rect 5238 -563 5244 -529
rect 5278 -563 5525 -529
rect 5590 -563 5596 -529
rect 5238 -575 5525 -563
rect 5577 -575 5596 -563
rect 5238 -593 5596 -575
rect 5238 -602 5525 -593
rect 5577 -602 5596 -593
rect 5238 -636 5244 -602
rect 5278 -636 5525 -602
rect 5590 -636 5596 -602
rect 5238 -645 5525 -636
rect 5577 -645 5596 -636
rect 5238 -664 5596 -645
rect 5238 -676 5525 -664
rect 5577 -676 5596 -664
rect 5148 -707 5200 -701
rect 5238 -710 5244 -676
rect 5278 -710 5525 -676
rect 5590 -710 5596 -676
rect 5238 -716 5525 -710
rect 5577 -716 5596 -710
rect 5238 -722 5596 -716
rect 5681 -523 6039 -517
rect 5681 -529 5801 -523
rect 5681 -563 5687 -529
rect 5721 -563 5801 -529
rect 5681 -575 5801 -563
rect 5853 -529 6039 -523
rect 5853 -563 5999 -529
rect 6033 -563 6039 -529
rect 5853 -575 6039 -563
rect 5681 -593 6039 -575
rect 5681 -602 5801 -593
rect 5681 -636 5687 -602
rect 5721 -636 5801 -602
rect 5681 -645 5801 -636
rect 5853 -602 6039 -593
rect 6419 -539 6471 -527
rect 6419 -597 6471 -591
rect 5853 -636 5999 -602
rect 6033 -636 6039 -602
rect 5853 -645 6039 -636
rect 5681 -664 6039 -645
rect 5681 -676 5801 -664
rect 5681 -710 5687 -676
rect 5721 -710 5801 -676
rect 5681 -716 5801 -710
rect 5853 -676 6039 -664
rect 5853 -710 5999 -676
rect 6033 -710 6039 -676
rect 5853 -716 6039 -710
rect 5681 -722 6039 -716
rect 5148 -771 5200 -759
rect 6009 -774 6061 -768
rect 5200 -791 6009 -779
rect 5200 -823 5400 -791
rect 5148 -825 5400 -823
rect 5434 -825 6009 -791
rect 5148 -826 6009 -825
rect 6061 -826 6715 -779
rect 5148 -829 6715 -826
rect 5394 -863 5440 -829
rect 5394 -897 5400 -863
rect 5434 -897 5440 -863
rect 6009 -838 6061 -829
rect 5394 -909 5440 -897
rect 5837 -877 5883 -865
rect 5837 -911 5843 -877
rect 5877 -911 5883 -877
rect 6009 -896 6061 -890
rect 6575 -891 6627 -885
rect 5837 -946 5883 -911
rect 6575 -946 6627 -943
rect 5163 -949 6627 -946
rect 5163 -952 5843 -949
rect 5215 -983 5843 -952
rect 5877 -955 6627 -949
rect 5877 -983 6575 -955
rect 5215 -996 6575 -983
rect 5163 -1016 5215 -1004
rect 6575 -1013 6627 -1007
rect 5163 -1074 5215 -1068
rect 5341 -1066 5730 -1060
rect 5393 -1118 5678 -1066
rect 5341 -1133 5393 -1118
tri 5393 -1142 5417 -1118 nw
tri 5649 -1142 5673 -1118 ne
rect 5673 -1133 5730 -1118
rect 5673 -1142 5678 -1133
tri 5673 -1147 5678 -1142 ne
rect 5341 -1191 5393 -1185
rect 5678 -1191 5730 -1185
rect 5289 -1238 6086 -1232
rect 5289 -1272 5301 -1238
rect 5335 -1272 5382 -1238
rect 5416 -1272 5462 -1238
rect 5496 -1272 5542 -1238
rect 5576 -1272 5622 -1238
rect 5656 -1272 5702 -1238
rect 5736 -1272 5782 -1238
rect 5816 -1272 5862 -1238
rect 5896 -1272 5942 -1238
rect 5976 -1272 6086 -1238
rect 5289 -1275 6086 -1272
tri 6086 -1275 6129 -1232 sw
rect 5289 -1278 6471 -1275
tri 6050 -1311 6083 -1278 ne
rect 6083 -1281 6471 -1278
rect 6083 -1311 6419 -1281
rect 5238 -1317 5596 -1311
rect 5238 -1323 5249 -1317
rect 5301 -1323 5596 -1317
rect 5238 -1357 5244 -1323
rect 5301 -1357 5556 -1323
rect 5590 -1357 5596 -1323
rect 5238 -1369 5249 -1357
rect 5301 -1369 5596 -1357
rect 5238 -1387 5596 -1369
rect 5238 -1396 5249 -1387
rect 5301 -1396 5596 -1387
rect 5238 -1430 5244 -1396
rect 5301 -1430 5556 -1396
rect 5590 -1430 5596 -1396
rect 5238 -1439 5249 -1430
rect 5301 -1439 5596 -1430
rect 5238 -1458 5596 -1439
rect 5238 -1470 5249 -1458
rect 5301 -1470 5596 -1458
rect 5149 -1503 5201 -1497
rect 5238 -1504 5244 -1470
rect 5301 -1504 5556 -1470
rect 5590 -1504 5596 -1470
rect 5238 -1510 5249 -1504
rect 5301 -1510 5596 -1504
rect 5238 -1516 5596 -1510
rect 5678 -1317 6039 -1311
tri 6083 -1313 6085 -1311 ne
rect 6085 -1313 6419 -1311
rect 5730 -1323 6039 -1317
rect 5730 -1357 5999 -1323
rect 6033 -1357 6039 -1323
rect 5730 -1369 6039 -1357
rect 5678 -1387 6039 -1369
rect 5730 -1396 6039 -1387
rect 5730 -1430 5999 -1396
rect 6033 -1430 6039 -1396
rect 6419 -1345 6471 -1333
rect 6419 -1403 6471 -1397
rect 5730 -1439 6039 -1430
rect 5678 -1458 6039 -1439
rect 5730 -1470 6039 -1458
rect 5730 -1504 5999 -1470
rect 6033 -1504 6039 -1470
rect 5730 -1510 6039 -1504
rect 5678 -1516 6039 -1510
rect 5149 -1567 5201 -1555
rect 6255 -1545 6307 -1539
rect 5201 -1587 6255 -1575
rect 5201 -1619 5400 -1587
rect 5149 -1621 5400 -1619
rect 5434 -1597 6255 -1587
rect 5434 -1609 6307 -1597
rect 5434 -1621 6255 -1609
rect 5149 -1625 6255 -1621
rect 5394 -1659 5440 -1625
rect 5394 -1693 5400 -1659
rect 5434 -1693 5440 -1659
rect 5394 -1705 5440 -1693
rect 5837 -1673 5883 -1661
rect 6255 -1667 6307 -1661
rect 5837 -1707 5843 -1673
rect 5877 -1707 5883 -1673
rect 5837 -1742 5883 -1707
rect 5163 -1745 6223 -1742
rect 5163 -1748 5843 -1745
rect 5215 -1779 5843 -1748
rect 5877 -1748 6223 -1745
rect 5877 -1779 6171 -1748
rect 5215 -1792 6171 -1779
rect 5163 -1812 5215 -1800
rect 5163 -1870 5215 -1864
rect 6171 -1812 6223 -1800
rect 6171 -1870 6223 -1864
rect 6419 -1952 6471 -1946
rect 6419 -2016 6471 -2004
rect 5289 -2034 6419 -2028
rect 5289 -2068 5301 -2034
rect 5335 -2068 5400 -2034
rect 5434 -2068 5499 -2034
rect 5533 -2068 6419 -2034
rect 5289 -2074 6471 -2068
rect 5238 -2125 5596 -2119
rect 5238 -2131 5433 -2125
rect 5238 -2165 5244 -2131
rect 5278 -2165 5433 -2131
rect 5238 -2177 5433 -2165
rect 5485 -2131 5596 -2125
rect 5485 -2165 5556 -2131
rect 5590 -2165 5596 -2131
rect 5485 -2177 5596 -2165
rect 5238 -2195 5596 -2177
rect 5238 -2204 5433 -2195
rect 5238 -2238 5244 -2204
rect 5278 -2238 5433 -2204
rect 5238 -2247 5433 -2238
rect 5485 -2204 5596 -2195
rect 5485 -2238 5556 -2204
rect 5590 -2238 5596 -2204
rect 5485 -2247 5596 -2238
rect 5238 -2266 5596 -2247
rect 5238 -2278 5433 -2266
rect 5238 -2312 5244 -2278
rect 5278 -2312 5433 -2278
rect 5238 -2318 5433 -2312
rect 5485 -2278 5596 -2266
rect 5485 -2312 5556 -2278
rect 5590 -2312 5596 -2278
rect 5485 -2318 5596 -2312
rect 5238 -2324 5596 -2318
rect 6337 -2308 6389 -2302
rect 5163 -2360 6337 -2356
rect 5163 -2362 6389 -2360
rect 5215 -2368 6389 -2362
rect 5215 -2402 5400 -2368
rect 5434 -2372 6389 -2368
rect 5434 -2402 6337 -2372
rect 5215 -2406 6337 -2402
rect 5163 -2426 5215 -2414
rect 5163 -2484 5215 -2478
rect 5394 -2440 5440 -2406
rect 6337 -2430 6389 -2424
rect 5394 -2474 5400 -2440
rect 5434 -2474 5440 -2440
rect 5394 -2486 5440 -2474
<< via1 >>
rect 5281 10811 5286 10817
rect 5286 10811 5330 10817
rect 5330 10811 5333 10817
rect 5374 10811 5408 10817
rect 5408 10811 5426 10817
rect 5467 10811 5486 10817
rect 5486 10811 5519 10817
rect 5281 10773 5333 10811
rect 5374 10773 5426 10811
rect 5467 10773 5519 10811
rect 5281 10765 5286 10773
rect 5286 10765 5330 10773
rect 5330 10765 5333 10773
rect 5374 10765 5408 10773
rect 5408 10765 5426 10773
rect 5467 10765 5486 10773
rect 5486 10765 5519 10773
rect 5357 10571 5409 10585
rect 5357 10537 5366 10571
rect 5366 10537 5400 10571
rect 5400 10537 5409 10571
rect 5357 10533 5409 10537
rect 5357 10499 5409 10521
rect 5357 10469 5366 10499
rect 5366 10469 5400 10499
rect 5400 10469 5409 10499
rect 5279 10033 5331 10085
rect 5279 9969 5331 10021
rect 5279 9905 5331 9957
rect 5513 10571 5565 10585
rect 5513 10537 5522 10571
rect 5522 10537 5556 10571
rect 5556 10537 5565 10571
rect 5513 10533 5565 10537
rect 5513 10499 5565 10521
rect 5513 10469 5522 10499
rect 5522 10469 5556 10499
rect 5556 10469 5565 10499
rect 5435 10371 5487 10423
rect 5435 10307 5487 10359
rect 5435 10243 5487 10295
rect 5279 9709 5331 9761
rect 5279 9645 5331 9697
rect 5279 9581 5331 9633
rect 5591 10033 5643 10085
rect 5591 9969 5643 10021
rect 5591 9905 5643 9957
rect 5435 9371 5487 9423
rect 5435 9307 5487 9359
rect 5435 9243 5487 9295
rect 5279 8569 5331 8621
rect 5279 8505 5331 8557
rect 5279 8441 5331 8493
rect 5591 9709 5643 9761
rect 5591 9645 5643 9697
rect 5591 9581 5643 9633
rect 5435 8907 5487 8959
rect 5435 8843 5487 8895
rect 5435 8779 5487 8831
rect 5279 8245 5331 8297
rect 5279 8181 5331 8233
rect 5279 8117 5331 8169
rect 5591 8569 5643 8621
rect 5591 8505 5643 8557
rect 5591 8441 5643 8493
rect 5435 7907 5487 7959
rect 5435 7843 5487 7895
rect 5435 7779 5487 7831
rect 5279 7105 5331 7157
rect 5279 7041 5331 7093
rect 5279 6977 5331 7029
rect 5591 8245 5643 8297
rect 5591 8181 5643 8233
rect 5591 8117 5643 8169
rect 5435 7443 5487 7495
rect 5435 7379 5487 7431
rect 5435 7315 5487 7367
rect 5279 6781 5331 6833
rect 5279 6717 5331 6769
rect 5279 6653 5331 6705
rect 5591 7105 5643 7157
rect 5591 7041 5643 7093
rect 5591 6977 5643 7029
rect 5435 6443 5487 6495
rect 5435 6379 5487 6431
rect 5435 6315 5487 6367
rect 5591 6781 5643 6833
rect 5591 6717 5643 6769
rect 5591 6653 5643 6705
rect 5435 5979 5487 6031
rect 5435 5915 5487 5967
rect 5435 5851 5487 5903
rect 5279 5641 5331 5693
rect 5279 5577 5331 5629
rect 5279 5513 5331 5565
rect 5525 5641 5577 5693
rect 5525 5577 5577 5629
rect 5525 5513 5577 5565
rect 6211 3175 6263 3227
rect 6275 3175 6327 3227
rect 6211 3100 6263 3152
rect 6275 3100 6327 3152
rect 5928 2819 5980 2871
rect 5928 2744 5980 2796
rect 6020 2766 6072 2818
rect 6020 2691 6072 2743
rect 5249 2428 5301 2480
rect 5249 2353 5301 2405
rect 6112 2766 6164 2818
rect 6112 2691 6164 2743
rect 5341 2428 5393 2480
rect 5341 2353 5393 2405
rect 5433 2426 5485 2478
rect 5433 2351 5485 2403
rect 5525 2159 5577 2211
rect 5525 2095 5577 2147
rect 20811 2089 20863 2141
rect 20875 2089 20927 2141
rect 21338 2038 21454 2154
rect 25670 2084 25722 2136
rect 25670 2020 25722 2072
rect 25766 2084 25818 2136
rect 25766 2020 25818 2072
rect 25847 2123 25899 2175
rect 25847 2059 25899 2111
rect 25927 2149 25979 2201
rect 25927 2085 25979 2137
rect 25517 1818 25633 1934
rect 20811 1516 20863 1568
rect 20875 1516 20927 1568
rect 26009 1517 26061 1569
rect 26073 1517 26125 1569
rect 5624 1441 5676 1493
rect 5688 1441 5740 1493
rect 26185 1441 26237 1493
rect 26249 1441 26301 1493
rect 5709 1122 5761 1174
rect 25892 1136 25944 1188
rect 25956 1136 26008 1188
rect 5709 1058 5761 1110
rect 5807 1054 5859 1106
rect 5871 1054 5923 1106
rect 26062 1060 26114 1112
rect 26126 1060 26178 1112
rect 6252 265 6304 317
rect 6316 265 6368 317
rect 5525 232 5577 238
rect 5525 198 5535 232
rect 5535 198 5569 232
rect 5569 198 5577 232
rect 5525 186 5577 198
rect 5525 159 5577 168
rect 5525 125 5535 159
rect 5535 125 5569 159
rect 5569 125 5577 159
rect 5525 116 5577 125
rect 5525 85 5577 97
rect 5525 51 5535 85
rect 5535 51 5569 85
rect 5569 51 5577 85
rect 5525 45 5577 51
rect 5617 81 5669 133
rect 5149 -29 5201 23
rect 5149 -93 5201 -41
rect 5617 -22 5669 30
rect 5148 -216 5200 -164
rect 5148 -280 5200 -228
rect 5525 -529 5577 -523
rect 5525 -563 5556 -529
rect 5556 -563 5577 -529
rect 5525 -575 5577 -563
rect 5525 -602 5577 -593
rect 5525 -636 5556 -602
rect 5556 -636 5577 -602
rect 5525 -645 5577 -636
rect 5525 -676 5577 -664
rect 5148 -759 5200 -707
rect 5525 -710 5556 -676
rect 5556 -710 5577 -676
rect 5525 -716 5577 -710
rect 5801 -575 5853 -523
rect 5801 -645 5853 -593
rect 6419 -527 6471 -475
rect 6419 -591 6471 -539
rect 5801 -716 5853 -664
rect 5148 -823 5200 -771
rect 6009 -826 6061 -774
rect 6009 -890 6061 -838
rect 6575 -943 6627 -891
rect 5163 -1004 5215 -952
rect 6575 -1007 6627 -955
rect 5163 -1068 5215 -1016
rect 5341 -1118 5393 -1066
rect 5678 -1118 5730 -1066
rect 5341 -1185 5393 -1133
rect 5678 -1185 5730 -1133
rect 5249 -1323 5301 -1317
rect 5249 -1357 5278 -1323
rect 5278 -1357 5301 -1323
rect 5249 -1369 5301 -1357
rect 5249 -1396 5301 -1387
rect 5249 -1430 5278 -1396
rect 5278 -1430 5301 -1396
rect 5249 -1439 5301 -1430
rect 5249 -1470 5301 -1458
rect 5149 -1555 5201 -1503
rect 5249 -1504 5278 -1470
rect 5278 -1504 5301 -1470
rect 5249 -1510 5301 -1504
rect 5678 -1323 5730 -1317
rect 5678 -1357 5687 -1323
rect 5687 -1357 5721 -1323
rect 5721 -1357 5730 -1323
rect 5678 -1369 5730 -1357
rect 5678 -1396 5730 -1387
rect 5678 -1430 5687 -1396
rect 5687 -1430 5721 -1396
rect 5721 -1430 5730 -1396
rect 6419 -1333 6471 -1281
rect 6419 -1397 6471 -1345
rect 5678 -1439 5730 -1430
rect 5678 -1470 5730 -1458
rect 5678 -1504 5687 -1470
rect 5687 -1504 5721 -1470
rect 5721 -1504 5730 -1470
rect 5678 -1510 5730 -1504
rect 5149 -1619 5201 -1567
rect 6255 -1597 6307 -1545
rect 6255 -1661 6307 -1609
rect 5163 -1800 5215 -1748
rect 5163 -1864 5215 -1812
rect 6171 -1800 6223 -1748
rect 6171 -1864 6223 -1812
rect 6419 -2004 6471 -1952
rect 6419 -2068 6471 -2016
rect 5433 -2177 5485 -2125
rect 5433 -2247 5485 -2195
rect 5433 -2318 5485 -2266
rect 6337 -2360 6389 -2308
rect 5163 -2414 5215 -2362
rect 5163 -2478 5215 -2426
rect 6337 -2424 6389 -2372
<< metal2 >>
rect 5093 10818 5525 10847
rect 5093 10762 5102 10818
rect 5158 10762 5199 10818
rect 5255 10817 5525 10818
rect 5255 10765 5281 10817
rect 5333 10765 5374 10817
rect 5426 10765 5467 10817
rect 5519 10765 5525 10817
rect 5255 10762 5525 10765
rect 5093 10735 5525 10762
rect 5357 10585 6335 10591
rect 5409 10533 5513 10585
rect 5565 10533 6335 10585
rect 5357 10521 6335 10533
rect 5409 10469 5513 10521
rect 5565 10469 6335 10521
rect 5357 10463 6335 10469
tri 6162 10429 6196 10463 ne
rect 6196 10429 6335 10463
rect 5435 10423 5487 10429
tri 6196 10421 6204 10429 ne
rect 5435 10359 5487 10371
rect 5435 10295 5487 10307
tri 5404 10187 5435 10218 se
rect 5435 10187 5487 10243
rect 5176 10135 5487 10187
tri 5151 9423 5176 9448 se
rect 5176 9423 5228 10135
tri 5228 10104 5259 10135 nw
rect 5279 10085 6164 10091
rect 5331 10033 5591 10085
rect 5643 10033 6164 10085
rect 5279 10021 6164 10033
rect 5331 9969 5591 10021
rect 5643 9969 6164 10021
rect 5279 9957 6164 9969
rect 5331 9905 5591 9957
rect 5643 9905 6164 9957
rect 5279 9899 6164 9905
tri 6089 9876 6112 9899 ne
rect 5279 9761 6072 9767
rect 5331 9709 5591 9761
rect 5643 9709 6072 9761
rect 5279 9697 6072 9709
rect 5331 9645 5591 9697
rect 5643 9645 6072 9697
rect 5279 9633 6072 9645
rect 5331 9581 5591 9633
rect 5643 9581 6072 9633
rect 5279 9575 6072 9581
tri 5997 9552 6020 9575 ne
tri 5145 9417 5151 9423 se
rect 5151 9417 5228 9423
rect 4449 9365 5228 9417
rect 5435 9423 5487 9429
rect 4449 9359 4527 9365
tri 4527 9359 4533 9365 nw
rect 5435 9359 5487 9371
tri 4422 4025 4449 4052 se
rect 4449 4025 4501 9359
tri 4501 9333 4527 9359 nw
tri 5418 9333 5435 9350 se
tri 5405 9320 5418 9333 se
rect 5418 9320 5435 9333
rect 4295 4010 4501 4025
rect 4295 3973 4464 4010
tri 4464 3973 4501 4010 nw
rect 4539 9307 5435 9320
rect 4539 9295 5487 9307
rect 4539 9268 5435 9295
rect 4539 9243 4598 9268
tri 4598 9243 4623 9268 nw
tri 5404 9243 5429 9268 ne
rect 5429 9243 5435 9268
rect 4295 -2356 4347 3973
rect 4539 3935 4591 9243
tri 4591 9236 4598 9243 nw
tri 5429 9237 5435 9243 ne
rect 5435 9237 5487 9243
rect 5435 8959 5487 8965
tri 5404 8920 5435 8951 se
rect 4379 3883 4591 3935
rect 4623 8907 5435 8920
rect 4623 8895 5487 8907
rect 4623 8868 5435 8895
rect 4623 8843 4682 8868
tri 4682 8843 4707 8868 nw
tri 5405 8843 5430 8868 ne
rect 5430 8843 5435 8868
rect 4379 -1672 4431 3883
rect 4623 3826 4675 8843
tri 4675 8836 4682 8843 nw
tri 5430 8838 5435 8843 ne
rect 5435 8831 5487 8843
rect 5435 8773 5487 8779
rect 5279 8621 5980 8627
rect 5331 8569 5591 8621
rect 5643 8569 5980 8621
rect 5279 8557 5980 8569
rect 5331 8505 5591 8557
rect 5643 8505 5980 8557
rect 5279 8493 5980 8505
rect 5331 8441 5591 8493
rect 5643 8441 5980 8493
rect 5279 8435 5980 8441
tri 5905 8412 5928 8435 ne
rect 5279 8297 5853 8303
rect 5331 8245 5591 8297
rect 5643 8245 5853 8297
rect 5279 8233 5853 8245
rect 5331 8181 5591 8233
rect 5643 8181 5853 8233
rect 5279 8169 5853 8181
rect 5331 8117 5591 8169
rect 5643 8117 5853 8169
rect 5279 8111 5853 8117
tri 5758 8068 5801 8111 ne
rect 5435 7959 5487 7965
tri 5430 7895 5435 7900 se
rect 5435 7895 5487 7907
tri 5405 7870 5430 7895 se
rect 5430 7870 5435 7895
rect 4463 3774 4675 3826
rect 4711 7843 5435 7870
rect 4711 7831 5487 7843
rect 4711 7818 5435 7831
rect 4463 -1570 4515 3774
rect 4711 -946 4763 7818
tri 4763 7786 4795 7818 nw
tri 5404 7787 5435 7818 ne
rect 5435 7773 5487 7779
rect 5435 7495 5487 7501
tri 5404 7456 5435 7487 se
rect 4795 7443 5435 7456
rect 4795 7431 5487 7443
rect 4795 7404 5435 7431
rect 4795 7379 4854 7404
tri 4854 7379 4879 7404 nw
tri 5405 7379 5430 7404 ne
rect 5430 7379 5435 7404
rect 4795 -701 4847 7379
tri 4847 7372 4854 7379 nw
tri 5430 7374 5435 7379 ne
rect 5435 7367 5487 7379
rect 5435 7309 5487 7315
rect 5279 7157 5761 7163
rect 5331 7105 5591 7157
rect 5643 7105 5761 7157
rect 5279 7093 5761 7105
rect 5331 7041 5591 7093
rect 5643 7041 5761 7093
rect 5279 7029 5761 7041
rect 5331 6977 5591 7029
rect 5643 6977 5761 7029
rect 5279 6971 5761 6977
rect 5279 6833 5669 6839
rect 5331 6781 5591 6833
rect 5643 6781 5669 6833
rect 5279 6769 5669 6781
rect 5331 6717 5591 6769
rect 5643 6717 5669 6769
rect 5279 6705 5669 6717
rect 5331 6653 5591 6705
rect 5643 6653 5669 6705
rect 5279 6647 5669 6653
rect 5435 6495 5487 6501
tri 5430 6431 5435 6436 se
rect 5435 6431 5487 6443
tri 5405 6406 5430 6431 se
rect 5430 6406 5435 6431
rect 4885 6379 5435 6406
rect 4885 6367 5487 6379
rect 4885 6354 5435 6367
rect 4885 -158 4937 6354
tri 4937 6325 4966 6354 nw
tri 5404 6325 5433 6354 ne
rect 5433 6325 5435 6354
tri 5433 6323 5435 6325 ne
rect 5435 6309 5487 6315
rect 5435 6031 5487 6037
tri 5404 5992 5435 6023 se
rect 4969 5979 5435 5992
rect 4969 5967 5487 5979
rect 4969 5940 5435 5967
rect 4969 5915 5026 5940
tri 5026 5915 5051 5940 nw
tri 5405 5915 5430 5940 ne
rect 5430 5915 5435 5940
rect 4969 29 5021 5915
tri 5021 5910 5026 5915 nw
tri 5430 5910 5435 5915 ne
rect 5435 5903 5487 5915
rect 5435 5845 5487 5851
rect 5279 5693 5577 5699
rect 5331 5641 5525 5693
rect 5279 5629 5577 5641
rect 5331 5577 5525 5629
rect 5279 5565 5577 5577
rect 5331 5513 5525 5565
rect 5279 5507 5577 5513
rect 5249 2480 5301 2486
rect 5249 2405 5301 2428
rect 5249 955 5301 2353
rect 5341 2480 5393 2486
rect 5341 2405 5393 2428
tri 5301 955 5313 967 sw
rect 5249 923 5313 955
tri 5249 911 5261 923 ne
tri 5249 610 5261 622 se
rect 5261 610 5313 923
rect 5249 578 5313 610
rect 4969 23 5201 29
rect 4969 -23 5149 23
rect 5149 -41 5201 -29
rect 5149 -99 5201 -93
rect 4885 -164 5200 -158
rect 4885 -210 5148 -164
rect 5148 -228 5200 -216
rect 5148 -286 5200 -280
rect 4795 -707 5200 -701
rect 4795 -753 5148 -707
rect 5148 -771 5200 -759
rect 5148 -829 5200 -823
rect 4711 -952 5215 -946
rect 4711 -998 5163 -952
rect 5163 -1016 5215 -1004
rect 5163 -1074 5215 -1068
rect 5249 -1317 5301 578
tri 5301 566 5313 578 nw
rect 5249 -1387 5301 -1369
rect 5249 -1458 5301 -1439
rect 5149 -1503 5201 -1497
rect 5149 -1567 5201 -1555
rect 4463 -1619 5149 -1570
rect 4463 -1622 5201 -1619
rect 5149 -1625 5201 -1622
rect 4379 -1724 5215 -1672
rect 5163 -1748 5215 -1724
rect 5163 -1812 5215 -1800
rect 5163 -1870 5215 -1864
rect 4295 -2362 5215 -2356
rect 4295 -2408 5163 -2362
rect 5163 -2426 5215 -2414
rect 5163 -2484 5215 -2478
rect 5249 -2554 5301 -1510
rect 5341 -1066 5393 2353
rect 5341 -1133 5393 -1118
rect 5341 -2548 5393 -1185
rect 5433 2478 5485 2484
rect 5433 2403 5485 2426
rect 5433 -2125 5485 2351
rect 5525 2211 5577 5507
rect 5525 2147 5577 2159
rect 5525 238 5577 2095
rect 5525 168 5577 186
rect 5525 97 5577 116
rect 5525 39 5577 45
rect 5617 1493 5669 6647
rect 5709 1652 5761 6971
rect 5801 1709 5853 8111
rect 5928 2871 5980 8435
rect 5928 2796 5980 2819
rect 5928 2738 5980 2744
rect 6020 2818 6072 9575
rect 6020 2743 6072 2766
rect 6020 2685 6072 2691
rect 6112 2818 6164 9899
rect 6204 3227 6335 10429
rect 6204 3175 6211 3227
rect 6263 3175 6275 3227
rect 6327 3175 6335 3227
rect 6204 3152 6335 3175
rect 6204 3100 6211 3152
rect 6263 3100 6275 3152
rect 6327 3100 6335 3152
rect 6204 3094 6335 3100
rect 6112 2743 6164 2766
rect 6112 2685 6164 2691
rect 25927 2201 25979 2207
rect 25847 2175 25899 2181
rect 21338 2154 21454 2160
rect 20805 2089 20811 2141
rect 20863 2089 20875 2141
rect 20927 2089 20933 2141
tri 5853 1709 5870 1726 sw
tri 5801 1708 5802 1709 ne
rect 5802 1708 5870 1709
tri 5870 1708 5871 1709 sw
tri 5802 1669 5841 1708 ne
rect 5841 1669 5871 1708
tri 5761 1652 5778 1669 sw
tri 5841 1652 5858 1669 ne
rect 5858 1663 5871 1669
tri 5871 1663 5916 1708 sw
rect 5858 1652 5916 1663
tri 5709 1585 5776 1652 ne
rect 5776 1639 5778 1652
tri 5778 1639 5791 1652 sw
tri 5858 1639 5871 1652 ne
rect 5776 1609 5791 1639
tri 5791 1609 5821 1639 sw
rect 5617 1441 5624 1493
rect 5676 1441 5688 1493
rect 5740 1441 5746 1493
rect 5617 133 5669 1441
rect 5617 30 5669 81
rect 5617 -28 5669 -22
tri 5709 1334 5776 1401 se
rect 5776 1374 5821 1609
rect 5776 1361 5808 1374
tri 5808 1361 5821 1374 nw
rect 5776 1354 5801 1361
tri 5801 1354 5808 1361 nw
tri 5864 1354 5871 1361 se
rect 5871 1354 5916 1652
rect 20805 1568 20933 2089
rect 21338 1934 21454 2038
rect 25670 2136 25722 2142
rect 25670 2072 25722 2084
tri 21454 1934 21511 1991 sw
rect 21338 1865 25517 1934
tri 21338 1818 21385 1865 ne
rect 21385 1818 25517 1865
rect 25633 1818 25639 1934
rect 20805 1516 20811 1568
rect 20863 1516 20875 1568
rect 20927 1516 20933 1568
rect 5776 1334 5781 1354
tri 5781 1334 5801 1354 nw
tri 5844 1334 5864 1354 se
rect 5864 1334 5916 1354
rect 5709 1329 5776 1334
tri 5776 1329 5781 1334 nw
tri 5839 1329 5844 1334 se
rect 5844 1329 5873 1334
rect 5709 1174 5761 1329
tri 5761 1314 5776 1329 nw
tri 5824 1314 5839 1329 se
rect 5839 1314 5873 1329
rect 5709 1110 5761 1122
tri 5626 -270 5709 -187 se
rect 5709 -218 5761 1058
tri 5801 1291 5824 1314 se
rect 5824 1291 5873 1314
tri 5873 1291 5916 1334 nw
rect 5801 1289 5871 1291
tri 5871 1289 5873 1291 nw
rect 5801 1106 5853 1289
tri 5853 1271 5871 1289 nw
rect 25670 1136 25722 2020
rect 25766 2136 25818 2142
rect 25766 2072 25818 2084
rect 25766 1188 25818 2020
rect 25847 2111 25899 2123
rect 25847 1517 25899 2059
rect 25927 2137 25979 2149
rect 25927 1569 25979 2085
tri 25979 1569 26031 1621 sw
rect 25927 1541 26009 1569
tri 25927 1523 25945 1541 ne
rect 25945 1523 26009 1541
tri 25899 1517 25905 1523 sw
tri 25945 1517 25951 1523 ne
rect 25951 1517 26009 1523
rect 26061 1517 26073 1569
rect 26125 1517 26131 1569
rect 25847 1493 25905 1517
tri 25905 1493 25929 1517 sw
rect 25847 1489 25929 1493
tri 25929 1489 25933 1493 sw
tri 26175 1489 26179 1493 se
rect 26179 1489 26185 1493
rect 25847 1441 26185 1489
rect 26237 1441 26249 1493
rect 26301 1441 26307 1493
tri 25818 1188 25856 1226 sw
rect 25766 1166 25892 1188
tri 25766 1142 25790 1166 ne
rect 25790 1142 25892 1166
tri 25722 1136 25728 1142 sw
tri 25790 1136 25796 1142 ne
rect 25796 1136 25892 1142
rect 25944 1136 25956 1188
rect 26008 1136 26014 1188
rect 25670 1112 25728 1136
tri 25728 1112 25752 1136 sw
rect 25670 1108 25752 1112
tri 25752 1108 25756 1112 sw
tri 26052 1108 26056 1112 se
rect 26056 1108 26062 1112
rect 5801 1054 5807 1106
rect 5859 1054 5871 1106
rect 5923 1054 5929 1106
rect 25670 1060 26062 1108
rect 26114 1060 26126 1112
rect 26178 1060 26184 1112
tri 5790 427 5801 438 se
rect 5801 427 5853 1054
rect 5790 375 5853 427
rect 5790 102 5836 375
tri 5836 358 5853 375 nw
rect 6246 265 6252 317
rect 6304 265 6316 317
rect 6368 265 6374 317
tri 5836 102 5853 119 sw
rect 5790 50 5853 102
tri 5790 39 5801 50 ne
tri 5709 -270 5761 -218 nw
tri 5543 -353 5626 -270 se
tri 5626 -353 5709 -270 nw
tri 5525 -371 5543 -353 se
rect 5543 -371 5608 -353
tri 5608 -371 5626 -353 nw
rect 5525 -523 5577 -371
tri 5577 -402 5608 -371 nw
rect 5525 -593 5577 -575
rect 5525 -664 5577 -645
rect 5525 -722 5577 -716
rect 5801 -523 5853 50
rect 5801 -593 5853 -575
rect 6419 -475 6471 -469
rect 6419 -539 6471 -527
rect 6419 -597 6471 -591
rect 5801 -664 5853 -645
rect 5801 -722 5853 -716
rect 6009 -774 6061 -768
rect 6009 -838 6061 -826
rect 6009 -896 6061 -890
rect 6575 -891 6627 -885
rect 6575 -955 6627 -943
rect 6575 -1013 6627 -1007
rect 5678 -1066 5730 -1060
rect 5678 -1133 5730 -1118
rect 5678 -1317 5730 -1185
rect 5678 -1387 5730 -1369
rect 6419 -1281 6471 -1275
rect 6419 -1345 6471 -1333
rect 6419 -1403 6471 -1397
rect 5678 -1458 5730 -1439
rect 5678 -1516 5730 -1510
rect 6255 -1545 6307 -1539
rect 6255 -1609 6307 -1597
rect 6255 -1667 6307 -1661
rect 6171 -1748 6223 -1742
rect 6171 -1812 6223 -1800
rect 6171 -1870 6223 -1864
rect 6419 -1952 6471 -1946
rect 6419 -2016 6471 -2004
rect 6419 -2074 6471 -2068
rect 5433 -2195 5485 -2177
rect 5433 -2266 5485 -2247
rect 5433 -2524 5485 -2318
rect 6337 -2308 6389 -2302
rect 6337 -2372 6389 -2360
rect 6337 -2430 6389 -2424
tri 5433 -2534 5443 -2524 ne
rect 5443 -2534 5485 -2524
tri 5485 -2534 5508 -2511 sw
tri 5301 -2554 5307 -2548 sw
tri 5341 -2554 5347 -2548 ne
rect 5347 -2554 5393 -2548
rect 5249 -2564 5307 -2554
tri 5249 -2594 5279 -2564 ne
rect 5279 -2585 5307 -2564
tri 5307 -2585 5338 -2554 sw
tri 5347 -2585 5378 -2554 ne
rect 5378 -2574 5393 -2554
tri 5393 -2574 5433 -2534 sw
tri 5443 -2573 5482 -2534 ne
rect 5482 -2573 5508 -2534
tri 5508 -2573 5547 -2534 sw
tri 5482 -2574 5483 -2573 ne
rect 5483 -2574 5547 -2573
rect 5378 -2576 5433 -2574
tri 5433 -2576 5435 -2574 sw
tri 5483 -2576 5485 -2574 ne
rect 5485 -2576 5547 -2574
rect 5378 -2585 5435 -2576
tri 5435 -2585 5444 -2576 sw
tri 5485 -2585 5494 -2576 ne
rect 5494 -2585 5547 -2576
tri 5547 -2585 5559 -2573 sw
rect 5279 -2594 5338 -2585
tri 5338 -2594 5347 -2585 sw
tri 5378 -2594 5387 -2585 ne
rect 5387 -2594 5444 -2585
tri 5279 -2616 5301 -2594 ne
rect 5301 -2600 5347 -2594
tri 5347 -2600 5353 -2594 sw
tri 5387 -2600 5393 -2594 ne
rect 5393 -2600 5444 -2594
rect 5301 -2616 5353 -2600
tri 5301 -2662 5347 -2616 ne
rect 5347 -2622 5353 -2616
tri 5353 -2622 5375 -2600 sw
tri 5393 -2622 5415 -2600 ne
rect 5415 -2622 5444 -2600
rect 5347 -2651 5375 -2622
tri 5375 -2651 5404 -2622 sw
tri 5415 -2651 5444 -2622 ne
tri 5444 -2626 5485 -2585 sw
tri 5494 -2626 5535 -2585 ne
rect 5535 -2626 5559 -2585
rect 5444 -2638 5485 -2626
tri 5485 -2638 5497 -2626 sw
tri 5535 -2638 5547 -2626 ne
rect 5547 -2638 5559 -2626
tri 5559 -2638 5612 -2585 sw
rect 5444 -2651 5497 -2638
tri 5497 -2651 5510 -2638 sw
tri 5547 -2651 5560 -2638 ne
rect 5560 -2651 5612 -2638
tri 5612 -2651 5625 -2638 sw
rect 5347 -2662 5404 -2651
tri 5404 -2662 5415 -2651 sw
tri 5444 -2662 5455 -2651 ne
rect 5455 -2662 5510 -2651
tri 5347 -2730 5415 -2662 ne
tri 5415 -2690 5443 -2662 sw
tri 5455 -2690 5483 -2662 ne
rect 5483 -2688 5510 -2662
tri 5510 -2688 5547 -2651 sw
tri 5560 -2688 5597 -2651 ne
rect 5597 -2688 5625 -2651
rect 5483 -2690 5547 -2688
rect 5415 -2717 5443 -2690
tri 5443 -2717 5470 -2690 sw
tri 5483 -2717 5510 -2690 ne
rect 5510 -2703 5547 -2690
tri 5547 -2703 5562 -2688 sw
tri 5597 -2703 5612 -2688 ne
rect 5612 -2703 5625 -2688
tri 5625 -2703 5677 -2651 sw
rect 5510 -2717 5562 -2703
tri 5562 -2717 5576 -2703 sw
tri 5612 -2717 5626 -2703 ne
rect 5626 -2717 6166 -2703
tri 6166 -2717 6180 -2703 sw
rect 5415 -2730 5470 -2717
tri 5470 -2730 5483 -2717 sw
tri 5510 -2730 5523 -2717 ne
rect 5523 -2730 5576 -2717
tri 5415 -2798 5483 -2730 ne
tri 5483 -2758 5511 -2730 sw
tri 5523 -2758 5551 -2730 ne
rect 5551 -2753 5576 -2730
tri 5576 -2753 5612 -2717 sw
tri 5626 -2753 5662 -2717 ne
rect 5662 -2753 6180 -2717
rect 5551 -2758 5612 -2753
rect 5483 -2783 5511 -2758
tri 5511 -2783 5536 -2758 sw
tri 5551 -2783 5576 -2758 ne
rect 5576 -2783 5612 -2758
tri 5612 -2783 5642 -2753 sw
tri 6136 -2759 6142 -2753 ne
rect 6142 -2759 6180 -2753
tri 6180 -2759 6222 -2717 sw
tri 6142 -2783 6166 -2759 ne
rect 6166 -2783 6222 -2759
rect 5483 -2798 5536 -2783
tri 5536 -2798 5551 -2783 sw
tri 5576 -2798 5591 -2783 ne
rect 5591 -2798 6099 -2783
tri 5483 -2866 5551 -2798 ne
tri 5551 -2814 5567 -2798 sw
tri 5591 -2814 5607 -2798 ne
rect 5607 -2814 6099 -2798
tri 6099 -2814 6130 -2783 sw
tri 6166 -2787 6170 -2783 ne
rect 5551 -2825 5567 -2814
tri 5567 -2825 5578 -2814 sw
tri 5607 -2825 5618 -2814 ne
rect 5618 -2825 6130 -2814
rect 5551 -2847 5578 -2825
tri 5578 -2847 5600 -2825 sw
tri 6056 -2847 6078 -2825 ne
rect 5551 -2866 5600 -2847
tri 5600 -2866 5619 -2847 sw
tri 5551 -2880 5565 -2866 ne
rect 5565 -2880 6024 -2866
tri 6024 -2880 6038 -2866 sw
tri 5565 -2920 5605 -2880 ne
rect 5605 -2920 6038 -2880
tri 5971 -2935 5986 -2920 ne
tri 5918 -5278 5986 -5210 se
rect 5986 -5226 6038 -2920
tri 5986 -5278 6038 -5226 nw
tri 5850 -5346 5918 -5278 se
tri 5918 -5346 5986 -5278 nw
tri 5831 -5365 5850 -5346 se
rect 5850 -5365 5899 -5346
tri 5899 -5365 5918 -5346 nw
tri 5782 -5414 5831 -5365 se
rect 5831 -5414 5850 -5365
tri 5850 -5414 5899 -5365 nw
tri 6029 -5414 6078 -5365 se
rect 6078 -5383 6130 -2825
tri 5761 -5435 5782 -5414 se
rect 5782 -5435 5829 -5414
tri 5829 -5435 5850 -5414 nw
tri 6008 -5435 6029 -5414 se
rect 6029 -5435 6078 -5414
tri 6078 -5435 6130 -5383 nw
tri 5714 -5482 5761 -5435 se
rect 5761 -5482 5782 -5435
tri 5782 -5482 5829 -5435 nw
tri 6002 -5441 6008 -5435 se
rect 6008 -5441 6072 -5435
tri 6072 -5441 6078 -5435 nw
tri 5667 -5529 5714 -5482 se
rect 5714 -5529 5735 -5482
tri 5735 -5529 5782 -5482 nw
rect 6002 -5529 6054 -5441
tri 6054 -5459 6072 -5441 nw
rect 6170 -5511 6222 -2783
tri 5646 -5550 5667 -5529 se
rect 5667 -5550 5714 -5529
tri 5714 -5550 5735 -5529 nw
tri 5578 -5618 5646 -5550 se
tri 5646 -5618 5714 -5550 nw
tri 5515 -5681 5578 -5618 se
rect 5578 -5681 5583 -5618
tri 5583 -5681 5646 -5618 nw
rect 5515 -5902 5567 -5681
tri 5567 -5697 5583 -5681 nw
<< via2 >>
rect 5102 10762 5158 10818
rect 5199 10762 5255 10818
<< metal3 >>
rect 5097 17584 5260 17585
rect 5020 17578 5260 17584
rect 5020 17514 5021 17578
rect 5085 17514 5105 17578
rect 5169 17514 5189 17578
rect 5253 17514 5260 17578
rect 5020 17498 5260 17514
rect 5020 17434 5021 17498
rect 5085 17434 5105 17498
rect 5169 17434 5189 17498
rect 5253 17434 5260 17498
rect 5020 17418 5260 17434
rect 5020 17354 5021 17418
rect 5085 17354 5105 17418
rect 5169 17354 5189 17418
rect 5253 17354 5260 17418
rect 5020 17338 5260 17354
rect 5020 17274 5021 17338
rect 5085 17274 5105 17338
rect 5169 17274 5189 17338
rect 5253 17274 5260 17338
rect 5020 17258 5260 17274
rect 5020 17194 5021 17258
rect 5085 17194 5105 17258
rect 5169 17194 5189 17258
rect 5253 17194 5260 17258
rect 5020 17178 5260 17194
rect 5020 17114 5021 17178
rect 5085 17114 5105 17178
rect 5169 17114 5189 17178
rect 5253 17114 5260 17178
rect 5020 17098 5260 17114
rect 5020 17034 5021 17098
rect 5085 17034 5105 17098
rect 5169 17034 5189 17098
rect 5253 17034 5260 17098
rect 5020 17018 5260 17034
rect 5020 16954 5021 17018
rect 5085 16954 5105 17018
rect 5169 16954 5189 17018
rect 5253 16954 5260 17018
rect 5020 16938 5260 16954
rect 5020 16874 5021 16938
rect 5085 16874 5105 16938
rect 5169 16874 5189 16938
rect 5253 16874 5260 16938
rect 5020 16858 5260 16874
rect 5020 16794 5021 16858
rect 5085 16794 5105 16858
rect 5169 16794 5189 16858
rect 5253 16794 5260 16858
rect 5020 16778 5260 16794
rect 5020 16714 5021 16778
rect 5085 16714 5105 16778
rect 5169 16714 5189 16778
rect 5253 16714 5260 16778
rect 5020 16698 5260 16714
rect 5020 16634 5021 16698
rect 5085 16634 5105 16698
rect 5169 16634 5189 16698
rect 5253 16634 5260 16698
rect 5020 16618 5260 16634
rect 5020 16554 5021 16618
rect 5085 16554 5105 16618
rect 5169 16554 5189 16618
rect 5253 16554 5260 16618
rect 5020 16538 5260 16554
rect 5020 16474 5021 16538
rect 5085 16474 5105 16538
rect 5169 16474 5189 16538
rect 5253 16474 5260 16538
rect 5020 16458 5260 16474
rect 5020 16394 5021 16458
rect 5085 16394 5105 16458
rect 5169 16394 5189 16458
rect 5253 16394 5260 16458
rect 5020 16378 5260 16394
rect 5020 16314 5021 16378
rect 5085 16314 5105 16378
rect 5169 16314 5189 16378
rect 5253 16314 5260 16378
rect 5020 16298 5260 16314
rect 5020 16234 5021 16298
rect 5085 16234 5105 16298
rect 5169 16234 5189 16298
rect 5253 16234 5260 16298
rect 5020 16218 5260 16234
rect 5020 16154 5021 16218
rect 5085 16154 5105 16218
rect 5169 16154 5189 16218
rect 5253 16154 5260 16218
rect 5020 16138 5260 16154
rect 5020 16074 5021 16138
rect 5085 16074 5105 16138
rect 5169 16074 5189 16138
rect 5253 16074 5260 16138
rect 5020 16058 5260 16074
rect 5020 15994 5021 16058
rect 5085 15994 5105 16058
rect 5169 15994 5189 16058
rect 5253 15994 5260 16058
rect 5020 15977 5260 15994
rect 5020 15913 5021 15977
rect 5085 15913 5105 15977
rect 5169 15913 5189 15977
rect 5253 15913 5260 15977
rect 5020 15896 5260 15913
rect 5020 15832 5021 15896
rect 5085 15832 5105 15896
rect 5169 15832 5189 15896
rect 5253 15832 5260 15896
rect 5020 15815 5260 15832
rect 5020 15751 5021 15815
rect 5085 15751 5105 15815
rect 5169 15751 5189 15815
rect 5253 15751 5260 15815
rect 5020 15734 5260 15751
rect 5020 15670 5021 15734
rect 5085 15670 5105 15734
rect 5169 15670 5189 15734
rect 5253 15670 5260 15734
rect 5020 15653 5260 15670
rect 5020 15589 5021 15653
rect 5085 15589 5105 15653
rect 5169 15589 5189 15653
rect 5253 15589 5260 15653
rect 5020 15572 5260 15589
rect 5020 15508 5021 15572
rect 5085 15508 5105 15572
rect 5169 15508 5189 15572
rect 5253 15508 5260 15572
rect 5020 15491 5260 15508
rect 5020 15427 5021 15491
rect 5085 15427 5105 15491
rect 5169 15427 5189 15491
rect 5253 15427 5260 15491
rect 5020 15410 5260 15427
rect 5020 15346 5021 15410
rect 5085 15346 5105 15410
rect 5169 15346 5189 15410
rect 5253 15346 5260 15410
rect 5020 15329 5260 15346
rect 5020 15265 5021 15329
rect 5085 15265 5105 15329
rect 5169 15265 5189 15329
rect 5253 15265 5260 15329
rect 5020 15248 5260 15265
rect 5020 15184 5021 15248
rect 5085 15184 5105 15248
rect 5169 15184 5189 15248
rect 5253 15184 5260 15248
rect 5020 15178 5260 15184
tri 5020 15101 5097 15178 ne
rect 5097 10818 5260 15178
rect 5097 10762 5102 10818
rect 5158 10762 5199 10818
rect 5255 10762 5260 10818
rect 5097 10730 5260 10762
<< via3 >>
rect 5021 17514 5085 17578
rect 5105 17514 5169 17578
rect 5189 17514 5253 17578
rect 5021 17434 5085 17498
rect 5105 17434 5169 17498
rect 5189 17434 5253 17498
rect 5021 17354 5085 17418
rect 5105 17354 5169 17418
rect 5189 17354 5253 17418
rect 5021 17274 5085 17338
rect 5105 17274 5169 17338
rect 5189 17274 5253 17338
rect 5021 17194 5085 17258
rect 5105 17194 5169 17258
rect 5189 17194 5253 17258
rect 5021 17114 5085 17178
rect 5105 17114 5169 17178
rect 5189 17114 5253 17178
rect 5021 17034 5085 17098
rect 5105 17034 5169 17098
rect 5189 17034 5253 17098
rect 5021 16954 5085 17018
rect 5105 16954 5169 17018
rect 5189 16954 5253 17018
rect 5021 16874 5085 16938
rect 5105 16874 5169 16938
rect 5189 16874 5253 16938
rect 5021 16794 5085 16858
rect 5105 16794 5169 16858
rect 5189 16794 5253 16858
rect 5021 16714 5085 16778
rect 5105 16714 5169 16778
rect 5189 16714 5253 16778
rect 5021 16634 5085 16698
rect 5105 16634 5169 16698
rect 5189 16634 5253 16698
rect 5021 16554 5085 16618
rect 5105 16554 5169 16618
rect 5189 16554 5253 16618
rect 5021 16474 5085 16538
rect 5105 16474 5169 16538
rect 5189 16474 5253 16538
rect 5021 16394 5085 16458
rect 5105 16394 5169 16458
rect 5189 16394 5253 16458
rect 5021 16314 5085 16378
rect 5105 16314 5169 16378
rect 5189 16314 5253 16378
rect 5021 16234 5085 16298
rect 5105 16234 5169 16298
rect 5189 16234 5253 16298
rect 5021 16154 5085 16218
rect 5105 16154 5169 16218
rect 5189 16154 5253 16218
rect 5021 16074 5085 16138
rect 5105 16074 5169 16138
rect 5189 16074 5253 16138
rect 5021 15994 5085 16058
rect 5105 15994 5169 16058
rect 5189 15994 5253 16058
rect 5021 15913 5085 15977
rect 5105 15913 5169 15977
rect 5189 15913 5253 15977
rect 5021 15832 5085 15896
rect 5105 15832 5169 15896
rect 5189 15832 5253 15896
rect 5021 15751 5085 15815
rect 5105 15751 5169 15815
rect 5189 15751 5253 15815
rect 5021 15670 5085 15734
rect 5105 15670 5169 15734
rect 5189 15670 5253 15734
rect 5021 15589 5085 15653
rect 5105 15589 5169 15653
rect 5189 15589 5253 15653
rect 5021 15508 5085 15572
rect 5105 15508 5169 15572
rect 5189 15508 5253 15572
rect 5021 15427 5085 15491
rect 5105 15427 5169 15491
rect 5189 15427 5253 15491
rect 5021 15346 5085 15410
rect 5105 15346 5169 15410
rect 5189 15346 5253 15410
rect 5021 15265 5085 15329
rect 5105 15265 5169 15329
rect 5189 15265 5253 15329
rect 5021 15184 5085 15248
rect 5105 15184 5169 15248
rect 5189 15184 5253 15248
<< metal4 >>
rect 5019 17578 5255 17579
rect 5019 17514 5021 17578
rect 5085 17514 5105 17578
rect 5169 17514 5189 17578
rect 5253 17514 5255 17578
rect 5019 17498 5255 17514
rect 5019 17434 5021 17498
rect 5085 17434 5105 17498
rect 5169 17434 5189 17498
rect 5253 17434 5255 17498
rect 5019 17418 5255 17434
rect 5019 17354 5021 17418
rect 5085 17354 5105 17418
rect 5169 17354 5189 17418
rect 5253 17354 5255 17418
rect 5019 17338 5255 17354
rect 5019 17274 5021 17338
rect 5085 17274 5105 17338
rect 5169 17274 5189 17338
rect 5253 17274 5255 17338
rect 5019 17258 5255 17274
rect 5019 17194 5021 17258
rect 5085 17194 5105 17258
rect 5169 17194 5189 17258
rect 5253 17194 5255 17258
rect 5019 17178 5255 17194
rect 5019 17114 5021 17178
rect 5085 17114 5105 17178
rect 5169 17114 5189 17178
rect 5253 17114 5255 17178
rect 5019 17098 5255 17114
rect 5019 17034 5021 17098
rect 5085 17034 5105 17098
rect 5169 17034 5189 17098
rect 5253 17034 5255 17098
rect 5019 17018 5255 17034
rect 5019 16954 5021 17018
rect 5085 16954 5105 17018
rect 5169 16954 5189 17018
rect 5253 16954 5255 17018
rect 5019 16938 5255 16954
rect 5019 16874 5021 16938
rect 5085 16874 5105 16938
rect 5169 16874 5189 16938
rect 5253 16874 5255 16938
rect 5019 16858 5255 16874
rect 5019 16794 5021 16858
rect 5085 16794 5105 16858
rect 5169 16794 5189 16858
rect 5253 16794 5255 16858
rect 5019 16778 5255 16794
rect 5019 16714 5021 16778
rect 5085 16714 5105 16778
rect 5169 16714 5189 16778
rect 5253 16714 5255 16778
rect 5019 16698 5255 16714
rect 5019 16634 5021 16698
rect 5085 16634 5105 16698
rect 5169 16634 5189 16698
rect 5253 16634 5255 16698
rect 5019 16618 5255 16634
rect 5019 16554 5021 16618
rect 5085 16554 5105 16618
rect 5169 16554 5189 16618
rect 5253 16554 5255 16618
rect 5019 16538 5255 16554
rect 5019 16474 5021 16538
rect 5085 16474 5105 16538
rect 5169 16474 5189 16538
rect 5253 16474 5255 16538
rect 5019 16458 5255 16474
rect 5019 16394 5021 16458
rect 5085 16394 5105 16458
rect 5169 16394 5189 16458
rect 5253 16394 5255 16458
rect 5019 16378 5255 16394
rect 5019 16314 5021 16378
rect 5085 16314 5105 16378
rect 5169 16314 5189 16378
rect 5253 16314 5255 16378
rect 5019 16298 5255 16314
rect 5019 16234 5021 16298
rect 5085 16234 5105 16298
rect 5169 16234 5189 16298
rect 5253 16234 5255 16298
rect 5019 16218 5255 16234
rect 5019 16154 5021 16218
rect 5085 16154 5105 16218
rect 5169 16154 5189 16218
rect 5253 16154 5255 16218
rect 5019 16138 5255 16154
rect 5019 16074 5021 16138
rect 5085 16074 5105 16138
rect 5169 16074 5189 16138
rect 5253 16074 5255 16138
rect 5019 16058 5255 16074
rect 5019 15994 5021 16058
rect 5085 15994 5105 16058
rect 5169 15994 5189 16058
rect 5253 15994 5255 16058
rect 5019 15977 5255 15994
rect 5019 15913 5021 15977
rect 5085 15913 5105 15977
rect 5169 15913 5189 15977
rect 5253 15913 5255 15977
rect 5019 15896 5255 15913
rect 5019 15832 5021 15896
rect 5085 15832 5105 15896
rect 5169 15832 5189 15896
rect 5253 15832 5255 15896
rect 5019 15815 5255 15832
rect 5019 15751 5021 15815
rect 5085 15751 5105 15815
rect 5169 15751 5189 15815
rect 5253 15751 5255 15815
rect 5019 15734 5255 15751
rect 5019 15670 5021 15734
rect 5085 15670 5105 15734
rect 5169 15670 5189 15734
rect 5253 15670 5255 15734
rect 5019 15653 5255 15670
rect 5019 15589 5021 15653
rect 5085 15589 5105 15653
rect 5169 15589 5189 15653
rect 5253 15589 5255 15653
rect 5019 15572 5255 15589
rect 5019 15508 5021 15572
rect 5085 15508 5105 15572
rect 5169 15508 5189 15572
rect 5253 15508 5255 15572
rect 5019 15491 5255 15508
rect 5019 15427 5021 15491
rect 5085 15427 5105 15491
rect 5169 15427 5189 15491
rect 5253 15427 5255 15491
rect 5019 15410 5255 15427
rect 5019 15346 5021 15410
rect 5085 15346 5105 15410
rect 5169 15346 5189 15410
rect 5253 15346 5255 15410
rect 5019 15329 5255 15346
rect 5019 15265 5021 15329
rect 5085 15265 5105 15329
rect 5169 15265 5189 15329
rect 5253 15265 5255 15329
rect 5019 15248 5255 15265
rect 5019 15184 5021 15248
rect 5085 15184 5105 15248
rect 5169 15184 5189 15248
rect 5253 15184 5255 15248
rect 5019 15183 5255 15184
<< labels >>
flabel comment s 26592 1852 26592 1852 0 FreeSans 400 0 0 0 NGHS_H
flabel comment s 6187 -5344 6187 -5344 0 FreeSans 200 90 0 0 PGB_PAD_VDDIOQ_H_N
flabel comment s 6094 -5235 6094 -5235 0 FreeSans 200 90 0 0 PGA_PAD_VDDIOQ_H_N
flabel comment s 5336 -871 5336 -871 0 FreeSans 600 0 0 0 <2>
flabel comment s 5539 -5746 5539 -5746 0 FreeSans 400 90 0 0 PU_CSD_H
flabel comment s 5053 10274 5053 10274 0 FreeSans 400 270 0 0 CONDIODE
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 43391508
string GDS_START 43232354
<< end >>
