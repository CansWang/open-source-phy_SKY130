magic
tech sky130A
magscale 1 2
timestamp 1619862920
<< checkpaint >>
rect -1260 -1250 1344 1275
<< labels >>
flabel comment s 36 13 36 13 2 FreeSans 50 0 0 0 EM1O
flabel comment s 24 15 24 15 0 FreeSans 50 0 0 0 A
flabel comment s 60 15 60 15 0 FreeSans 50 0 0 0 B
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 9213680
string GDS_START 9212912
<< end >>
