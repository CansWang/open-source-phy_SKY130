// Level triggered programmable counter
// 
module moduleName (
    ports
);
    
endmodule