magic
tech sky130A
magscale 1 2
timestamp 1619862920
<< checkpaint >>
rect -1260 -1396 17264 41260
<< metal1 >>
tri 3115 39968 3147 40000 se
rect 2697 39916 2703 39968
rect 2755 39916 2793 39968
rect 2845 39916 2883 39968
rect 2935 39916 2973 39968
rect 3025 39916 3063 39968
rect 3115 39916 3158 39968
rect 2697 39876 3158 39916
rect 2697 39824 2703 39876
rect 2755 39824 2793 39876
rect 2845 39824 2883 39876
rect 2935 39824 2973 39876
rect 3025 39824 3063 39876
rect 3115 39824 3158 39876
rect 2697 39784 3158 39824
rect 2697 39732 2703 39784
rect 2755 39732 2793 39784
rect 2845 39732 2883 39784
rect 2935 39732 2973 39784
rect 3025 39732 3063 39784
rect 3115 39732 3158 39784
rect 3342 39782 3799 39961
rect 15429 39770 15848 39986
tri 3115 39700 3147 39732 ne
rect 954 38664 960 38716
rect 1012 38664 1024 38716
rect 1076 38664 2546 38716
tri 2460 38630 2494 38664 ne
rect 1014 38387 1020 38439
rect 1072 38387 1084 38439
rect 1136 38387 2466 38439
tri 2380 38353 2414 38387 ne
rect 2414 38204 2466 38387
rect 2494 38322 2546 38664
rect 3449 38545 3455 38597
rect 3507 38545 3519 38597
rect 3571 38545 3577 38597
tri 2546 38322 2580 38356 sw
rect 2494 38270 3455 38322
rect 3507 38270 3519 38322
rect 3571 38270 3577 38322
tri 2466 38204 2500 38238 sw
rect 2414 38152 3210 38204
rect 3262 38152 3274 38204
rect 3326 38152 3332 38204
rect 2470 38107 3333 38113
rect 2522 38061 3333 38107
rect 2470 38043 2522 38055
tri 2522 38027 2556 38061 nw
rect 15862 38051 15914 38057
tri 15846 38027 15862 38043 se
tri 15828 38009 15846 38027 se
rect 15846 38009 15862 38027
rect 2470 37985 2522 37991
rect 2774 37907 2780 37959
rect 2832 37907 2844 37959
rect 2896 37958 2902 37959
tri 2902 37958 2903 37959 sw
rect 2896 37907 8463 37958
rect 13588 37929 13594 37981
rect 13646 37929 13660 37981
rect 13712 37929 13718 37981
rect 15473 37934 15595 38006
rect 15818 37999 15862 38009
rect 15818 37987 15914 37999
rect 15818 37935 15862 37987
rect 15818 37929 15914 37935
rect 2774 37906 8463 37907
rect 2774 37897 8521 37906
tri 8521 37897 8530 37906 nw
rect 2774 37894 8463 37897
rect 2774 37891 8341 37894
rect 2774 37839 2780 37891
rect 2832 37839 2844 37891
rect 2896 37842 8341 37891
rect 8393 37842 8405 37894
rect 8457 37842 8463 37894
rect 2896 37839 8463 37842
tri 8463 37839 8521 37897 nw
rect 2550 37664 2556 37716
rect 2608 37664 2620 37716
rect 2672 37664 4271 37716
rect 4323 37664 4335 37716
rect 4387 37664 4395 37716
rect 2390 37407 2442 37413
rect 3301 37377 3307 37429
rect 3359 37377 3371 37429
rect 3423 37377 3429 37429
rect 2390 37343 2442 37355
tri 2442 37337 2476 37371 sw
rect 2442 37291 3333 37337
rect 2390 37285 3333 37291
tri 15426 37210 15460 37244 ne
rect 2435 37101 2902 37124
rect 2435 37049 2780 37101
rect 2832 37049 2844 37101
rect 2896 37049 2902 37101
rect 2435 37028 2902 37049
rect 13866 37101 13918 37107
rect 15723 37101 15775 37107
rect 13866 37037 13918 37049
rect 2435 36998 2521 37028
tri 2521 36998 2551 37028 nw
rect 1284 36946 2058 36998
rect 2162 36482 2259 36998
rect 2131 36459 2137 36482
tri 2024 36354 2129 36459 ne
rect 2129 36430 2137 36459
rect 2189 36430 2201 36482
rect 2253 36430 2259 36482
rect 2129 36406 2259 36430
rect 2129 36354 2137 36406
rect 2189 36354 2201 36406
rect 2253 36354 2259 36406
tri 2401 36222 2435 36256 se
rect 2435 36222 2517 36998
tri 2517 36994 2521 36998 nw
tri 13918 37031 13952 37065 sw
tri 15689 37031 15723 37065 se
rect 15723 37037 15775 37049
rect 13918 36985 15723 37031
rect 13866 36979 15775 36985
rect 794 36203 2517 36222
rect 794 36151 800 36203
rect 852 36151 864 36203
rect 916 36151 2517 36203
rect 2612 36202 3014 36319
rect 794 36140 2517 36151
rect 0 36079 3141 36080
rect 0 36074 397 36079
rect 0 36022 157 36074
rect 209 36022 269 36074
rect 321 36027 397 36074
rect 449 36027 489 36079
rect 541 36027 581 36079
rect 633 36027 673 36079
rect 725 36074 3141 36079
rect 725 36027 2131 36074
rect 321 36022 2131 36027
rect 2183 36022 2207 36074
rect 2259 36022 3141 36074
rect 0 35997 3141 36022
rect 0 35996 397 35997
rect 0 35944 157 35996
rect 209 35944 269 35996
rect 321 35945 397 35996
rect 449 35945 489 35997
rect 541 35945 581 35997
rect 633 35945 673 35997
rect 725 35996 3141 35997
rect 725 35945 2131 35996
rect 321 35944 2131 35945
rect 2183 35944 2207 35996
rect 2259 35944 3141 35996
rect 0 35917 3141 35944
rect 0 35865 157 35917
rect 209 35865 269 35917
rect 321 35915 2131 35917
rect 321 35865 397 35915
rect 0 35863 397 35865
rect 449 35863 489 35915
rect 541 35863 581 35915
rect 633 35863 673 35915
rect 725 35865 2131 35915
rect 2183 35865 2207 35917
rect 2259 35865 3141 35917
rect 725 35863 3141 35865
rect 0 35838 3141 35863
rect 0 35786 157 35838
rect 209 35786 269 35838
rect 321 35833 2131 35838
rect 321 35786 397 35833
rect 0 35781 397 35786
rect 449 35781 489 35833
rect 541 35781 581 35833
rect 633 35781 673 35833
rect 725 35786 2131 35833
rect 2183 35786 2207 35838
rect 2259 35786 3141 35838
rect 725 35781 3141 35786
rect 0 35780 3141 35781
tri 2058 35701 2064 35707 se
rect 2064 35655 2070 35707
rect 2122 35655 2149 35707
rect 2201 35655 2227 35707
rect 2279 35655 2305 35707
rect 2357 35655 2363 35707
tri 2363 35701 2369 35707 sw
tri 5489 3800 5496 3807 se
rect 5496 3800 8566 3807
tri 8566 3800 8573 3807 sw
rect 1090 3770 1142 3776
tri 1142 3731 1185 3774 sw
tri 1844 3731 1878 3765 se
rect 1878 3760 2175 3800
tri 5453 3764 5489 3800 se
rect 5489 3767 8573 3800
rect 5489 3764 5498 3767
rect 1878 3731 1923 3760
tri 1923 3731 1952 3760 nw
tri 2101 3751 2110 3760 ne
rect 2110 3751 2175 3760
tri 2175 3751 2188 3764 sw
tri 5440 3751 5453 3764 se
rect 5453 3751 5498 3764
tri 5498 3751 5514 3767 nw
tri 8548 3751 8564 3767 ne
rect 8564 3764 8573 3767
tri 8573 3764 8609 3800 sw
rect 8564 3751 8609 3764
tri 8609 3751 8622 3764 sw
tri 2110 3731 2130 3751 ne
rect 2130 3731 2188 3751
rect 1142 3718 1918 3731
tri 1918 3726 1923 3731 nw
tri 2130 3726 2135 3731 ne
rect 2135 3730 2188 3731
tri 2188 3730 2209 3751 sw
tri 5438 3749 5440 3751 se
rect 5440 3749 5496 3751
tri 5496 3749 5498 3751 nw
tri 8564 3749 8566 3751 ne
rect 8566 3749 8764 3751
tri 5419 3730 5438 3749 se
rect 5438 3730 5477 3749
tri 5477 3730 5496 3749 nw
tri 8566 3730 8585 3749 ne
rect 8585 3730 8764 3749
rect 1090 3706 1918 3718
rect 1142 3691 1918 3706
rect 2135 3699 5446 3730
tri 5446 3699 5477 3730 nw
tri 8585 3699 8616 3730 ne
rect 8616 3699 8764 3730
rect 8816 3699 8828 3751
rect 8880 3699 8886 3751
rect 1090 3648 1142 3654
tri 1142 3648 1185 3691 nw
rect 2135 3690 5437 3699
tri 5437 3690 5446 3699 nw
rect 1134 3460 1140 3512
rect 1192 3460 1204 3512
rect 1256 3509 1262 3512
tri 1262 3509 1265 3512 sw
tri 9503 3509 9505 3511 se
rect 9505 3509 9511 3511
rect 1256 3469 9511 3509
rect 1256 3464 1266 3469
tri 1266 3464 1271 3469 nw
tri 9500 3464 9505 3469 ne
rect 1256 3460 1262 3464
tri 1262 3460 1266 3464 nw
rect 9505 3459 9511 3469
rect 9563 3459 9575 3511
rect 9627 3459 9633 3511
tri 1340 3432 1344 3436 se
rect 1344 3432 9298 3436
rect 1073 3380 1079 3432
rect 1131 3380 1143 3432
rect 1195 3431 9298 3432
tri 9298 3431 9303 3436 sw
rect 1195 3396 9434 3431
rect 1195 3392 1384 3396
tri 1384 3392 1388 3396 nw
tri 9253 3392 9257 3396 ne
rect 9257 3392 9434 3396
rect 1195 3380 1201 3392
tri 1201 3380 1213 3392 nw
tri 9257 3391 9258 3392 ne
rect 9258 3391 9434 3392
tri 9421 3384 9428 3391 ne
rect 9428 3379 9434 3391
rect 9486 3379 9498 3431
rect 9550 3379 9556 3431
rect 9334 910 9654 1086
rect 9602 789 9654 795
rect 9143 710 9195 737
rect 9330 687 9363 788
rect 9602 725 9654 737
rect 9786 678 9818 789
rect 9602 667 9654 673
rect 9143 646 9195 658
rect 10320 642 10351 759
rect 11416 728 11524 760
rect 11816 725 11876 762
rect 12069 729 12160 763
rect 9143 588 9195 594
rect 10972 361 11001 477
rect 9008 285 9360 337
rect 9412 285 9445 337
rect 9497 285 9503 337
rect 10366 69 10823 248
<< via1 >>
rect 2703 39916 2755 39968
rect 2793 39916 2845 39968
rect 2883 39916 2935 39968
rect 2973 39916 3025 39968
rect 3063 39916 3115 39968
rect 2703 39824 2755 39876
rect 2793 39824 2845 39876
rect 2883 39824 2935 39876
rect 2973 39824 3025 39876
rect 3063 39824 3115 39876
rect 2703 39732 2755 39784
rect 2793 39732 2845 39784
rect 2883 39732 2935 39784
rect 2973 39732 3025 39784
rect 3063 39732 3115 39784
rect 960 38664 1012 38716
rect 1024 38664 1076 38716
rect 1020 38387 1072 38439
rect 1084 38387 1136 38439
rect 3455 38545 3507 38597
rect 3519 38545 3571 38597
rect 3455 38270 3507 38322
rect 3519 38270 3571 38322
rect 3210 38152 3262 38204
rect 3274 38152 3326 38204
rect 2470 38055 2522 38107
rect 2470 37991 2522 38043
rect 2780 37907 2832 37959
rect 2844 37907 2896 37959
rect 13594 37929 13646 37981
rect 13660 37929 13712 37981
rect 15862 37999 15914 38051
rect 15862 37935 15914 37987
rect 2780 37839 2832 37891
rect 2844 37839 2896 37891
rect 8341 37842 8393 37894
rect 8405 37842 8457 37894
rect 2556 37664 2608 37716
rect 2620 37664 2672 37716
rect 4271 37664 4323 37716
rect 4335 37664 4387 37716
rect 2390 37355 2442 37407
rect 3307 37377 3359 37429
rect 3371 37377 3423 37429
rect 2390 37291 2442 37343
rect 2780 37049 2832 37101
rect 2844 37049 2896 37101
rect 13866 37049 13918 37101
rect 2137 36430 2189 36482
rect 2201 36430 2253 36482
rect 2137 36354 2189 36406
rect 2201 36354 2253 36406
rect 13866 36985 13918 37037
rect 15723 37049 15775 37101
rect 15723 36985 15775 37037
rect 800 36151 852 36203
rect 864 36151 916 36203
rect 157 36022 209 36074
rect 269 36022 321 36074
rect 397 36027 449 36079
rect 489 36027 541 36079
rect 581 36027 633 36079
rect 673 36027 725 36079
rect 2131 36022 2183 36074
rect 2207 36022 2259 36074
rect 157 35944 209 35996
rect 269 35944 321 35996
rect 397 35945 449 35997
rect 489 35945 541 35997
rect 581 35945 633 35997
rect 673 35945 725 35997
rect 2131 35944 2183 35996
rect 2207 35944 2259 35996
rect 157 35865 209 35917
rect 269 35865 321 35917
rect 397 35863 449 35915
rect 489 35863 541 35915
rect 581 35863 633 35915
rect 673 35863 725 35915
rect 2131 35865 2183 35917
rect 2207 35865 2259 35917
rect 157 35786 209 35838
rect 269 35786 321 35838
rect 397 35781 449 35833
rect 489 35781 541 35833
rect 581 35781 633 35833
rect 673 35781 725 35833
rect 2131 35786 2183 35838
rect 2207 35786 2259 35838
rect 2070 35655 2122 35707
rect 2149 35655 2201 35707
rect 2227 35655 2279 35707
rect 2305 35655 2357 35707
rect 1090 3718 1142 3770
rect 1090 3654 1142 3706
rect 8764 3699 8816 3751
rect 8828 3699 8880 3751
rect 1140 3460 1192 3512
rect 1204 3460 1256 3512
rect 9511 3459 9563 3511
rect 9575 3459 9627 3511
rect 1079 3380 1131 3432
rect 1143 3380 1195 3432
rect 9434 3379 9486 3431
rect 9498 3379 9550 3431
rect 9143 658 9195 710
rect 9602 737 9654 789
rect 9602 673 9654 725
rect 9143 594 9195 646
rect 9360 285 9412 337
rect 9445 285 9497 337
<< metal2 >>
rect 1351 39916 2703 39968
rect 2755 39916 2793 39968
rect 2845 39916 2883 39968
rect 2935 39916 2973 39968
rect 3025 39916 3063 39968
rect 3115 39916 3121 39968
rect 1351 39876 3121 39916
rect 1351 39824 2703 39876
rect 2755 39824 2793 39876
rect 2845 39824 2883 39876
rect 2935 39824 2973 39876
rect 3025 39824 3063 39876
rect 3115 39824 3121 39876
rect 1351 39784 3121 39824
rect 1351 39732 2703 39784
rect 2755 39732 2793 39784
rect 2845 39732 2883 39784
rect 2935 39732 2973 39784
rect 3025 39732 3063 39784
rect 3115 39732 3121 39784
tri 1752 39524 1960 39732 nw
rect 954 38664 960 38716
rect 1012 38664 1024 38716
rect 1076 38664 1082 38716
rect 8392 38683 8418 38696
tri 225 37101 359 37235 se
rect 359 37101 457 37152
tri 457 37101 508 37152 nw
tri 204 37080 225 37101 se
rect 225 37080 436 37101
tri 436 37080 457 37101 nw
tri 173 37049 204 37080 se
rect 204 37049 405 37080
tri 405 37049 436 37080 nw
tri 549 37049 580 37080 se
rect 580 37049 921 37050
tri 161 37037 173 37049 se
rect 173 37037 393 37049
tri 393 37037 405 37049 nw
tri 537 37037 549 37049 se
rect 549 37037 921 37049
tri 157 37033 161 37037 se
rect 161 37033 389 37037
tri 389 37033 393 37037 nw
tri 533 37033 537 37037 se
rect 537 37033 921 37037
rect 157 36985 341 37033
tri 341 36985 389 37033 nw
tri 485 36985 533 37033 se
rect 533 36985 921 37033
rect 157 36074 321 36985
tri 321 36965 341 36985 nw
tri 465 36965 485 36985 se
rect 485 36965 921 36985
rect 209 36022 269 36074
rect 157 35996 321 36022
rect 209 35944 269 35996
rect 157 35917 321 35944
rect 209 35865 269 35917
rect 157 35838 321 35865
rect 209 35786 269 35838
rect 157 35780 321 35786
tri 391 36891 465 36965 se
rect 465 36891 921 36965
rect 391 36528 921 36891
rect 391 36482 875 36528
tri 875 36482 921 36528 nw
rect 391 36430 823 36482
tri 823 36430 875 36482 nw
rect 391 36406 799 36430
tri 799 36406 823 36430 nw
rect 391 36354 747 36406
tri 747 36354 799 36406 nw
rect 391 36079 731 36354
tri 731 36338 747 36354 nw
rect 794 36151 800 36203
rect 852 36151 864 36203
rect 916 36151 922 36203
tri 794 36123 822 36151 ne
rect 391 36027 397 36079
rect 449 36027 489 36079
rect 541 36027 581 36079
rect 633 36027 673 36079
rect 725 36027 731 36079
rect 391 35997 731 36027
rect 391 35945 397 35997
rect 449 35945 489 35997
rect 541 35945 581 35997
rect 633 35945 673 35997
rect 725 35945 731 35997
rect 391 35915 731 35945
rect 391 35863 397 35915
rect 449 35863 489 35915
rect 541 35863 581 35915
rect 633 35863 673 35915
rect 725 35863 731 35915
rect 391 35833 731 35863
rect 391 35781 397 35833
rect 449 35781 489 35833
rect 541 35781 581 35833
rect 633 35781 673 35833
rect 725 35781 731 35833
rect 391 35780 731 35781
rect 822 35669 922 36151
rect 954 7453 986 38664
tri 986 38630 1020 38664 nw
rect 1014 38387 1020 38439
rect 1072 38387 1084 38439
rect 1136 38387 1142 38439
rect 1014 7499 1046 38387
tri 1046 38353 1080 38387 nw
rect 3204 38204 3332 38639
rect 3449 38545 3455 38597
rect 3507 38545 3519 38597
rect 3571 38545 3577 38597
rect 3449 38322 3577 38545
rect 3449 38270 3455 38322
rect 3507 38270 3519 38322
rect 3571 38270 3577 38322
rect 3204 38152 3210 38204
rect 3262 38152 3274 38204
rect 3326 38152 3332 38204
rect 2470 38107 2522 38113
rect 2470 38043 2522 38055
rect 2390 37407 2442 37413
rect 2390 37343 2442 37355
tri 2356 36879 2390 36913 se
rect 2390 36831 2442 37291
tri 2454 36793 2470 36809 se
rect 2470 36793 2522 37991
rect 15848 38051 15914 38057
rect 15848 38048 15862 38051
rect 15848 37992 15853 38048
rect 15909 37992 15914 37999
rect 15848 37987 15914 37992
rect 2774 37907 2780 37959
rect 2832 37907 2844 37959
rect 2896 37907 2902 37959
rect 13588 37929 13594 37981
rect 13646 37929 13660 37981
rect 13712 37929 13718 37981
tri 13632 37916 13645 37929 ne
rect 13645 37916 13718 37929
rect 2774 37891 2902 37907
rect 2774 37839 2780 37891
rect 2832 37839 2844 37891
rect 2896 37839 2902 37891
rect 8335 37894 8463 37916
tri 13645 37895 13666 37916 ne
rect 8335 37842 8341 37894
rect 8393 37842 8405 37894
rect 8457 37842 8463 37894
rect 8335 37839 8463 37842
tri 2017 36779 2031 36793 se
tri 2440 36779 2454 36793 se
rect 2454 36779 2522 36793
rect 1621 36711 2048 36779
tri 2436 36775 2440 36779 se
rect 2440 36775 2522 36779
rect 2470 36728 2522 36775
rect 2550 37664 2556 37716
rect 2608 37664 2620 37716
rect 2672 37664 2678 37716
tri 1587 36207 1621 36241 se
rect 1621 36207 1653 36711
tri 1653 36677 1687 36711 nw
tri 1997 36677 2031 36711 ne
tri 2516 36623 2550 36657 se
rect 2550 36575 2602 37664
tri 2602 37630 2636 37664 nw
rect 2774 37101 2902 37839
rect 4265 37664 4271 37716
rect 4323 37664 4335 37716
rect 4387 37664 4393 37716
rect 3301 37377 3307 37429
rect 3359 37377 3371 37429
rect 3423 37377 3429 37429
tri 3363 37343 3397 37377 ne
rect 2774 37049 2780 37101
rect 2832 37049 2844 37101
rect 2896 37049 2902 37101
rect 2774 37028 2902 37049
tri 3395 36575 3397 36577 se
rect 3397 36575 3429 37377
rect 13666 37317 13718 37916
rect 15848 37968 15862 37987
rect 15848 37912 15853 37968
rect 15909 37912 15914 37935
rect 15848 37903 15914 37912
tri 13666 37287 13696 37317 ne
rect 13696 37287 13718 37317
tri 13718 37287 13770 37339 sw
tri 13696 37265 13718 37287 ne
rect 13718 37265 13770 37287
tri 13718 37213 13770 37265 ne
tri 13770 37213 13844 37287 sw
rect 15184 37213 15187 37244
tri 15187 37213 15218 37244 nw
tri 13770 37139 13844 37213 ne
tri 13844 37139 13918 37213 sw
tri 15184 37210 15187 37213 nw
tri 13844 37117 13866 37139 ne
rect 13866 37101 13918 37139
rect 13866 37037 13918 37049
rect 13866 36979 13918 36985
rect 15721 37101 15777 37107
rect 15721 37091 15723 37101
rect 15775 37091 15777 37101
rect 15721 37011 15723 37035
rect 15775 37011 15777 37035
rect 15721 36946 15777 36955
tri 15184 36845 15218 36879 sw
tri 3363 36543 3395 36575 se
rect 3395 36543 3429 36575
tri 2017 36497 2063 36543 se
rect 2063 36511 3429 36543
tri 2063 36497 2077 36511 nw
tri 2002 36482 2017 36497 se
rect 2017 36482 2048 36497
tri 2048 36482 2063 36497 nw
tri 1971 36451 2002 36482 se
rect 2002 36451 2017 36482
tri 2017 36451 2048 36482 nw
tri 1950 36430 1971 36451 se
rect 1971 36430 1996 36451
tri 1996 36430 2017 36451 nw
rect 2131 36430 2137 36482
rect 2189 36430 2201 36482
rect 2253 36430 2259 36482
tri 1926 36406 1950 36430 se
rect 1950 36406 1972 36430
tri 1972 36406 1996 36430 nw
rect 2131 36406 2259 36430
tri 1925 36405 1926 36406 se
rect 1926 36405 1971 36406
tri 1971 36405 1972 36406 nw
tri 1879 36359 1925 36405 se
tri 1925 36359 1971 36405 nw
tri 1874 36354 1879 36359 se
rect 1879 36354 1920 36359
tri 1920 36354 1925 36359 nw
rect 2131 36354 2137 36406
rect 2189 36354 2201 36406
rect 2253 36354 2259 36406
tri 1833 36313 1874 36354 se
rect 1874 36313 1879 36354
tri 1879 36313 1920 36354 nw
tri 1787 36267 1833 36313 se
tri 1833 36267 1879 36313 nw
tri 1741 36221 1787 36267 se
tri 1787 36221 1833 36267 nw
rect 1074 36175 1653 36207
tri 1695 36175 1741 36221 se
tri 1741 36175 1787 36221 nw
rect 1074 7537 1104 36175
tri 1104 36141 1138 36175 nw
tri 1661 36141 1695 36175 se
rect 1695 36141 1707 36175
tri 1707 36141 1741 36175 nw
tri 1142 36095 1188 36141 se
rect 1188 36109 1675 36141
tri 1675 36109 1707 36141 nw
tri 1188 36095 1202 36109 nw
tri 1133 36086 1142 36095 se
rect 1142 36086 1179 36095
tri 1179 36086 1188 36095 nw
rect 1133 36074 1167 36086
tri 1167 36074 1179 36086 nw
rect 2131 36074 2259 36354
rect 1133 7603 1165 36074
tri 1165 36072 1167 36074 nw
rect 2183 36022 2207 36074
rect 2131 35996 2259 36022
rect 2183 35944 2207 35996
rect 2131 35917 2259 35944
rect 2183 35865 2207 35917
rect 2131 35838 2259 35865
rect 2183 35786 2207 35838
rect 2131 35780 2259 35786
rect 2064 35655 2070 35707
rect 2122 35655 2149 35707
rect 2201 35655 2227 35707
rect 2279 35655 2305 35707
rect 2357 35655 2363 35707
tri 1165 7603 1179 7617 sw
tri 1133 7557 1179 7603 ne
tri 1179 7557 1225 7603 sw
tri 1179 7549 1187 7557 ne
rect 1187 7549 1225 7557
tri 1104 7537 1116 7549 sw
tri 1187 7537 1199 7549 ne
rect 1199 7537 1225 7549
tri 1074 7503 1108 7537 ne
rect 1108 7503 1116 7537
tri 1046 7499 1050 7503 sw
tri 1108 7499 1112 7503 ne
rect 1112 7499 1116 7503
rect 1014 7495 1050 7499
tri 1050 7495 1054 7499 sw
tri 1112 7495 1116 7499 ne
tri 1116 7495 1158 7537 sw
tri 1199 7511 1225 7537 ne
tri 1225 7520 1262 7557 sw
rect 1225 7511 1262 7520
tri 1225 7506 1230 7511 ne
rect 1014 7489 1054 7495
tri 1014 7459 1044 7489 ne
rect 1044 7459 1054 7489
tri 1054 7459 1090 7495 sw
tri 1116 7459 1152 7495 ne
rect 1152 7482 1158 7495
tri 1158 7482 1171 7495 sw
rect 1152 7459 1171 7482
tri 986 7453 992 7459 sw
tri 1044 7453 1050 7459 ne
rect 1050 7453 1090 7459
tri 1090 7453 1096 7459 sw
tri 1152 7453 1158 7459 ne
rect 1158 7453 1171 7459
tri 1171 7453 1200 7482 sw
rect 954 7445 992 7453
tri 954 7429 970 7445 ne
rect 970 7429 992 7445
tri 992 7429 1016 7453 sw
tri 1050 7429 1074 7453 ne
rect 1074 7429 1096 7453
tri 1096 7429 1120 7453 sw
tri 1158 7440 1171 7453 ne
rect 1171 7452 1200 7453
tri 1200 7452 1201 7453 sw
tri 970 7413 986 7429 ne
rect 986 7413 1016 7429
tri 986 7383 1016 7413 ne
tri 1016 7407 1038 7429 sw
tri 1074 7407 1096 7429 ne
rect 1096 7407 1120 7429
tri 1120 7407 1142 7429 sw
rect 1016 7383 1038 7407
tri 1038 7383 1062 7407 sw
tri 1096 7393 1110 7407 ne
tri 1016 7369 1030 7383 ne
rect 1030 4044 1062 7383
rect 1110 4285 1142 7407
rect 1171 4377 1201 7452
rect 1230 4518 1262 7511
tri 1262 4518 1287 4543 sw
rect 1230 4486 1287 4518
tri 1230 4461 1255 4486 ne
tri 1201 4377 1226 4402 sw
rect 1171 4363 1226 4377
tri 1171 4338 1196 4363 ne
tri 1142 4285 1167 4310 sw
rect 1110 4253 1167 4285
tri 1110 4228 1135 4253 ne
tri 1110 3943 1135 3968 se
rect 1135 3943 1167 4253
rect 1110 3911 1167 3943
tri 1090 3776 1110 3796 se
rect 1110 3776 1142 3911
tri 1142 3886 1167 3911 nw
rect 1090 3770 1142 3776
rect 1090 3706 1142 3718
rect 1090 3648 1142 3654
tri 1171 3854 1196 3879 se
rect 1196 3854 1226 4363
rect 1171 3824 1226 3854
tri 1129 3595 1171 3637 se
rect 1171 3625 1201 3824
tri 1201 3799 1226 3824 nw
tri 1251 3799 1255 3803 se
rect 1255 3799 1287 4486
tri 1171 3595 1201 3625 nw
tri 1230 3778 1251 3799 se
rect 1251 3778 1287 3799
rect 1230 3746 1287 3778
tri 1087 3553 1129 3595 se
tri 1129 3553 1171 3595 nw
tri 1051 3517 1087 3553 se
rect 1087 3517 1093 3553
tri 1093 3517 1129 3553 nw
tri 1208 3517 1230 3539 se
rect 1230 3517 1262 3746
tri 1262 3721 1287 3746 nw
rect 8758 3699 8764 3751
rect 8816 3699 8828 3751
rect 8880 3699 9689 3751
tri 9606 3644 9661 3699 ne
rect 1051 3512 1088 3517
tri 1088 3512 1093 3517 nw
tri 1203 3512 1208 3517 se
rect 1208 3512 1262 3517
rect 1051 3460 1081 3512
tri 1081 3505 1088 3512 nw
tri 1081 3460 1084 3463 sw
rect 1134 3460 1140 3512
rect 1192 3460 1204 3512
rect 1256 3460 1262 3512
rect 1051 3459 1084 3460
tri 1084 3459 1085 3460 sw
rect 9505 3459 9511 3511
rect 9563 3459 9575 3511
rect 9627 3459 9633 3511
rect 1051 3432 1085 3459
tri 1085 3432 1112 3459 sw
tri 9578 3432 9605 3459 ne
rect 1051 3380 1079 3432
rect 1131 3380 1143 3432
rect 1195 3380 1201 3432
rect 9428 3379 9434 3431
rect 9486 3379 9498 3431
rect 9550 3384 9556 3431
tri 9556 3384 9571 3399 sw
rect 9550 3379 9571 3384
tri 9510 3346 9543 3379 ne
tri 9513 973 9543 1003 se
rect 9543 973 9571 3379
rect 9143 945 9571 973
rect 9143 710 9195 945
tri 9195 911 9229 945 nw
tri 9581 911 9605 935 se
rect 9605 911 9633 3459
tri 9575 905 9581 911 se
rect 9581 905 9633 911
rect 9143 646 9195 658
rect 9143 588 9195 594
rect 9475 877 9633 905
tri 9441 337 9475 371 se
rect 9475 337 9503 877
tri 9503 843 9537 877 nw
tri 9643 843 9661 861 se
rect 9661 843 9689 3699
tri 9627 827 9643 843 se
rect 9643 827 9689 843
rect 9602 795 9689 827
rect 9602 789 9654 795
tri 9654 761 9688 795 nw
rect 9602 725 9654 737
rect 9602 667 9654 673
rect 9354 285 9360 337
rect 9412 285 9445 337
rect 9497 285 9503 337
<< via2 >>
rect 15853 37999 15862 38048
rect 15862 37999 15909 38048
rect 15853 37992 15909 37999
rect 15853 37935 15862 37968
rect 15862 37935 15909 37968
rect 15853 37912 15909 37935
rect 15721 37049 15723 37091
rect 15723 37049 15775 37091
rect 15775 37049 15777 37091
rect 15721 37037 15777 37049
rect 15721 37035 15723 37037
rect 15723 37035 15775 37037
rect 15775 37035 15777 37037
rect 15721 36985 15723 37011
rect 15723 36985 15775 37011
rect 15775 36985 15777 37011
rect 15721 36955 15777 36985
<< metal3 >>
rect 15848 38048 15914 38053
rect 15848 37992 15853 38048
rect 15909 37992 15914 38048
rect 15848 37968 15914 37992
rect 15848 37912 15853 37968
rect 15909 37912 15914 37968
rect 15716 37091 15782 37107
rect 15716 37035 15721 37091
rect 15777 37035 15782 37091
rect 15716 37011 15782 37035
rect 15716 36955 15721 37011
rect 15777 36955 15782 37011
rect 15716 35292 15782 36955
rect 15848 35292 15914 37912
use sky130_fd_io__gpiov2_ictl_logic  sky130_fd_io__gpiov2_ictl_logic_0
timestamp 1619862920
transform -1 0 12264 0 -1 1116
box -34 10 3321 1116
use sky130_fd_io__gpiov2_buf_localesd  sky130_fd_io__gpiov2_buf_localesd_0
timestamp 1619862920
transform -1 0 3161 0 1 36196
box 146 0 3161 3800
use sky130_fd_io__gpiov2_ibuf_se  sky130_fd_io__gpiov2_ibuf_se_0
timestamp 1619862920
transform 1 0 3079 0 1 36000
box -467 -220 12925 4000
<< labels >>
flabel metal3 s 15726 35819 15775 36078 3 FreeSans 200 0 0 0 ENABLE_VDDIO_LV
port 1 nsew
flabel metal2 s 824 35975 904 36127 3 FreeSans 400 180 0 0 OUT_H
port 2 nsew
flabel metal2 s 1042 4136 1042 4136 0 FreeSans 200 90 0 0 MODE_VCCHIB_N
port 3 nsew
flabel metal1 s 10245 704 10245 704 0 FreeSans 200 90 0 0 MODE_VCCHIB_N
port 3 nsew
flabel metal1 s 15429 39770 15848 39986 3 FreeSans 400 180 0 0 VCCHIB
port 4 nsew
flabel metal1 s 3342 39782 3799 39961 3 FreeSans 400 180 0 0 VDDIO_Q
port 5 nsew
flabel metal1 s 911 35817 1231 36038 3 FreeSans 400 180 0 0 VSSD
port 6 nsew
flabel metal1 s 2702 36238 2938 36301 3 FreeSans 400 180 0 0 PAD
port 7 nsew
flabel metal1 s 15473 37934 15595 38006 3 FreeSans 400 180 0 0 OUT
port 8 nsew
flabel metal1 s 12069 729 12160 763 3 FreeSans 200 0 0 0 DM_H_N[1]
port 9 nsew
flabel metal1 s 11816 725 11876 762 3 FreeSans 200 0 0 0 DM_H_N[0]
port 10 nsew
flabel metal1 s 11416 728 11524 760 3 FreeSans 200 0 0 0 DM_H_N[2]
port 11 nsew
flabel metal1 s 10972 361 11001 477 3 FreeSans 200 0 0 0 INP_DIS_H_N
port 12 nsew
flabel metal1 s 10320 642 10351 759 3 FreeSans 200 0 0 0 IB_MODE_SEL_H
port 13 nsew
flabel metal1 s 9786 678 9818 789 3 FreeSans 200 0 0 0 IB_MODE_SEL_H_N
port 14 nsew
flabel metal1 s 9330 687 9363 788 3 FreeSans 200 0 0 0 VTRIP_SEL_H_N
port 15 nsew
flabel metal1 s 9334 910 9654 1086 3 FreeSans 400 180 0 0 VSSD
port 6 nsew
flabel metal1 s 10366 69 10823 248 3 FreeSans 400 180 0 0 VDDIO_Q
port 5 nsew
flabel comment s 13712 38624 13712 38624 0 FreeSans 440 0 0 0 LV_NET
flabel comment s 1148 35565 1148 35565 0 FreeSans 200 90 0 0 TRIPSEL_I_H_N
flabel comment s 1084 35565 1084 35565 0 FreeSans 200 90 0 0 VTRIP_SEL_H
flabel comment s 1026 35565 1026 35565 0 FreeSans 200 90 0 0 MODE_NORMAL_N
flabel comment s 967 35565 967 35565 0 FreeSans 200 90 0 0 MODE_VCCHIB_N
flabel comment s 15882 35630 15882 35630 0 FreeSans 400 0 0 0 OUT
flabel comment s 15740 35546 15740 35546 0 FreeSans 400 90 0 0 ENABLE_VDDIO_LV
flabel comment s 870 35708 870 35708 0 FreeSans 400 0 0 0 OUT_H
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 6287526
string GDS_START 6266328
<< end >>
