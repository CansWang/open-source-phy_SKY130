# Created by MC2 : Version 2013.12.00.f on 2020/05/11, 12:57:42

#*********************************************************************************************************************/
# Technology     : TSMC 16nm CMOS Logic FinFet Compact (FFC) Low Leakage HKMG  						*/
# Memory Type    : TSMC 16nm FFC High Density Single Port Single-Bank SRAM Compiler with d0734 bit cell	 				*/
# Library Name   : ts1n16ffcllsblvtc1024x144m4sw (user specify : ts1n16ffcllsblvtc1024x144m4sw)			*/
# Library Version: 130a												*/
# Generated Time : 2020/05/11, 12:57:39										*/
#*********************************************************************************************************************/
#															*/
# STATEMENT OF USE													*/
#															*/
# This information contains confidential and proprietary information of TSMC.					*/
# No part of this information may be reproduced, transmitted, transcribed,						*/
# stored in a retrieval system, or translated into any human or computer						*/
# language, in any form or by any means, electronic, mechanical, magnetic,						*/
# optical, chemical, manual, or otherwise, without the prior written permission					*/
# of TSMC. This information was prepared for informational purpose and is for					*/
# use by TSMC's customers only. TSMC reserves the right to make changes in the					*/
# information at any time and without notice.									*/
#															*/
#*********************************************************************************************************************/
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO TS1N16FFCLLSBLVTC1024X144M4SW
	CLASS BLOCK ;
	FOREIGN TS1N16FFCLLSBLVTC1024X144M4SW 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 64.175 BY 249.840 ;
	SYMMETRY X Y ;
	PIN A[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 120.200 64.175 120.280 ;
			LAYER M2 ;
			RECT 63.927 120.200 64.175 120.280 ;
			LAYER M3 ;
			RECT 63.927 120.200 64.175 120.280 ;
		END
		ANTENNAGATEAREA 0.006480 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.067800 LAYER M1 ;
		ANTENNAMAXAREACAR 4.009920 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.152040 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006480 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.075600 LAYER M2 ;
		ANTENNAMAXAREACAR 9.319320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.304200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006480 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.134280 LAYER M3 ;
		ANTENNAMAXAREACAR 21.482600 LAYER M3 ;
	END A[0]

	PIN A[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 118.856 64.175 118.936 ;
			LAYER M2 ;
			RECT 63.927 118.856 64.175 118.936 ;
			LAYER M3 ;
			RECT 63.927 118.856 64.175 118.936 ;
		END
		ANTENNAGATEAREA 0.006480 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.067800 LAYER M1 ;
		ANTENNAMAXAREACAR 4.009920 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.152040 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006480 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.075600 LAYER M2 ;
		ANTENNAMAXAREACAR 9.319320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.304200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006480 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.134280 LAYER M3 ;
		ANTENNAMAXAREACAR 21.482600 LAYER M3 ;
	END A[1]

	PIN A[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 129.224 64.175 129.304 ;
			LAYER M2 ;
			RECT 63.927 129.224 64.175 129.304 ;
			LAYER M3 ;
			RECT 63.927 129.224 64.175 129.304 ;
		END
		ANTENNAGATEAREA 0.006480 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.067800 LAYER M1 ;
		ANTENNAMAXAREACAR 4.009920 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.152040 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006480 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.075600 LAYER M2 ;
		ANTENNAMAXAREACAR 9.319320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.304200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006480 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.134280 LAYER M3 ;
		ANTENNAMAXAREACAR 21.482600 LAYER M3 ;
	END A[2]

	PIN A[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 128.456 64.175 128.536 ;
			LAYER M2 ;
			RECT 63.927 128.456 64.175 128.536 ;
			LAYER M3 ;
			RECT 63.927 128.456 64.175 128.536 ;
		END
		ANTENNAGATEAREA 0.006480 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.067800 LAYER M1 ;
		ANTENNAMAXAREACAR 4.009920 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.152040 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006480 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.075600 LAYER M2 ;
		ANTENNAMAXAREACAR 9.319320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.304200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006480 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.134280 LAYER M3 ;
		ANTENNAMAXAREACAR 21.482600 LAYER M3 ;
	END A[3]

	PIN A[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 127.880 64.175 127.960 ;
			LAYER M2 ;
			RECT 63.927 127.880 64.175 127.960 ;
			LAYER M3 ;
			RECT 63.927 127.880 64.175 127.960 ;
		END
		ANTENNAGATEAREA 0.006480 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.067800 LAYER M1 ;
		ANTENNAMAXAREACAR 4.009920 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.152040 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006480 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.075600 LAYER M2 ;
		ANTENNAMAXAREACAR 9.319320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.304200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006480 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.134280 LAYER M3 ;
		ANTENNAMAXAREACAR 21.482600 LAYER M3 ;
	END A[4]

	PIN A[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 125.192 64.175 125.272 ;
			LAYER M2 ;
			RECT 63.927 125.192 64.175 125.272 ;
			LAYER M3 ;
			RECT 63.927 125.192 64.175 125.272 ;
		END
		ANTENNAGATEAREA 0.006480 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.067800 LAYER M1 ;
		ANTENNAMAXAREACAR 4.009920 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.152040 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006480 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.075600 LAYER M2 ;
		ANTENNAMAXAREACAR 9.319320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.304200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006480 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.134280 LAYER M3 ;
		ANTENNAMAXAREACAR 21.482600 LAYER M3 ;
	END A[5]

	PIN A[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 125.960 64.175 126.040 ;
			LAYER M2 ;
			RECT 63.927 125.960 64.175 126.040 ;
			LAYER M3 ;
			RECT 63.927 125.960 64.175 126.040 ;
		END
		ANTENNAGATEAREA 0.006480 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.067800 LAYER M1 ;
		ANTENNAMAXAREACAR 4.009920 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.152040 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006480 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.075600 LAYER M2 ;
		ANTENNAMAXAREACAR 9.319320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.304200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006480 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.134280 LAYER M3 ;
		ANTENNAMAXAREACAR 21.482600 LAYER M3 ;
	END A[6]

	PIN A[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 127.112 64.175 127.192 ;
			LAYER M2 ;
			RECT 63.927 127.112 64.175 127.192 ;
			LAYER M3 ;
			RECT 63.927 127.112 64.175 127.192 ;
		END
		ANTENNAGATEAREA 0.006480 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.067800 LAYER M1 ;
		ANTENNAMAXAREACAR 4.009920 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.152040 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006480 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.075600 LAYER M2 ;
		ANTENNAMAXAREACAR 9.319320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.304200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006480 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.134280 LAYER M3 ;
		ANTENNAMAXAREACAR 21.482600 LAYER M3 ;
	END A[7]

	PIN A[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 121.736 64.175 121.816 ;
			LAYER M2 ;
			RECT 63.927 121.736 64.175 121.816 ;
			LAYER M3 ;
			RECT 63.927 121.736 64.175 121.816 ;
		END
		ANTENNAGATEAREA 0.006480 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.067800 LAYER M1 ;
		ANTENNAMAXAREACAR 4.009920 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.152040 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006480 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.075600 LAYER M2 ;
		ANTENNAMAXAREACAR 9.319320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.304200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006480 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.134280 LAYER M3 ;
		ANTENNAMAXAREACAR 21.482600 LAYER M3 ;
	END A[8]

	PIN A[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 120.392 64.175 120.472 ;
			LAYER M2 ;
			RECT 63.927 120.392 64.175 120.472 ;
			LAYER M3 ;
			RECT 63.927 120.392 64.175 120.472 ;
		END
		ANTENNAGATEAREA 0.006480 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.067800 LAYER M1 ;
		ANTENNAMAXAREACAR 4.009920 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.152040 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006480 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.075600 LAYER M2 ;
		ANTENNAMAXAREACAR 9.319320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.304200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006480 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.134280 LAYER M3 ;
		ANTENNAMAXAREACAR 21.482600 LAYER M3 ;
	END A[9]

	PIN BWEB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 2.120 64.175 2.200 ;
			LAYER M2 ;
			RECT 63.927 2.120 64.175 2.200 ;
			LAYER M3 ;
			RECT 63.927 2.120 64.175 2.200 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[0]

	PIN BWEB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 3.752 64.175 3.832 ;
			LAYER M2 ;
			RECT 63.927 3.752 64.175 3.832 ;
			LAYER M3 ;
			RECT 63.927 3.752 64.175 3.832 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[1]

	PIN BWEB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 5.384 64.175 5.464 ;
			LAYER M2 ;
			RECT 63.927 5.384 64.175 5.464 ;
			LAYER M3 ;
			RECT 63.927 5.384 64.175 5.464 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[2]

	PIN BWEB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 7.016 64.175 7.096 ;
			LAYER M2 ;
			RECT 63.927 7.016 64.175 7.096 ;
			LAYER M3 ;
			RECT 63.927 7.016 64.175 7.096 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[3]

	PIN BWEB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 8.648 64.175 8.728 ;
			LAYER M2 ;
			RECT 63.927 8.648 64.175 8.728 ;
			LAYER M3 ;
			RECT 63.927 8.648 64.175 8.728 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[4]

	PIN BWEB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 10.280 64.175 10.360 ;
			LAYER M2 ;
			RECT 63.927 10.280 64.175 10.360 ;
			LAYER M3 ;
			RECT 63.927 10.280 64.175 10.360 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[5]

	PIN BWEB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 11.912 64.175 11.992 ;
			LAYER M2 ;
			RECT 63.927 11.912 64.175 11.992 ;
			LAYER M3 ;
			RECT 63.927 11.912 64.175 11.992 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[6]

	PIN BWEB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 13.544 64.175 13.624 ;
			LAYER M2 ;
			RECT 63.927 13.544 64.175 13.624 ;
			LAYER M3 ;
			RECT 63.927 13.544 64.175 13.624 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[7]

	PIN BWEB[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 15.176 64.175 15.256 ;
			LAYER M2 ;
			RECT 63.927 15.176 64.175 15.256 ;
			LAYER M3 ;
			RECT 63.927 15.176 64.175 15.256 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[8]

	PIN BWEB[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 16.808 64.175 16.888 ;
			LAYER M2 ;
			RECT 63.927 16.808 64.175 16.888 ;
			LAYER M3 ;
			RECT 63.927 16.808 64.175 16.888 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[9]

	PIN BWEB[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 18.440 64.175 18.520 ;
			LAYER M2 ;
			RECT 63.927 18.440 64.175 18.520 ;
			LAYER M3 ;
			RECT 63.927 18.440 64.175 18.520 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[10]

	PIN BWEB[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 20.072 64.175 20.152 ;
			LAYER M2 ;
			RECT 63.927 20.072 64.175 20.152 ;
			LAYER M3 ;
			RECT 63.927 20.072 64.175 20.152 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[11]

	PIN BWEB[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 21.704 64.175 21.784 ;
			LAYER M2 ;
			RECT 63.927 21.704 64.175 21.784 ;
			LAYER M3 ;
			RECT 63.927 21.704 64.175 21.784 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[12]

	PIN BWEB[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 23.336 64.175 23.416 ;
			LAYER M2 ;
			RECT 63.927 23.336 64.175 23.416 ;
			LAYER M3 ;
			RECT 63.927 23.336 64.175 23.416 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[13]

	PIN BWEB[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 24.968 64.175 25.048 ;
			LAYER M2 ;
			RECT 63.927 24.968 64.175 25.048 ;
			LAYER M3 ;
			RECT 63.927 24.968 64.175 25.048 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[14]

	PIN BWEB[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 26.600 64.175 26.680 ;
			LAYER M2 ;
			RECT 63.927 26.600 64.175 26.680 ;
			LAYER M3 ;
			RECT 63.927 26.600 64.175 26.680 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[15]

	PIN BWEB[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 28.232 64.175 28.312 ;
			LAYER M2 ;
			RECT 63.927 28.232 64.175 28.312 ;
			LAYER M3 ;
			RECT 63.927 28.232 64.175 28.312 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[16]

	PIN BWEB[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 29.864 64.175 29.944 ;
			LAYER M2 ;
			RECT 63.927 29.864 64.175 29.944 ;
			LAYER M3 ;
			RECT 63.927 29.864 64.175 29.944 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[17]

	PIN BWEB[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 31.496 64.175 31.576 ;
			LAYER M2 ;
			RECT 63.927 31.496 64.175 31.576 ;
			LAYER M3 ;
			RECT 63.927 31.496 64.175 31.576 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[18]

	PIN BWEB[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 33.128 64.175 33.208 ;
			LAYER M2 ;
			RECT 63.927 33.128 64.175 33.208 ;
			LAYER M3 ;
			RECT 63.927 33.128 64.175 33.208 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[19]

	PIN BWEB[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 34.760 64.175 34.840 ;
			LAYER M2 ;
			RECT 63.927 34.760 64.175 34.840 ;
			LAYER M3 ;
			RECT 63.927 34.760 64.175 34.840 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[20]

	PIN BWEB[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 36.392 64.175 36.472 ;
			LAYER M2 ;
			RECT 63.927 36.392 64.175 36.472 ;
			LAYER M3 ;
			RECT 63.927 36.392 64.175 36.472 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[21]

	PIN BWEB[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 38.024 64.175 38.104 ;
			LAYER M2 ;
			RECT 63.927 38.024 64.175 38.104 ;
			LAYER M3 ;
			RECT 63.927 38.024 64.175 38.104 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[22]

	PIN BWEB[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 39.656 64.175 39.736 ;
			LAYER M2 ;
			RECT 63.927 39.656 64.175 39.736 ;
			LAYER M3 ;
			RECT 63.927 39.656 64.175 39.736 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[23]

	PIN BWEB[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 41.288 64.175 41.368 ;
			LAYER M2 ;
			RECT 63.927 41.288 64.175 41.368 ;
			LAYER M3 ;
			RECT 63.927 41.288 64.175 41.368 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[24]

	PIN BWEB[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 42.920 64.175 43.000 ;
			LAYER M2 ;
			RECT 63.927 42.920 64.175 43.000 ;
			LAYER M3 ;
			RECT 63.927 42.920 64.175 43.000 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[25]

	PIN BWEB[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 44.552 64.175 44.632 ;
			LAYER M2 ;
			RECT 63.927 44.552 64.175 44.632 ;
			LAYER M3 ;
			RECT 63.927 44.552 64.175 44.632 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[26]

	PIN BWEB[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 46.184 64.175 46.264 ;
			LAYER M2 ;
			RECT 63.927 46.184 64.175 46.264 ;
			LAYER M3 ;
			RECT 63.927 46.184 64.175 46.264 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[27]

	PIN BWEB[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 47.816 64.175 47.896 ;
			LAYER M2 ;
			RECT 63.927 47.816 64.175 47.896 ;
			LAYER M3 ;
			RECT 63.927 47.816 64.175 47.896 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[28]

	PIN BWEB[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 49.448 64.175 49.528 ;
			LAYER M2 ;
			RECT 63.927 49.448 64.175 49.528 ;
			LAYER M3 ;
			RECT 63.927 49.448 64.175 49.528 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[29]

	PIN BWEB[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 51.080 64.175 51.160 ;
			LAYER M2 ;
			RECT 63.927 51.080 64.175 51.160 ;
			LAYER M3 ;
			RECT 63.927 51.080 64.175 51.160 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[30]

	PIN BWEB[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 52.712 64.175 52.792 ;
			LAYER M2 ;
			RECT 63.927 52.712 64.175 52.792 ;
			LAYER M3 ;
			RECT 63.927 52.712 64.175 52.792 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[31]

	PIN BWEB[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 54.344 64.175 54.424 ;
			LAYER M2 ;
			RECT 63.927 54.344 64.175 54.424 ;
			LAYER M3 ;
			RECT 63.927 54.344 64.175 54.424 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[32]

	PIN BWEB[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 55.976 64.175 56.056 ;
			LAYER M2 ;
			RECT 63.927 55.976 64.175 56.056 ;
			LAYER M3 ;
			RECT 63.927 55.976 64.175 56.056 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[33]

	PIN BWEB[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 57.608 64.175 57.688 ;
			LAYER M2 ;
			RECT 63.927 57.608 64.175 57.688 ;
			LAYER M3 ;
			RECT 63.927 57.608 64.175 57.688 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[34]

	PIN BWEB[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 59.240 64.175 59.320 ;
			LAYER M2 ;
			RECT 63.927 59.240 64.175 59.320 ;
			LAYER M3 ;
			RECT 63.927 59.240 64.175 59.320 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[35]

	PIN BWEB[36]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 60.872 64.175 60.952 ;
			LAYER M2 ;
			RECT 63.927 60.872 64.175 60.952 ;
			LAYER M3 ;
			RECT 63.927 60.872 64.175 60.952 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[36]

	PIN BWEB[37]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 62.504 64.175 62.584 ;
			LAYER M2 ;
			RECT 63.927 62.504 64.175 62.584 ;
			LAYER M3 ;
			RECT 63.927 62.504 64.175 62.584 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[37]

	PIN BWEB[38]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 64.136 64.175 64.216 ;
			LAYER M2 ;
			RECT 63.927 64.136 64.175 64.216 ;
			LAYER M3 ;
			RECT 63.927 64.136 64.175 64.216 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[38]

	PIN BWEB[39]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 65.768 64.175 65.848 ;
			LAYER M2 ;
			RECT 63.927 65.768 64.175 65.848 ;
			LAYER M3 ;
			RECT 63.927 65.768 64.175 65.848 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[39]

	PIN BWEB[40]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 67.400 64.175 67.480 ;
			LAYER M2 ;
			RECT 63.927 67.400 64.175 67.480 ;
			LAYER M3 ;
			RECT 63.927 67.400 64.175 67.480 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[40]

	PIN BWEB[41]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 69.032 64.175 69.112 ;
			LAYER M2 ;
			RECT 63.927 69.032 64.175 69.112 ;
			LAYER M3 ;
			RECT 63.927 69.032 64.175 69.112 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[41]

	PIN BWEB[42]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 70.664 64.175 70.744 ;
			LAYER M2 ;
			RECT 63.927 70.664 64.175 70.744 ;
			LAYER M3 ;
			RECT 63.927 70.664 64.175 70.744 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[42]

	PIN BWEB[43]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 72.296 64.175 72.376 ;
			LAYER M2 ;
			RECT 63.927 72.296 64.175 72.376 ;
			LAYER M3 ;
			RECT 63.927 72.296 64.175 72.376 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[43]

	PIN BWEB[44]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 73.928 64.175 74.008 ;
			LAYER M2 ;
			RECT 63.927 73.928 64.175 74.008 ;
			LAYER M3 ;
			RECT 63.927 73.928 64.175 74.008 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[44]

	PIN BWEB[45]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 75.560 64.175 75.640 ;
			LAYER M2 ;
			RECT 63.927 75.560 64.175 75.640 ;
			LAYER M3 ;
			RECT 63.927 75.560 64.175 75.640 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[45]

	PIN BWEB[46]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 77.192 64.175 77.272 ;
			LAYER M2 ;
			RECT 63.927 77.192 64.175 77.272 ;
			LAYER M3 ;
			RECT 63.927 77.192 64.175 77.272 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[46]

	PIN BWEB[47]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 78.824 64.175 78.904 ;
			LAYER M2 ;
			RECT 63.927 78.824 64.175 78.904 ;
			LAYER M3 ;
			RECT 63.927 78.824 64.175 78.904 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[47]

	PIN BWEB[48]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 80.456 64.175 80.536 ;
			LAYER M2 ;
			RECT 63.927 80.456 64.175 80.536 ;
			LAYER M3 ;
			RECT 63.927 80.456 64.175 80.536 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[48]

	PIN BWEB[49]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 82.088 64.175 82.168 ;
			LAYER M2 ;
			RECT 63.927 82.088 64.175 82.168 ;
			LAYER M3 ;
			RECT 63.927 82.088 64.175 82.168 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[49]

	PIN BWEB[50]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 83.720 64.175 83.800 ;
			LAYER M2 ;
			RECT 63.927 83.720 64.175 83.800 ;
			LAYER M3 ;
			RECT 63.927 83.720 64.175 83.800 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[50]

	PIN BWEB[51]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 85.352 64.175 85.432 ;
			LAYER M2 ;
			RECT 63.927 85.352 64.175 85.432 ;
			LAYER M3 ;
			RECT 63.927 85.352 64.175 85.432 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[51]

	PIN BWEB[52]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 86.984 64.175 87.064 ;
			LAYER M2 ;
			RECT 63.927 86.984 64.175 87.064 ;
			LAYER M3 ;
			RECT 63.927 86.984 64.175 87.064 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[52]

	PIN BWEB[53]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 88.616 64.175 88.696 ;
			LAYER M2 ;
			RECT 63.927 88.616 64.175 88.696 ;
			LAYER M3 ;
			RECT 63.927 88.616 64.175 88.696 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[53]

	PIN BWEB[54]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 90.248 64.175 90.328 ;
			LAYER M2 ;
			RECT 63.927 90.248 64.175 90.328 ;
			LAYER M3 ;
			RECT 63.927 90.248 64.175 90.328 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[54]

	PIN BWEB[55]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 91.880 64.175 91.960 ;
			LAYER M2 ;
			RECT 63.927 91.880 64.175 91.960 ;
			LAYER M3 ;
			RECT 63.927 91.880 64.175 91.960 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[55]

	PIN BWEB[56]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 93.512 64.175 93.592 ;
			LAYER M2 ;
			RECT 63.927 93.512 64.175 93.592 ;
			LAYER M3 ;
			RECT 63.927 93.512 64.175 93.592 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[56]

	PIN BWEB[57]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 95.144 64.175 95.224 ;
			LAYER M2 ;
			RECT 63.927 95.144 64.175 95.224 ;
			LAYER M3 ;
			RECT 63.927 95.144 64.175 95.224 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[57]

	PIN BWEB[58]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 96.776 64.175 96.856 ;
			LAYER M2 ;
			RECT 63.927 96.776 64.175 96.856 ;
			LAYER M3 ;
			RECT 63.927 96.776 64.175 96.856 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[58]

	PIN BWEB[59]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 98.408 64.175 98.488 ;
			LAYER M2 ;
			RECT 63.927 98.408 64.175 98.488 ;
			LAYER M3 ;
			RECT 63.927 98.408 64.175 98.488 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[59]

	PIN BWEB[60]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 100.040 64.175 100.120 ;
			LAYER M2 ;
			RECT 63.927 100.040 64.175 100.120 ;
			LAYER M3 ;
			RECT 63.927 100.040 64.175 100.120 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[60]

	PIN BWEB[61]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 101.672 64.175 101.752 ;
			LAYER M2 ;
			RECT 63.927 101.672 64.175 101.752 ;
			LAYER M3 ;
			RECT 63.927 101.672 64.175 101.752 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[61]

	PIN BWEB[62]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 103.304 64.175 103.384 ;
			LAYER M2 ;
			RECT 63.927 103.304 64.175 103.384 ;
			LAYER M3 ;
			RECT 63.927 103.304 64.175 103.384 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[62]

	PIN BWEB[63]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 104.936 64.175 105.016 ;
			LAYER M2 ;
			RECT 63.927 104.936 64.175 105.016 ;
			LAYER M3 ;
			RECT 63.927 104.936 64.175 105.016 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[63]

	PIN BWEB[64]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 106.568 64.175 106.648 ;
			LAYER M2 ;
			RECT 63.927 106.568 64.175 106.648 ;
			LAYER M3 ;
			RECT 63.927 106.568 64.175 106.648 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[64]

	PIN BWEB[65]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 108.200 64.175 108.280 ;
			LAYER M2 ;
			RECT 63.927 108.200 64.175 108.280 ;
			LAYER M3 ;
			RECT 63.927 108.200 64.175 108.280 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[65]

	PIN BWEB[66]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 109.832 64.175 109.912 ;
			LAYER M2 ;
			RECT 63.927 109.832 64.175 109.912 ;
			LAYER M3 ;
			RECT 63.927 109.832 64.175 109.912 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[66]

	PIN BWEB[67]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 111.464 64.175 111.544 ;
			LAYER M2 ;
			RECT 63.927 111.464 64.175 111.544 ;
			LAYER M3 ;
			RECT 63.927 111.464 64.175 111.544 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[67]

	PIN BWEB[68]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 113.096 64.175 113.176 ;
			LAYER M2 ;
			RECT 63.927 113.096 64.175 113.176 ;
			LAYER M3 ;
			RECT 63.927 113.096 64.175 113.176 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[68]

	PIN BWEB[69]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 114.728 64.175 114.808 ;
			LAYER M2 ;
			RECT 63.927 114.728 64.175 114.808 ;
			LAYER M3 ;
			RECT 63.927 114.728 64.175 114.808 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[69]

	PIN BWEB[70]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 116.360 64.175 116.440 ;
			LAYER M2 ;
			RECT 63.927 116.360 64.175 116.440 ;
			LAYER M3 ;
			RECT 63.927 116.360 64.175 116.440 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[70]

	PIN BWEB[71]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 117.992 64.175 118.072 ;
			LAYER M2 ;
			RECT 63.927 117.992 64.175 118.072 ;
			LAYER M3 ;
			RECT 63.927 117.992 64.175 118.072 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[71]

	PIN BWEB[72]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 132.488 64.175 132.568 ;
			LAYER M2 ;
			RECT 63.927 132.488 64.175 132.568 ;
			LAYER M3 ;
			RECT 63.927 132.488 64.175 132.568 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[72]

	PIN BWEB[73]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 134.120 64.175 134.200 ;
			LAYER M2 ;
			RECT 63.927 134.120 64.175 134.200 ;
			LAYER M3 ;
			RECT 63.927 134.120 64.175 134.200 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[73]

	PIN BWEB[74]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 135.752 64.175 135.832 ;
			LAYER M2 ;
			RECT 63.927 135.752 64.175 135.832 ;
			LAYER M3 ;
			RECT 63.927 135.752 64.175 135.832 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[74]

	PIN BWEB[75]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 137.384 64.175 137.464 ;
			LAYER M2 ;
			RECT 63.927 137.384 64.175 137.464 ;
			LAYER M3 ;
			RECT 63.927 137.384 64.175 137.464 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[75]

	PIN BWEB[76]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 139.016 64.175 139.096 ;
			LAYER M2 ;
			RECT 63.927 139.016 64.175 139.096 ;
			LAYER M3 ;
			RECT 63.927 139.016 64.175 139.096 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[76]

	PIN BWEB[77]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 140.648 64.175 140.728 ;
			LAYER M2 ;
			RECT 63.927 140.648 64.175 140.728 ;
			LAYER M3 ;
			RECT 63.927 140.648 64.175 140.728 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[77]

	PIN BWEB[78]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 142.280 64.175 142.360 ;
			LAYER M2 ;
			RECT 63.927 142.280 64.175 142.360 ;
			LAYER M3 ;
			RECT 63.927 142.280 64.175 142.360 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[78]

	PIN BWEB[79]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 143.912 64.175 143.992 ;
			LAYER M2 ;
			RECT 63.927 143.912 64.175 143.992 ;
			LAYER M3 ;
			RECT 63.927 143.912 64.175 143.992 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[79]

	PIN BWEB[80]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 145.544 64.175 145.624 ;
			LAYER M2 ;
			RECT 63.927 145.544 64.175 145.624 ;
			LAYER M3 ;
			RECT 63.927 145.544 64.175 145.624 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[80]

	PIN BWEB[81]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 147.176 64.175 147.256 ;
			LAYER M2 ;
			RECT 63.927 147.176 64.175 147.256 ;
			LAYER M3 ;
			RECT 63.927 147.176 64.175 147.256 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[81]

	PIN BWEB[82]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 148.808 64.175 148.888 ;
			LAYER M2 ;
			RECT 63.927 148.808 64.175 148.888 ;
			LAYER M3 ;
			RECT 63.927 148.808 64.175 148.888 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[82]

	PIN BWEB[83]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 150.440 64.175 150.520 ;
			LAYER M2 ;
			RECT 63.927 150.440 64.175 150.520 ;
			LAYER M3 ;
			RECT 63.927 150.440 64.175 150.520 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[83]

	PIN BWEB[84]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 152.072 64.175 152.152 ;
			LAYER M2 ;
			RECT 63.927 152.072 64.175 152.152 ;
			LAYER M3 ;
			RECT 63.927 152.072 64.175 152.152 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[84]

	PIN BWEB[85]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 153.704 64.175 153.784 ;
			LAYER M2 ;
			RECT 63.927 153.704 64.175 153.784 ;
			LAYER M3 ;
			RECT 63.927 153.704 64.175 153.784 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[85]

	PIN BWEB[86]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 155.336 64.175 155.416 ;
			LAYER M2 ;
			RECT 63.927 155.336 64.175 155.416 ;
			LAYER M3 ;
			RECT 63.927 155.336 64.175 155.416 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[86]

	PIN BWEB[87]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 156.968 64.175 157.048 ;
			LAYER M2 ;
			RECT 63.927 156.968 64.175 157.048 ;
			LAYER M3 ;
			RECT 63.927 156.968 64.175 157.048 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[87]

	PIN BWEB[88]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 158.600 64.175 158.680 ;
			LAYER M2 ;
			RECT 63.927 158.600 64.175 158.680 ;
			LAYER M3 ;
			RECT 63.927 158.600 64.175 158.680 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[88]

	PIN BWEB[89]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 160.232 64.175 160.312 ;
			LAYER M2 ;
			RECT 63.927 160.232 64.175 160.312 ;
			LAYER M3 ;
			RECT 63.927 160.232 64.175 160.312 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[89]

	PIN BWEB[90]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 161.864 64.175 161.944 ;
			LAYER M2 ;
			RECT 63.927 161.864 64.175 161.944 ;
			LAYER M3 ;
			RECT 63.927 161.864 64.175 161.944 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[90]

	PIN BWEB[91]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 163.496 64.175 163.576 ;
			LAYER M2 ;
			RECT 63.927 163.496 64.175 163.576 ;
			LAYER M3 ;
			RECT 63.927 163.496 64.175 163.576 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[91]

	PIN BWEB[92]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 165.128 64.175 165.208 ;
			LAYER M2 ;
			RECT 63.927 165.128 64.175 165.208 ;
			LAYER M3 ;
			RECT 63.927 165.128 64.175 165.208 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[92]

	PIN BWEB[93]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 166.760 64.175 166.840 ;
			LAYER M2 ;
			RECT 63.927 166.760 64.175 166.840 ;
			LAYER M3 ;
			RECT 63.927 166.760 64.175 166.840 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[93]

	PIN BWEB[94]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 168.392 64.175 168.472 ;
			LAYER M2 ;
			RECT 63.927 168.392 64.175 168.472 ;
			LAYER M3 ;
			RECT 63.927 168.392 64.175 168.472 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[94]

	PIN BWEB[95]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 170.024 64.175 170.104 ;
			LAYER M2 ;
			RECT 63.927 170.024 64.175 170.104 ;
			LAYER M3 ;
			RECT 63.927 170.024 64.175 170.104 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[95]

	PIN BWEB[96]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 171.656 64.175 171.736 ;
			LAYER M2 ;
			RECT 63.927 171.656 64.175 171.736 ;
			LAYER M3 ;
			RECT 63.927 171.656 64.175 171.736 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[96]

	PIN BWEB[97]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 173.288 64.175 173.368 ;
			LAYER M2 ;
			RECT 63.927 173.288 64.175 173.368 ;
			LAYER M3 ;
			RECT 63.927 173.288 64.175 173.368 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[97]

	PIN BWEB[98]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 174.920 64.175 175.000 ;
			LAYER M2 ;
			RECT 63.927 174.920 64.175 175.000 ;
			LAYER M3 ;
			RECT 63.927 174.920 64.175 175.000 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[98]

	PIN BWEB[99]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 176.552 64.175 176.632 ;
			LAYER M2 ;
			RECT 63.927 176.552 64.175 176.632 ;
			LAYER M3 ;
			RECT 63.927 176.552 64.175 176.632 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[99]

	PIN BWEB[100]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 178.184 64.175 178.264 ;
			LAYER M2 ;
			RECT 63.927 178.184 64.175 178.264 ;
			LAYER M3 ;
			RECT 63.927 178.184 64.175 178.264 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[100]

	PIN BWEB[101]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 179.816 64.175 179.896 ;
			LAYER M2 ;
			RECT 63.927 179.816 64.175 179.896 ;
			LAYER M3 ;
			RECT 63.927 179.816 64.175 179.896 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[101]

	PIN BWEB[102]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 181.448 64.175 181.528 ;
			LAYER M2 ;
			RECT 63.927 181.448 64.175 181.528 ;
			LAYER M3 ;
			RECT 63.927 181.448 64.175 181.528 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[102]

	PIN BWEB[103]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 183.080 64.175 183.160 ;
			LAYER M2 ;
			RECT 63.927 183.080 64.175 183.160 ;
			LAYER M3 ;
			RECT 63.927 183.080 64.175 183.160 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[103]

	PIN BWEB[104]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 184.712 64.175 184.792 ;
			LAYER M2 ;
			RECT 63.927 184.712 64.175 184.792 ;
			LAYER M3 ;
			RECT 63.927 184.712 64.175 184.792 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[104]

	PIN BWEB[105]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 186.344 64.175 186.424 ;
			LAYER M2 ;
			RECT 63.927 186.344 64.175 186.424 ;
			LAYER M3 ;
			RECT 63.927 186.344 64.175 186.424 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[105]

	PIN BWEB[106]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 187.976 64.175 188.056 ;
			LAYER M2 ;
			RECT 63.927 187.976 64.175 188.056 ;
			LAYER M3 ;
			RECT 63.927 187.976 64.175 188.056 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[106]

	PIN BWEB[107]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 189.608 64.175 189.688 ;
			LAYER M2 ;
			RECT 63.927 189.608 64.175 189.688 ;
			LAYER M3 ;
			RECT 63.927 189.608 64.175 189.688 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[107]

	PIN BWEB[108]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 191.240 64.175 191.320 ;
			LAYER M2 ;
			RECT 63.927 191.240 64.175 191.320 ;
			LAYER M3 ;
			RECT 63.927 191.240 64.175 191.320 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[108]

	PIN BWEB[109]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 192.872 64.175 192.952 ;
			LAYER M2 ;
			RECT 63.927 192.872 64.175 192.952 ;
			LAYER M3 ;
			RECT 63.927 192.872 64.175 192.952 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[109]

	PIN BWEB[110]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 194.504 64.175 194.584 ;
			LAYER M2 ;
			RECT 63.927 194.504 64.175 194.584 ;
			LAYER M3 ;
			RECT 63.927 194.504 64.175 194.584 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[110]

	PIN BWEB[111]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 196.136 64.175 196.216 ;
			LAYER M2 ;
			RECT 63.927 196.136 64.175 196.216 ;
			LAYER M3 ;
			RECT 63.927 196.136 64.175 196.216 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[111]

	PIN BWEB[112]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 197.768 64.175 197.848 ;
			LAYER M2 ;
			RECT 63.927 197.768 64.175 197.848 ;
			LAYER M3 ;
			RECT 63.927 197.768 64.175 197.848 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[112]

	PIN BWEB[113]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 199.400 64.175 199.480 ;
			LAYER M2 ;
			RECT 63.927 199.400 64.175 199.480 ;
			LAYER M3 ;
			RECT 63.927 199.400 64.175 199.480 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[113]

	PIN BWEB[114]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 201.032 64.175 201.112 ;
			LAYER M2 ;
			RECT 63.927 201.032 64.175 201.112 ;
			LAYER M3 ;
			RECT 63.927 201.032 64.175 201.112 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[114]

	PIN BWEB[115]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 202.664 64.175 202.744 ;
			LAYER M2 ;
			RECT 63.927 202.664 64.175 202.744 ;
			LAYER M3 ;
			RECT 63.927 202.664 64.175 202.744 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[115]

	PIN BWEB[116]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 204.296 64.175 204.376 ;
			LAYER M2 ;
			RECT 63.927 204.296 64.175 204.376 ;
			LAYER M3 ;
			RECT 63.927 204.296 64.175 204.376 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[116]

	PIN BWEB[117]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 205.928 64.175 206.008 ;
			LAYER M2 ;
			RECT 63.927 205.928 64.175 206.008 ;
			LAYER M3 ;
			RECT 63.927 205.928 64.175 206.008 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[117]

	PIN BWEB[118]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 207.560 64.175 207.640 ;
			LAYER M2 ;
			RECT 63.927 207.560 64.175 207.640 ;
			LAYER M3 ;
			RECT 63.927 207.560 64.175 207.640 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[118]

	PIN BWEB[119]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 209.192 64.175 209.272 ;
			LAYER M2 ;
			RECT 63.927 209.192 64.175 209.272 ;
			LAYER M3 ;
			RECT 63.927 209.192 64.175 209.272 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[119]

	PIN BWEB[120]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 210.824 64.175 210.904 ;
			LAYER M2 ;
			RECT 63.927 210.824 64.175 210.904 ;
			LAYER M3 ;
			RECT 63.927 210.824 64.175 210.904 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[120]

	PIN BWEB[121]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 212.456 64.175 212.536 ;
			LAYER M2 ;
			RECT 63.927 212.456 64.175 212.536 ;
			LAYER M3 ;
			RECT 63.927 212.456 64.175 212.536 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[121]

	PIN BWEB[122]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 214.088 64.175 214.168 ;
			LAYER M2 ;
			RECT 63.927 214.088 64.175 214.168 ;
			LAYER M3 ;
			RECT 63.927 214.088 64.175 214.168 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[122]

	PIN BWEB[123]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 215.720 64.175 215.800 ;
			LAYER M2 ;
			RECT 63.927 215.720 64.175 215.800 ;
			LAYER M3 ;
			RECT 63.927 215.720 64.175 215.800 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[123]

	PIN BWEB[124]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 217.352 64.175 217.432 ;
			LAYER M2 ;
			RECT 63.927 217.352 64.175 217.432 ;
			LAYER M3 ;
			RECT 63.927 217.352 64.175 217.432 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[124]

	PIN BWEB[125]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 218.984 64.175 219.064 ;
			LAYER M2 ;
			RECT 63.927 218.984 64.175 219.064 ;
			LAYER M3 ;
			RECT 63.927 218.984 64.175 219.064 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[125]

	PIN BWEB[126]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 220.616 64.175 220.696 ;
			LAYER M2 ;
			RECT 63.927 220.616 64.175 220.696 ;
			LAYER M3 ;
			RECT 63.927 220.616 64.175 220.696 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[126]

	PIN BWEB[127]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 222.248 64.175 222.328 ;
			LAYER M2 ;
			RECT 63.927 222.248 64.175 222.328 ;
			LAYER M3 ;
			RECT 63.927 222.248 64.175 222.328 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[127]

	PIN BWEB[128]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 223.880 64.175 223.960 ;
			LAYER M2 ;
			RECT 63.927 223.880 64.175 223.960 ;
			LAYER M3 ;
			RECT 63.927 223.880 64.175 223.960 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[128]

	PIN BWEB[129]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 225.512 64.175 225.592 ;
			LAYER M2 ;
			RECT 63.927 225.512 64.175 225.592 ;
			LAYER M3 ;
			RECT 63.927 225.512 64.175 225.592 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[129]

	PIN BWEB[130]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 227.144 64.175 227.224 ;
			LAYER M2 ;
			RECT 63.927 227.144 64.175 227.224 ;
			LAYER M3 ;
			RECT 63.927 227.144 64.175 227.224 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[130]

	PIN BWEB[131]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 228.776 64.175 228.856 ;
			LAYER M2 ;
			RECT 63.927 228.776 64.175 228.856 ;
			LAYER M3 ;
			RECT 63.927 228.776 64.175 228.856 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[131]

	PIN BWEB[132]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 230.408 64.175 230.488 ;
			LAYER M2 ;
			RECT 63.927 230.408 64.175 230.488 ;
			LAYER M3 ;
			RECT 63.927 230.408 64.175 230.488 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[132]

	PIN BWEB[133]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 232.040 64.175 232.120 ;
			LAYER M2 ;
			RECT 63.927 232.040 64.175 232.120 ;
			LAYER M3 ;
			RECT 63.927 232.040 64.175 232.120 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[133]

	PIN BWEB[134]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 233.672 64.175 233.752 ;
			LAYER M2 ;
			RECT 63.927 233.672 64.175 233.752 ;
			LAYER M3 ;
			RECT 63.927 233.672 64.175 233.752 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[134]

	PIN BWEB[135]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 235.304 64.175 235.384 ;
			LAYER M2 ;
			RECT 63.927 235.304 64.175 235.384 ;
			LAYER M3 ;
			RECT 63.927 235.304 64.175 235.384 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[135]

	PIN BWEB[136]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 236.936 64.175 237.016 ;
			LAYER M2 ;
			RECT 63.927 236.936 64.175 237.016 ;
			LAYER M3 ;
			RECT 63.927 236.936 64.175 237.016 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[136]

	PIN BWEB[137]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 238.568 64.175 238.648 ;
			LAYER M2 ;
			RECT 63.927 238.568 64.175 238.648 ;
			LAYER M3 ;
			RECT 63.927 238.568 64.175 238.648 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[137]

	PIN BWEB[138]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 240.200 64.175 240.280 ;
			LAYER M2 ;
			RECT 63.927 240.200 64.175 240.280 ;
			LAYER M3 ;
			RECT 63.927 240.200 64.175 240.280 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[138]

	PIN BWEB[139]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 241.832 64.175 241.912 ;
			LAYER M2 ;
			RECT 63.927 241.832 64.175 241.912 ;
			LAYER M3 ;
			RECT 63.927 241.832 64.175 241.912 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[139]

	PIN BWEB[140]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 243.464 64.175 243.544 ;
			LAYER M2 ;
			RECT 63.927 243.464 64.175 243.544 ;
			LAYER M3 ;
			RECT 63.927 243.464 64.175 243.544 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[140]

	PIN BWEB[141]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 245.096 64.175 245.176 ;
			LAYER M2 ;
			RECT 63.927 245.096 64.175 245.176 ;
			LAYER M3 ;
			RECT 63.927 245.096 64.175 245.176 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[141]

	PIN BWEB[142]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 246.728 64.175 246.808 ;
			LAYER M2 ;
			RECT 63.927 246.728 64.175 246.808 ;
			LAYER M3 ;
			RECT 63.927 246.728 64.175 246.808 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[142]

	PIN BWEB[143]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 248.360 64.175 248.440 ;
			LAYER M2 ;
			RECT 63.927 248.360 64.175 248.440 ;
			LAYER M3 ;
			RECT 63.927 248.360 64.175 248.440 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.072960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.598900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.104640 LAYER M2 ;
		ANTENNAMAXAREACAR 22.892000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.154080 LAYER M3 ;
		ANTENNAMAXAREACAR 89.305900 LAYER M3 ;
	END BWEB[143]

	PIN CEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 121.928 64.175 122.008 ;
			LAYER M2 ;
			RECT 63.927 121.928 64.175 122.008 ;
			LAYER M3 ;
			RECT 63.927 121.928 64.175 122.008 ;
		END
		ANTENNAGATEAREA 0.008000 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.067560 LAYER M1 ;
		ANTENNAMAXAREACAR 3.216000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.122880 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008000 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.089760 LAYER M2 ;
		ANTENNAMAXAREACAR 7.464000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.245760 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008000 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.109800 LAYER M3 ;
		ANTENNAMAXAREACAR 15.642000 LAYER M3 ;
	END CEB

	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 124.232 64.175 124.312 ;
			LAYER M2 ;
			RECT 63.927 124.232 64.175 124.312 ;
			LAYER M3 ;
			RECT 63.927 124.232 64.175 124.312 ;
		END
		ANTENNAGATEAREA 0.014160 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.083640 LAYER M1 ;
		ANTENNAMAXAREACAR 2.732280 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.069480 LAYER VIA1 ;
		ANTENNAGATEAREA 0.014160 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.449760 LAYER M2 ;
		ANTENNAMAXAREACAR 25.547500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.243240 LAYER VIA2 ;
		ANTENNAGATEAREA 0.014160 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.503600 LAYER M3 ;
		ANTENNAMAXAREACAR 110.593000 LAYER M3 ;
	END CLK

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 1.448 64.175 1.528 ;
			LAYER M2 ;
			RECT 63.927 1.448 64.175 1.528 ;
			LAYER M3 ;
			RECT 63.927 1.448 64.175 1.528 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[0]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 3.080 64.175 3.160 ;
			LAYER M2 ;
			RECT 63.927 3.080 64.175 3.160 ;
			LAYER M3 ;
			RECT 63.927 3.080 64.175 3.160 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[1]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 4.712 64.175 4.792 ;
			LAYER M2 ;
			RECT 63.927 4.712 64.175 4.792 ;
			LAYER M3 ;
			RECT 63.927 4.712 64.175 4.792 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[2]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 6.344 64.175 6.424 ;
			LAYER M2 ;
			RECT 63.927 6.344 64.175 6.424 ;
			LAYER M3 ;
			RECT 63.927 6.344 64.175 6.424 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[3]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 7.976 64.175 8.056 ;
			LAYER M2 ;
			RECT 63.927 7.976 64.175 8.056 ;
			LAYER M3 ;
			RECT 63.927 7.976 64.175 8.056 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[4]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 9.608 64.175 9.688 ;
			LAYER M2 ;
			RECT 63.927 9.608 64.175 9.688 ;
			LAYER M3 ;
			RECT 63.927 9.608 64.175 9.688 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[5]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 11.240 64.175 11.320 ;
			LAYER M2 ;
			RECT 63.927 11.240 64.175 11.320 ;
			LAYER M3 ;
			RECT 63.927 11.240 64.175 11.320 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 12.872 64.175 12.952 ;
			LAYER M2 ;
			RECT 63.927 12.872 64.175 12.952 ;
			LAYER M3 ;
			RECT 63.927 12.872 64.175 12.952 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[7]

	PIN D[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 14.504 64.175 14.584 ;
			LAYER M2 ;
			RECT 63.927 14.504 64.175 14.584 ;
			LAYER M3 ;
			RECT 63.927 14.504 64.175 14.584 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[8]

	PIN D[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 16.136 64.175 16.216 ;
			LAYER M2 ;
			RECT 63.927 16.136 64.175 16.216 ;
			LAYER M3 ;
			RECT 63.927 16.136 64.175 16.216 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[9]

	PIN D[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 17.768 64.175 17.848 ;
			LAYER M2 ;
			RECT 63.927 17.768 64.175 17.848 ;
			LAYER M3 ;
			RECT 63.927 17.768 64.175 17.848 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[10]

	PIN D[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 19.400 64.175 19.480 ;
			LAYER M2 ;
			RECT 63.927 19.400 64.175 19.480 ;
			LAYER M3 ;
			RECT 63.927 19.400 64.175 19.480 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[11]

	PIN D[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 21.032 64.175 21.112 ;
			LAYER M2 ;
			RECT 63.927 21.032 64.175 21.112 ;
			LAYER M3 ;
			RECT 63.927 21.032 64.175 21.112 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[12]

	PIN D[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 22.664 64.175 22.744 ;
			LAYER M2 ;
			RECT 63.927 22.664 64.175 22.744 ;
			LAYER M3 ;
			RECT 63.927 22.664 64.175 22.744 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[13]

	PIN D[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 24.296 64.175 24.376 ;
			LAYER M2 ;
			RECT 63.927 24.296 64.175 24.376 ;
			LAYER M3 ;
			RECT 63.927 24.296 64.175 24.376 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[14]

	PIN D[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 25.928 64.175 26.008 ;
			LAYER M2 ;
			RECT 63.927 25.928 64.175 26.008 ;
			LAYER M3 ;
			RECT 63.927 25.928 64.175 26.008 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[15]

	PIN D[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 27.560 64.175 27.640 ;
			LAYER M2 ;
			RECT 63.927 27.560 64.175 27.640 ;
			LAYER M3 ;
			RECT 63.927 27.560 64.175 27.640 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[16]

	PIN D[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 29.192 64.175 29.272 ;
			LAYER M2 ;
			RECT 63.927 29.192 64.175 29.272 ;
			LAYER M3 ;
			RECT 63.927 29.192 64.175 29.272 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[17]

	PIN D[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 30.824 64.175 30.904 ;
			LAYER M2 ;
			RECT 63.927 30.824 64.175 30.904 ;
			LAYER M3 ;
			RECT 63.927 30.824 64.175 30.904 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[18]

	PIN D[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 32.456 64.175 32.536 ;
			LAYER M2 ;
			RECT 63.927 32.456 64.175 32.536 ;
			LAYER M3 ;
			RECT 63.927 32.456 64.175 32.536 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[19]

	PIN D[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 34.088 64.175 34.168 ;
			LAYER M2 ;
			RECT 63.927 34.088 64.175 34.168 ;
			LAYER M3 ;
			RECT 63.927 34.088 64.175 34.168 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[20]

	PIN D[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 35.720 64.175 35.800 ;
			LAYER M2 ;
			RECT 63.927 35.720 64.175 35.800 ;
			LAYER M3 ;
			RECT 63.927 35.720 64.175 35.800 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[21]

	PIN D[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 37.352 64.175 37.432 ;
			LAYER M2 ;
			RECT 63.927 37.352 64.175 37.432 ;
			LAYER M3 ;
			RECT 63.927 37.352 64.175 37.432 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[22]

	PIN D[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 38.984 64.175 39.064 ;
			LAYER M2 ;
			RECT 63.927 38.984 64.175 39.064 ;
			LAYER M3 ;
			RECT 63.927 38.984 64.175 39.064 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[23]

	PIN D[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 40.616 64.175 40.696 ;
			LAYER M2 ;
			RECT 63.927 40.616 64.175 40.696 ;
			LAYER M3 ;
			RECT 63.927 40.616 64.175 40.696 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[24]

	PIN D[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 42.248 64.175 42.328 ;
			LAYER M2 ;
			RECT 63.927 42.248 64.175 42.328 ;
			LAYER M3 ;
			RECT 63.927 42.248 64.175 42.328 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[25]

	PIN D[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 43.880 64.175 43.960 ;
			LAYER M2 ;
			RECT 63.927 43.880 64.175 43.960 ;
			LAYER M3 ;
			RECT 63.927 43.880 64.175 43.960 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[26]

	PIN D[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 45.512 64.175 45.592 ;
			LAYER M2 ;
			RECT 63.927 45.512 64.175 45.592 ;
			LAYER M3 ;
			RECT 63.927 45.512 64.175 45.592 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[27]

	PIN D[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 47.144 64.175 47.224 ;
			LAYER M2 ;
			RECT 63.927 47.144 64.175 47.224 ;
			LAYER M3 ;
			RECT 63.927 47.144 64.175 47.224 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[28]

	PIN D[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 48.776 64.175 48.856 ;
			LAYER M2 ;
			RECT 63.927 48.776 64.175 48.856 ;
			LAYER M3 ;
			RECT 63.927 48.776 64.175 48.856 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[29]

	PIN D[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 50.408 64.175 50.488 ;
			LAYER M2 ;
			RECT 63.927 50.408 64.175 50.488 ;
			LAYER M3 ;
			RECT 63.927 50.408 64.175 50.488 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[30]

	PIN D[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 52.040 64.175 52.120 ;
			LAYER M2 ;
			RECT 63.927 52.040 64.175 52.120 ;
			LAYER M3 ;
			RECT 63.927 52.040 64.175 52.120 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[31]

	PIN D[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 53.672 64.175 53.752 ;
			LAYER M2 ;
			RECT 63.927 53.672 64.175 53.752 ;
			LAYER M3 ;
			RECT 63.927 53.672 64.175 53.752 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[32]

	PIN D[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 55.304 64.175 55.384 ;
			LAYER M2 ;
			RECT 63.927 55.304 64.175 55.384 ;
			LAYER M3 ;
			RECT 63.927 55.304 64.175 55.384 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[33]

	PIN D[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 56.936 64.175 57.016 ;
			LAYER M2 ;
			RECT 63.927 56.936 64.175 57.016 ;
			LAYER M3 ;
			RECT 63.927 56.936 64.175 57.016 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[34]

	PIN D[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 58.568 64.175 58.648 ;
			LAYER M2 ;
			RECT 63.927 58.568 64.175 58.648 ;
			LAYER M3 ;
			RECT 63.927 58.568 64.175 58.648 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[35]

	PIN D[36]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 60.200 64.175 60.280 ;
			LAYER M2 ;
			RECT 63.927 60.200 64.175 60.280 ;
			LAYER M3 ;
			RECT 63.927 60.200 64.175 60.280 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[36]

	PIN D[37]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 61.832 64.175 61.912 ;
			LAYER M2 ;
			RECT 63.927 61.832 64.175 61.912 ;
			LAYER M3 ;
			RECT 63.927 61.832 64.175 61.912 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[37]

	PIN D[38]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 63.464 64.175 63.544 ;
			LAYER M2 ;
			RECT 63.927 63.464 64.175 63.544 ;
			LAYER M3 ;
			RECT 63.927 63.464 64.175 63.544 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[38]

	PIN D[39]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 65.096 64.175 65.176 ;
			LAYER M2 ;
			RECT 63.927 65.096 64.175 65.176 ;
			LAYER M3 ;
			RECT 63.927 65.096 64.175 65.176 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[39]

	PIN D[40]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 66.728 64.175 66.808 ;
			LAYER M2 ;
			RECT 63.927 66.728 64.175 66.808 ;
			LAYER M3 ;
			RECT 63.927 66.728 64.175 66.808 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[40]

	PIN D[41]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 68.360 64.175 68.440 ;
			LAYER M2 ;
			RECT 63.927 68.360 64.175 68.440 ;
			LAYER M3 ;
			RECT 63.927 68.360 64.175 68.440 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[41]

	PIN D[42]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 69.992 64.175 70.072 ;
			LAYER M2 ;
			RECT 63.927 69.992 64.175 70.072 ;
			LAYER M3 ;
			RECT 63.927 69.992 64.175 70.072 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[42]

	PIN D[43]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 71.624 64.175 71.704 ;
			LAYER M2 ;
			RECT 63.927 71.624 64.175 71.704 ;
			LAYER M3 ;
			RECT 63.927 71.624 64.175 71.704 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[43]

	PIN D[44]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 73.256 64.175 73.336 ;
			LAYER M2 ;
			RECT 63.927 73.256 64.175 73.336 ;
			LAYER M3 ;
			RECT 63.927 73.256 64.175 73.336 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[44]

	PIN D[45]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 74.888 64.175 74.968 ;
			LAYER M2 ;
			RECT 63.927 74.888 64.175 74.968 ;
			LAYER M3 ;
			RECT 63.927 74.888 64.175 74.968 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[45]

	PIN D[46]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 76.520 64.175 76.600 ;
			LAYER M2 ;
			RECT 63.927 76.520 64.175 76.600 ;
			LAYER M3 ;
			RECT 63.927 76.520 64.175 76.600 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[46]

	PIN D[47]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 78.152 64.175 78.232 ;
			LAYER M2 ;
			RECT 63.927 78.152 64.175 78.232 ;
			LAYER M3 ;
			RECT 63.927 78.152 64.175 78.232 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[47]

	PIN D[48]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 79.784 64.175 79.864 ;
			LAYER M2 ;
			RECT 63.927 79.784 64.175 79.864 ;
			LAYER M3 ;
			RECT 63.927 79.784 64.175 79.864 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[48]

	PIN D[49]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 81.416 64.175 81.496 ;
			LAYER M2 ;
			RECT 63.927 81.416 64.175 81.496 ;
			LAYER M3 ;
			RECT 63.927 81.416 64.175 81.496 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[49]

	PIN D[50]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 83.048 64.175 83.128 ;
			LAYER M2 ;
			RECT 63.927 83.048 64.175 83.128 ;
			LAYER M3 ;
			RECT 63.927 83.048 64.175 83.128 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[50]

	PIN D[51]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 84.680 64.175 84.760 ;
			LAYER M2 ;
			RECT 63.927 84.680 64.175 84.760 ;
			LAYER M3 ;
			RECT 63.927 84.680 64.175 84.760 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[51]

	PIN D[52]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 86.312 64.175 86.392 ;
			LAYER M2 ;
			RECT 63.927 86.312 64.175 86.392 ;
			LAYER M3 ;
			RECT 63.927 86.312 64.175 86.392 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[52]

	PIN D[53]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 87.944 64.175 88.024 ;
			LAYER M2 ;
			RECT 63.927 87.944 64.175 88.024 ;
			LAYER M3 ;
			RECT 63.927 87.944 64.175 88.024 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[53]

	PIN D[54]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 89.576 64.175 89.656 ;
			LAYER M2 ;
			RECT 63.927 89.576 64.175 89.656 ;
			LAYER M3 ;
			RECT 63.927 89.576 64.175 89.656 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[54]

	PIN D[55]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 91.208 64.175 91.288 ;
			LAYER M2 ;
			RECT 63.927 91.208 64.175 91.288 ;
			LAYER M3 ;
			RECT 63.927 91.208 64.175 91.288 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[55]

	PIN D[56]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 92.840 64.175 92.920 ;
			LAYER M2 ;
			RECT 63.927 92.840 64.175 92.920 ;
			LAYER M3 ;
			RECT 63.927 92.840 64.175 92.920 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[56]

	PIN D[57]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 94.472 64.175 94.552 ;
			LAYER M2 ;
			RECT 63.927 94.472 64.175 94.552 ;
			LAYER M3 ;
			RECT 63.927 94.472 64.175 94.552 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[57]

	PIN D[58]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 96.104 64.175 96.184 ;
			LAYER M2 ;
			RECT 63.927 96.104 64.175 96.184 ;
			LAYER M3 ;
			RECT 63.927 96.104 64.175 96.184 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[58]

	PIN D[59]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 97.736 64.175 97.816 ;
			LAYER M2 ;
			RECT 63.927 97.736 64.175 97.816 ;
			LAYER M3 ;
			RECT 63.927 97.736 64.175 97.816 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[59]

	PIN D[60]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 99.368 64.175 99.448 ;
			LAYER M2 ;
			RECT 63.927 99.368 64.175 99.448 ;
			LAYER M3 ;
			RECT 63.927 99.368 64.175 99.448 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[60]

	PIN D[61]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 101.000 64.175 101.080 ;
			LAYER M2 ;
			RECT 63.927 101.000 64.175 101.080 ;
			LAYER M3 ;
			RECT 63.927 101.000 64.175 101.080 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[61]

	PIN D[62]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 102.632 64.175 102.712 ;
			LAYER M2 ;
			RECT 63.927 102.632 64.175 102.712 ;
			LAYER M3 ;
			RECT 63.927 102.632 64.175 102.712 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[62]

	PIN D[63]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 104.264 64.175 104.344 ;
			LAYER M2 ;
			RECT 63.927 104.264 64.175 104.344 ;
			LAYER M3 ;
			RECT 63.927 104.264 64.175 104.344 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[63]

	PIN D[64]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 105.896 64.175 105.976 ;
			LAYER M2 ;
			RECT 63.927 105.896 64.175 105.976 ;
			LAYER M3 ;
			RECT 63.927 105.896 64.175 105.976 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[64]

	PIN D[65]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 107.528 64.175 107.608 ;
			LAYER M2 ;
			RECT 63.927 107.528 64.175 107.608 ;
			LAYER M3 ;
			RECT 63.927 107.528 64.175 107.608 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[65]

	PIN D[66]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 109.160 64.175 109.240 ;
			LAYER M2 ;
			RECT 63.927 109.160 64.175 109.240 ;
			LAYER M3 ;
			RECT 63.927 109.160 64.175 109.240 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[66]

	PIN D[67]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 110.792 64.175 110.872 ;
			LAYER M2 ;
			RECT 63.927 110.792 64.175 110.872 ;
			LAYER M3 ;
			RECT 63.927 110.792 64.175 110.872 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[67]

	PIN D[68]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 112.424 64.175 112.504 ;
			LAYER M2 ;
			RECT 63.927 112.424 64.175 112.504 ;
			LAYER M3 ;
			RECT 63.927 112.424 64.175 112.504 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[68]

	PIN D[69]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 114.056 64.175 114.136 ;
			LAYER M2 ;
			RECT 63.927 114.056 64.175 114.136 ;
			LAYER M3 ;
			RECT 63.927 114.056 64.175 114.136 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[69]

	PIN D[70]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 115.688 64.175 115.768 ;
			LAYER M2 ;
			RECT 63.927 115.688 64.175 115.768 ;
			LAYER M3 ;
			RECT 63.927 115.688 64.175 115.768 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[70]

	PIN D[71]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 117.320 64.175 117.400 ;
			LAYER M2 ;
			RECT 63.927 117.320 64.175 117.400 ;
			LAYER M3 ;
			RECT 63.927 117.320 64.175 117.400 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[71]

	PIN D[72]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 131.816 64.175 131.896 ;
			LAYER M2 ;
			RECT 63.927 131.816 64.175 131.896 ;
			LAYER M3 ;
			RECT 63.927 131.816 64.175 131.896 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[72]

	PIN D[73]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 133.448 64.175 133.528 ;
			LAYER M2 ;
			RECT 63.927 133.448 64.175 133.528 ;
			LAYER M3 ;
			RECT 63.927 133.448 64.175 133.528 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[73]

	PIN D[74]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 135.080 64.175 135.160 ;
			LAYER M2 ;
			RECT 63.927 135.080 64.175 135.160 ;
			LAYER M3 ;
			RECT 63.927 135.080 64.175 135.160 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[74]

	PIN D[75]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 136.712 64.175 136.792 ;
			LAYER M2 ;
			RECT 63.927 136.712 64.175 136.792 ;
			LAYER M3 ;
			RECT 63.927 136.712 64.175 136.792 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[75]

	PIN D[76]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 138.344 64.175 138.424 ;
			LAYER M2 ;
			RECT 63.927 138.344 64.175 138.424 ;
			LAYER M3 ;
			RECT 63.927 138.344 64.175 138.424 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[76]

	PIN D[77]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 139.976 64.175 140.056 ;
			LAYER M2 ;
			RECT 63.927 139.976 64.175 140.056 ;
			LAYER M3 ;
			RECT 63.927 139.976 64.175 140.056 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[77]

	PIN D[78]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 141.608 64.175 141.688 ;
			LAYER M2 ;
			RECT 63.927 141.608 64.175 141.688 ;
			LAYER M3 ;
			RECT 63.927 141.608 64.175 141.688 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[78]

	PIN D[79]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 143.240 64.175 143.320 ;
			LAYER M2 ;
			RECT 63.927 143.240 64.175 143.320 ;
			LAYER M3 ;
			RECT 63.927 143.240 64.175 143.320 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[79]

	PIN D[80]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 144.872 64.175 144.952 ;
			LAYER M2 ;
			RECT 63.927 144.872 64.175 144.952 ;
			LAYER M3 ;
			RECT 63.927 144.872 64.175 144.952 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[80]

	PIN D[81]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 146.504 64.175 146.584 ;
			LAYER M2 ;
			RECT 63.927 146.504 64.175 146.584 ;
			LAYER M3 ;
			RECT 63.927 146.504 64.175 146.584 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[81]

	PIN D[82]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 148.136 64.175 148.216 ;
			LAYER M2 ;
			RECT 63.927 148.136 64.175 148.216 ;
			LAYER M3 ;
			RECT 63.927 148.136 64.175 148.216 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[82]

	PIN D[83]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 149.768 64.175 149.848 ;
			LAYER M2 ;
			RECT 63.927 149.768 64.175 149.848 ;
			LAYER M3 ;
			RECT 63.927 149.768 64.175 149.848 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[83]

	PIN D[84]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 151.400 64.175 151.480 ;
			LAYER M2 ;
			RECT 63.927 151.400 64.175 151.480 ;
			LAYER M3 ;
			RECT 63.927 151.400 64.175 151.480 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[84]

	PIN D[85]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 153.032 64.175 153.112 ;
			LAYER M2 ;
			RECT 63.927 153.032 64.175 153.112 ;
			LAYER M3 ;
			RECT 63.927 153.032 64.175 153.112 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[85]

	PIN D[86]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 154.664 64.175 154.744 ;
			LAYER M2 ;
			RECT 63.927 154.664 64.175 154.744 ;
			LAYER M3 ;
			RECT 63.927 154.664 64.175 154.744 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[86]

	PIN D[87]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 156.296 64.175 156.376 ;
			LAYER M2 ;
			RECT 63.927 156.296 64.175 156.376 ;
			LAYER M3 ;
			RECT 63.927 156.296 64.175 156.376 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[87]

	PIN D[88]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 157.928 64.175 158.008 ;
			LAYER M2 ;
			RECT 63.927 157.928 64.175 158.008 ;
			LAYER M3 ;
			RECT 63.927 157.928 64.175 158.008 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[88]

	PIN D[89]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 159.560 64.175 159.640 ;
			LAYER M2 ;
			RECT 63.927 159.560 64.175 159.640 ;
			LAYER M3 ;
			RECT 63.927 159.560 64.175 159.640 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[89]

	PIN D[90]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 161.192 64.175 161.272 ;
			LAYER M2 ;
			RECT 63.927 161.192 64.175 161.272 ;
			LAYER M3 ;
			RECT 63.927 161.192 64.175 161.272 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[90]

	PIN D[91]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 162.824 64.175 162.904 ;
			LAYER M2 ;
			RECT 63.927 162.824 64.175 162.904 ;
			LAYER M3 ;
			RECT 63.927 162.824 64.175 162.904 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[91]

	PIN D[92]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 164.456 64.175 164.536 ;
			LAYER M2 ;
			RECT 63.927 164.456 64.175 164.536 ;
			LAYER M3 ;
			RECT 63.927 164.456 64.175 164.536 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[92]

	PIN D[93]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 166.088 64.175 166.168 ;
			LAYER M2 ;
			RECT 63.927 166.088 64.175 166.168 ;
			LAYER M3 ;
			RECT 63.927 166.088 64.175 166.168 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[93]

	PIN D[94]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 167.720 64.175 167.800 ;
			LAYER M2 ;
			RECT 63.927 167.720 64.175 167.800 ;
			LAYER M3 ;
			RECT 63.927 167.720 64.175 167.800 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[94]

	PIN D[95]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 169.352 64.175 169.432 ;
			LAYER M2 ;
			RECT 63.927 169.352 64.175 169.432 ;
			LAYER M3 ;
			RECT 63.927 169.352 64.175 169.432 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[95]

	PIN D[96]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 170.984 64.175 171.064 ;
			LAYER M2 ;
			RECT 63.927 170.984 64.175 171.064 ;
			LAYER M3 ;
			RECT 63.927 170.984 64.175 171.064 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[96]

	PIN D[97]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 172.616 64.175 172.696 ;
			LAYER M2 ;
			RECT 63.927 172.616 64.175 172.696 ;
			LAYER M3 ;
			RECT 63.927 172.616 64.175 172.696 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[97]

	PIN D[98]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 174.248 64.175 174.328 ;
			LAYER M2 ;
			RECT 63.927 174.248 64.175 174.328 ;
			LAYER M3 ;
			RECT 63.927 174.248 64.175 174.328 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[98]

	PIN D[99]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 175.880 64.175 175.960 ;
			LAYER M2 ;
			RECT 63.927 175.880 64.175 175.960 ;
			LAYER M3 ;
			RECT 63.927 175.880 64.175 175.960 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[99]

	PIN D[100]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 177.512 64.175 177.592 ;
			LAYER M2 ;
			RECT 63.927 177.512 64.175 177.592 ;
			LAYER M3 ;
			RECT 63.927 177.512 64.175 177.592 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[100]

	PIN D[101]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 179.144 64.175 179.224 ;
			LAYER M2 ;
			RECT 63.927 179.144 64.175 179.224 ;
			LAYER M3 ;
			RECT 63.927 179.144 64.175 179.224 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[101]

	PIN D[102]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 180.776 64.175 180.856 ;
			LAYER M2 ;
			RECT 63.927 180.776 64.175 180.856 ;
			LAYER M3 ;
			RECT 63.927 180.776 64.175 180.856 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[102]

	PIN D[103]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 182.408 64.175 182.488 ;
			LAYER M2 ;
			RECT 63.927 182.408 64.175 182.488 ;
			LAYER M3 ;
			RECT 63.927 182.408 64.175 182.488 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[103]

	PIN D[104]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 184.040 64.175 184.120 ;
			LAYER M2 ;
			RECT 63.927 184.040 64.175 184.120 ;
			LAYER M3 ;
			RECT 63.927 184.040 64.175 184.120 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[104]

	PIN D[105]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 185.672 64.175 185.752 ;
			LAYER M2 ;
			RECT 63.927 185.672 64.175 185.752 ;
			LAYER M3 ;
			RECT 63.927 185.672 64.175 185.752 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[105]

	PIN D[106]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 187.304 64.175 187.384 ;
			LAYER M2 ;
			RECT 63.927 187.304 64.175 187.384 ;
			LAYER M3 ;
			RECT 63.927 187.304 64.175 187.384 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[106]

	PIN D[107]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 188.936 64.175 189.016 ;
			LAYER M2 ;
			RECT 63.927 188.936 64.175 189.016 ;
			LAYER M3 ;
			RECT 63.927 188.936 64.175 189.016 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[107]

	PIN D[108]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 190.568 64.175 190.648 ;
			LAYER M2 ;
			RECT 63.927 190.568 64.175 190.648 ;
			LAYER M3 ;
			RECT 63.927 190.568 64.175 190.648 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[108]

	PIN D[109]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 192.200 64.175 192.280 ;
			LAYER M2 ;
			RECT 63.927 192.200 64.175 192.280 ;
			LAYER M3 ;
			RECT 63.927 192.200 64.175 192.280 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[109]

	PIN D[110]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 193.832 64.175 193.912 ;
			LAYER M2 ;
			RECT 63.927 193.832 64.175 193.912 ;
			LAYER M3 ;
			RECT 63.927 193.832 64.175 193.912 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[110]

	PIN D[111]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 195.464 64.175 195.544 ;
			LAYER M2 ;
			RECT 63.927 195.464 64.175 195.544 ;
			LAYER M3 ;
			RECT 63.927 195.464 64.175 195.544 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[111]

	PIN D[112]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 197.096 64.175 197.176 ;
			LAYER M2 ;
			RECT 63.927 197.096 64.175 197.176 ;
			LAYER M3 ;
			RECT 63.927 197.096 64.175 197.176 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[112]

	PIN D[113]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 198.728 64.175 198.808 ;
			LAYER M2 ;
			RECT 63.927 198.728 64.175 198.808 ;
			LAYER M3 ;
			RECT 63.927 198.728 64.175 198.808 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[113]

	PIN D[114]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 200.360 64.175 200.440 ;
			LAYER M2 ;
			RECT 63.927 200.360 64.175 200.440 ;
			LAYER M3 ;
			RECT 63.927 200.360 64.175 200.440 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[114]

	PIN D[115]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 201.992 64.175 202.072 ;
			LAYER M2 ;
			RECT 63.927 201.992 64.175 202.072 ;
			LAYER M3 ;
			RECT 63.927 201.992 64.175 202.072 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[115]

	PIN D[116]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 203.624 64.175 203.704 ;
			LAYER M2 ;
			RECT 63.927 203.624 64.175 203.704 ;
			LAYER M3 ;
			RECT 63.927 203.624 64.175 203.704 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[116]

	PIN D[117]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 205.256 64.175 205.336 ;
			LAYER M2 ;
			RECT 63.927 205.256 64.175 205.336 ;
			LAYER M3 ;
			RECT 63.927 205.256 64.175 205.336 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[117]

	PIN D[118]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 206.888 64.175 206.968 ;
			LAYER M2 ;
			RECT 63.927 206.888 64.175 206.968 ;
			LAYER M3 ;
			RECT 63.927 206.888 64.175 206.968 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[118]

	PIN D[119]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 208.520 64.175 208.600 ;
			LAYER M2 ;
			RECT 63.927 208.520 64.175 208.600 ;
			LAYER M3 ;
			RECT 63.927 208.520 64.175 208.600 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[119]

	PIN D[120]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 210.152 64.175 210.232 ;
			LAYER M2 ;
			RECT 63.927 210.152 64.175 210.232 ;
			LAYER M3 ;
			RECT 63.927 210.152 64.175 210.232 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[120]

	PIN D[121]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 211.784 64.175 211.864 ;
			LAYER M2 ;
			RECT 63.927 211.784 64.175 211.864 ;
			LAYER M3 ;
			RECT 63.927 211.784 64.175 211.864 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[121]

	PIN D[122]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 213.416 64.175 213.496 ;
			LAYER M2 ;
			RECT 63.927 213.416 64.175 213.496 ;
			LAYER M3 ;
			RECT 63.927 213.416 64.175 213.496 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[122]

	PIN D[123]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 215.048 64.175 215.128 ;
			LAYER M2 ;
			RECT 63.927 215.048 64.175 215.128 ;
			LAYER M3 ;
			RECT 63.927 215.048 64.175 215.128 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[123]

	PIN D[124]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 216.680 64.175 216.760 ;
			LAYER M2 ;
			RECT 63.927 216.680 64.175 216.760 ;
			LAYER M3 ;
			RECT 63.927 216.680 64.175 216.760 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[124]

	PIN D[125]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 218.312 64.175 218.392 ;
			LAYER M2 ;
			RECT 63.927 218.312 64.175 218.392 ;
			LAYER M3 ;
			RECT 63.927 218.312 64.175 218.392 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[125]

	PIN D[126]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 219.944 64.175 220.024 ;
			LAYER M2 ;
			RECT 63.927 219.944 64.175 220.024 ;
			LAYER M3 ;
			RECT 63.927 219.944 64.175 220.024 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[126]

	PIN D[127]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 221.576 64.175 221.656 ;
			LAYER M2 ;
			RECT 63.927 221.576 64.175 221.656 ;
			LAYER M3 ;
			RECT 63.927 221.576 64.175 221.656 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[127]

	PIN D[128]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 223.208 64.175 223.288 ;
			LAYER M2 ;
			RECT 63.927 223.208 64.175 223.288 ;
			LAYER M3 ;
			RECT 63.927 223.208 64.175 223.288 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[128]

	PIN D[129]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 224.840 64.175 224.920 ;
			LAYER M2 ;
			RECT 63.927 224.840 64.175 224.920 ;
			LAYER M3 ;
			RECT 63.927 224.840 64.175 224.920 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[129]

	PIN D[130]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 226.472 64.175 226.552 ;
			LAYER M2 ;
			RECT 63.927 226.472 64.175 226.552 ;
			LAYER M3 ;
			RECT 63.927 226.472 64.175 226.552 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[130]

	PIN D[131]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 228.104 64.175 228.184 ;
			LAYER M2 ;
			RECT 63.927 228.104 64.175 228.184 ;
			LAYER M3 ;
			RECT 63.927 228.104 64.175 228.184 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[131]

	PIN D[132]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 229.736 64.175 229.816 ;
			LAYER M2 ;
			RECT 63.927 229.736 64.175 229.816 ;
			LAYER M3 ;
			RECT 63.927 229.736 64.175 229.816 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[132]

	PIN D[133]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 231.368 64.175 231.448 ;
			LAYER M2 ;
			RECT 63.927 231.368 64.175 231.448 ;
			LAYER M3 ;
			RECT 63.927 231.368 64.175 231.448 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[133]

	PIN D[134]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 233.000 64.175 233.080 ;
			LAYER M2 ;
			RECT 63.927 233.000 64.175 233.080 ;
			LAYER M3 ;
			RECT 63.927 233.000 64.175 233.080 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[134]

	PIN D[135]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 234.632 64.175 234.712 ;
			LAYER M2 ;
			RECT 63.927 234.632 64.175 234.712 ;
			LAYER M3 ;
			RECT 63.927 234.632 64.175 234.712 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[135]

	PIN D[136]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 236.264 64.175 236.344 ;
			LAYER M2 ;
			RECT 63.927 236.264 64.175 236.344 ;
			LAYER M3 ;
			RECT 63.927 236.264 64.175 236.344 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[136]

	PIN D[137]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 237.896 64.175 237.976 ;
			LAYER M2 ;
			RECT 63.927 237.896 64.175 237.976 ;
			LAYER M3 ;
			RECT 63.927 237.896 64.175 237.976 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[137]

	PIN D[138]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 239.528 64.175 239.608 ;
			LAYER M2 ;
			RECT 63.927 239.528 64.175 239.608 ;
			LAYER M3 ;
			RECT 63.927 239.528 64.175 239.608 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[138]

	PIN D[139]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 241.160 64.175 241.240 ;
			LAYER M2 ;
			RECT 63.927 241.160 64.175 241.240 ;
			LAYER M3 ;
			RECT 63.927 241.160 64.175 241.240 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[139]

	PIN D[140]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 242.792 64.175 242.872 ;
			LAYER M2 ;
			RECT 63.927 242.792 64.175 242.872 ;
			LAYER M3 ;
			RECT 63.927 242.792 64.175 242.872 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[140]

	PIN D[141]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 244.424 64.175 244.504 ;
			LAYER M2 ;
			RECT 63.927 244.424 64.175 244.504 ;
			LAYER M3 ;
			RECT 63.927 244.424 64.175 244.504 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[141]

	PIN D[142]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 246.056 64.175 246.136 ;
			LAYER M2 ;
			RECT 63.927 246.056 64.175 246.136 ;
			LAYER M3 ;
			RECT 63.927 246.056 64.175 246.136 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[142]

	PIN D[143]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 247.688 64.175 247.768 ;
			LAYER M2 ;
			RECT 63.927 247.688 64.175 247.768 ;
			LAYER M3 ;
			RECT 63.927 247.688 64.175 247.768 ;
		END
		ANTENNAGATEAREA 0.001840 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100920 LAYER M1 ;
		ANTENNAMAXAREACAR 15.881400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001840 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.174240 LAYER M2 ;
		ANTENNAMAXAREACAR 37.580600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001840 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121320 LAYER M3 ;
		ANTENNAMAXAREACAR 89.873800 LAYER M3 ;
	END D[143]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 1.784 64.175 1.864 ;
			LAYER M2 ;
			RECT 63.927 1.784 64.175 1.864 ;
			LAYER M3 ;
			RECT 63.927 1.784 64.175 1.864 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[0]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 3.416 64.175 3.496 ;
			LAYER M2 ;
			RECT 63.927 3.416 64.175 3.496 ;
			LAYER M3 ;
			RECT 63.927 3.416 64.175 3.496 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[1]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 5.048 64.175 5.128 ;
			LAYER M2 ;
			RECT 63.927 5.048 64.175 5.128 ;
			LAYER M3 ;
			RECT 63.927 5.048 64.175 5.128 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[2]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 6.680 64.175 6.760 ;
			LAYER M2 ;
			RECT 63.927 6.680 64.175 6.760 ;
			LAYER M3 ;
			RECT 63.927 6.680 64.175 6.760 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[3]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 8.312 64.175 8.392 ;
			LAYER M2 ;
			RECT 63.927 8.312 64.175 8.392 ;
			LAYER M3 ;
			RECT 63.927 8.312 64.175 8.392 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[4]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 9.944 64.175 10.024 ;
			LAYER M2 ;
			RECT 63.927 9.944 64.175 10.024 ;
			LAYER M3 ;
			RECT 63.927 9.944 64.175 10.024 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[5]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 11.576 64.175 11.656 ;
			LAYER M2 ;
			RECT 63.927 11.576 64.175 11.656 ;
			LAYER M3 ;
			RECT 63.927 11.576 64.175 11.656 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 13.208 64.175 13.288 ;
			LAYER M2 ;
			RECT 63.927 13.208 64.175 13.288 ;
			LAYER M3 ;
			RECT 63.927 13.208 64.175 13.288 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[7]

	PIN Q[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 14.840 64.175 14.920 ;
			LAYER M2 ;
			RECT 63.927 14.840 64.175 14.920 ;
			LAYER M3 ;
			RECT 63.927 14.840 64.175 14.920 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[8]

	PIN Q[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 16.472 64.175 16.552 ;
			LAYER M2 ;
			RECT 63.927 16.472 64.175 16.552 ;
			LAYER M3 ;
			RECT 63.927 16.472 64.175 16.552 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[9]

	PIN Q[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 18.104 64.175 18.184 ;
			LAYER M2 ;
			RECT 63.927 18.104 64.175 18.184 ;
			LAYER M3 ;
			RECT 63.927 18.104 64.175 18.184 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[10]

	PIN Q[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 19.736 64.175 19.816 ;
			LAYER M2 ;
			RECT 63.927 19.736 64.175 19.816 ;
			LAYER M3 ;
			RECT 63.927 19.736 64.175 19.816 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[11]

	PIN Q[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 21.368 64.175 21.448 ;
			LAYER M2 ;
			RECT 63.927 21.368 64.175 21.448 ;
			LAYER M3 ;
			RECT 63.927 21.368 64.175 21.448 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[12]

	PIN Q[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 23.000 64.175 23.080 ;
			LAYER M2 ;
			RECT 63.927 23.000 64.175 23.080 ;
			LAYER M3 ;
			RECT 63.927 23.000 64.175 23.080 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[13]

	PIN Q[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 24.632 64.175 24.712 ;
			LAYER M2 ;
			RECT 63.927 24.632 64.175 24.712 ;
			LAYER M3 ;
			RECT 63.927 24.632 64.175 24.712 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[14]

	PIN Q[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 26.264 64.175 26.344 ;
			LAYER M2 ;
			RECT 63.927 26.264 64.175 26.344 ;
			LAYER M3 ;
			RECT 63.927 26.264 64.175 26.344 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[15]

	PIN Q[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 27.896 64.175 27.976 ;
			LAYER M2 ;
			RECT 63.927 27.896 64.175 27.976 ;
			LAYER M3 ;
			RECT 63.927 27.896 64.175 27.976 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[16]

	PIN Q[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 29.528 64.175 29.608 ;
			LAYER M2 ;
			RECT 63.927 29.528 64.175 29.608 ;
			LAYER M3 ;
			RECT 63.927 29.528 64.175 29.608 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[17]

	PIN Q[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 31.160 64.175 31.240 ;
			LAYER M2 ;
			RECT 63.927 31.160 64.175 31.240 ;
			LAYER M3 ;
			RECT 63.927 31.160 64.175 31.240 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[18]

	PIN Q[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 32.792 64.175 32.872 ;
			LAYER M2 ;
			RECT 63.927 32.792 64.175 32.872 ;
			LAYER M3 ;
			RECT 63.927 32.792 64.175 32.872 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[19]

	PIN Q[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 34.424 64.175 34.504 ;
			LAYER M2 ;
			RECT 63.927 34.424 64.175 34.504 ;
			LAYER M3 ;
			RECT 63.927 34.424 64.175 34.504 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[20]

	PIN Q[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 36.056 64.175 36.136 ;
			LAYER M2 ;
			RECT 63.927 36.056 64.175 36.136 ;
			LAYER M3 ;
			RECT 63.927 36.056 64.175 36.136 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[21]

	PIN Q[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 37.688 64.175 37.768 ;
			LAYER M2 ;
			RECT 63.927 37.688 64.175 37.768 ;
			LAYER M3 ;
			RECT 63.927 37.688 64.175 37.768 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[22]

	PIN Q[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 39.320 64.175 39.400 ;
			LAYER M2 ;
			RECT 63.927 39.320 64.175 39.400 ;
			LAYER M3 ;
			RECT 63.927 39.320 64.175 39.400 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[23]

	PIN Q[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 40.952 64.175 41.032 ;
			LAYER M2 ;
			RECT 63.927 40.952 64.175 41.032 ;
			LAYER M3 ;
			RECT 63.927 40.952 64.175 41.032 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[24]

	PIN Q[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 42.584 64.175 42.664 ;
			LAYER M2 ;
			RECT 63.927 42.584 64.175 42.664 ;
			LAYER M3 ;
			RECT 63.927 42.584 64.175 42.664 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[25]

	PIN Q[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 44.216 64.175 44.296 ;
			LAYER M2 ;
			RECT 63.927 44.216 64.175 44.296 ;
			LAYER M3 ;
			RECT 63.927 44.216 64.175 44.296 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[26]

	PIN Q[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 45.848 64.175 45.928 ;
			LAYER M2 ;
			RECT 63.927 45.848 64.175 45.928 ;
			LAYER M3 ;
			RECT 63.927 45.848 64.175 45.928 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[27]

	PIN Q[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 47.480 64.175 47.560 ;
			LAYER M2 ;
			RECT 63.927 47.480 64.175 47.560 ;
			LAYER M3 ;
			RECT 63.927 47.480 64.175 47.560 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[28]

	PIN Q[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 49.112 64.175 49.192 ;
			LAYER M2 ;
			RECT 63.927 49.112 64.175 49.192 ;
			LAYER M3 ;
			RECT 63.927 49.112 64.175 49.192 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[29]

	PIN Q[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 50.744 64.175 50.824 ;
			LAYER M2 ;
			RECT 63.927 50.744 64.175 50.824 ;
			LAYER M3 ;
			RECT 63.927 50.744 64.175 50.824 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[30]

	PIN Q[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 52.376 64.175 52.456 ;
			LAYER M2 ;
			RECT 63.927 52.376 64.175 52.456 ;
			LAYER M3 ;
			RECT 63.927 52.376 64.175 52.456 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[31]

	PIN Q[32]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 54.008 64.175 54.088 ;
			LAYER M2 ;
			RECT 63.927 54.008 64.175 54.088 ;
			LAYER M3 ;
			RECT 63.927 54.008 64.175 54.088 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[32]

	PIN Q[33]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 55.640 64.175 55.720 ;
			LAYER M2 ;
			RECT 63.927 55.640 64.175 55.720 ;
			LAYER M3 ;
			RECT 63.927 55.640 64.175 55.720 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[33]

	PIN Q[34]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 57.272 64.175 57.352 ;
			LAYER M2 ;
			RECT 63.927 57.272 64.175 57.352 ;
			LAYER M3 ;
			RECT 63.927 57.272 64.175 57.352 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[34]

	PIN Q[35]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 58.904 64.175 58.984 ;
			LAYER M2 ;
			RECT 63.927 58.904 64.175 58.984 ;
			LAYER M3 ;
			RECT 63.927 58.904 64.175 58.984 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[35]

	PIN Q[36]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 60.536 64.175 60.616 ;
			LAYER M2 ;
			RECT 63.927 60.536 64.175 60.616 ;
			LAYER M3 ;
			RECT 63.927 60.536 64.175 60.616 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[36]

	PIN Q[37]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 62.168 64.175 62.248 ;
			LAYER M2 ;
			RECT 63.927 62.168 64.175 62.248 ;
			LAYER M3 ;
			RECT 63.927 62.168 64.175 62.248 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[37]

	PIN Q[38]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 63.800 64.175 63.880 ;
			LAYER M2 ;
			RECT 63.927 63.800 64.175 63.880 ;
			LAYER M3 ;
			RECT 63.927 63.800 64.175 63.880 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[38]

	PIN Q[39]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 65.432 64.175 65.512 ;
			LAYER M2 ;
			RECT 63.927 65.432 64.175 65.512 ;
			LAYER M3 ;
			RECT 63.927 65.432 64.175 65.512 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[39]

	PIN Q[40]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 67.064 64.175 67.144 ;
			LAYER M2 ;
			RECT 63.927 67.064 64.175 67.144 ;
			LAYER M3 ;
			RECT 63.927 67.064 64.175 67.144 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[40]

	PIN Q[41]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 68.696 64.175 68.776 ;
			LAYER M2 ;
			RECT 63.927 68.696 64.175 68.776 ;
			LAYER M3 ;
			RECT 63.927 68.696 64.175 68.776 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[41]

	PIN Q[42]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 70.328 64.175 70.408 ;
			LAYER M2 ;
			RECT 63.927 70.328 64.175 70.408 ;
			LAYER M3 ;
			RECT 63.927 70.328 64.175 70.408 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[42]

	PIN Q[43]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 71.960 64.175 72.040 ;
			LAYER M2 ;
			RECT 63.927 71.960 64.175 72.040 ;
			LAYER M3 ;
			RECT 63.927 71.960 64.175 72.040 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[43]

	PIN Q[44]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 73.592 64.175 73.672 ;
			LAYER M2 ;
			RECT 63.927 73.592 64.175 73.672 ;
			LAYER M3 ;
			RECT 63.927 73.592 64.175 73.672 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[44]

	PIN Q[45]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 75.224 64.175 75.304 ;
			LAYER M2 ;
			RECT 63.927 75.224 64.175 75.304 ;
			LAYER M3 ;
			RECT 63.927 75.224 64.175 75.304 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[45]

	PIN Q[46]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 76.856 64.175 76.936 ;
			LAYER M2 ;
			RECT 63.927 76.856 64.175 76.936 ;
			LAYER M3 ;
			RECT 63.927 76.856 64.175 76.936 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[46]

	PIN Q[47]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 78.488 64.175 78.568 ;
			LAYER M2 ;
			RECT 63.927 78.488 64.175 78.568 ;
			LAYER M3 ;
			RECT 63.927 78.488 64.175 78.568 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[47]

	PIN Q[48]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 80.120 64.175 80.200 ;
			LAYER M2 ;
			RECT 63.927 80.120 64.175 80.200 ;
			LAYER M3 ;
			RECT 63.927 80.120 64.175 80.200 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[48]

	PIN Q[49]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 81.752 64.175 81.832 ;
			LAYER M2 ;
			RECT 63.927 81.752 64.175 81.832 ;
			LAYER M3 ;
			RECT 63.927 81.752 64.175 81.832 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[49]

	PIN Q[50]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 83.384 64.175 83.464 ;
			LAYER M2 ;
			RECT 63.927 83.384 64.175 83.464 ;
			LAYER M3 ;
			RECT 63.927 83.384 64.175 83.464 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[50]

	PIN Q[51]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 85.016 64.175 85.096 ;
			LAYER M2 ;
			RECT 63.927 85.016 64.175 85.096 ;
			LAYER M3 ;
			RECT 63.927 85.016 64.175 85.096 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[51]

	PIN Q[52]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 86.648 64.175 86.728 ;
			LAYER M2 ;
			RECT 63.927 86.648 64.175 86.728 ;
			LAYER M3 ;
			RECT 63.927 86.648 64.175 86.728 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[52]

	PIN Q[53]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 88.280 64.175 88.360 ;
			LAYER M2 ;
			RECT 63.927 88.280 64.175 88.360 ;
			LAYER M3 ;
			RECT 63.927 88.280 64.175 88.360 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[53]

	PIN Q[54]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 89.912 64.175 89.992 ;
			LAYER M2 ;
			RECT 63.927 89.912 64.175 89.992 ;
			LAYER M3 ;
			RECT 63.927 89.912 64.175 89.992 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[54]

	PIN Q[55]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 91.544 64.175 91.624 ;
			LAYER M2 ;
			RECT 63.927 91.544 64.175 91.624 ;
			LAYER M3 ;
			RECT 63.927 91.544 64.175 91.624 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[55]

	PIN Q[56]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 93.176 64.175 93.256 ;
			LAYER M2 ;
			RECT 63.927 93.176 64.175 93.256 ;
			LAYER M3 ;
			RECT 63.927 93.176 64.175 93.256 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[56]

	PIN Q[57]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 94.808 64.175 94.888 ;
			LAYER M2 ;
			RECT 63.927 94.808 64.175 94.888 ;
			LAYER M3 ;
			RECT 63.927 94.808 64.175 94.888 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[57]

	PIN Q[58]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 96.440 64.175 96.520 ;
			LAYER M2 ;
			RECT 63.927 96.440 64.175 96.520 ;
			LAYER M3 ;
			RECT 63.927 96.440 64.175 96.520 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[58]

	PIN Q[59]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 98.072 64.175 98.152 ;
			LAYER M2 ;
			RECT 63.927 98.072 64.175 98.152 ;
			LAYER M3 ;
			RECT 63.927 98.072 64.175 98.152 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[59]

	PIN Q[60]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 99.704 64.175 99.784 ;
			LAYER M2 ;
			RECT 63.927 99.704 64.175 99.784 ;
			LAYER M3 ;
			RECT 63.927 99.704 64.175 99.784 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[60]

	PIN Q[61]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 101.336 64.175 101.416 ;
			LAYER M2 ;
			RECT 63.927 101.336 64.175 101.416 ;
			LAYER M3 ;
			RECT 63.927 101.336 64.175 101.416 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[61]

	PIN Q[62]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 102.968 64.175 103.048 ;
			LAYER M2 ;
			RECT 63.927 102.968 64.175 103.048 ;
			LAYER M3 ;
			RECT 63.927 102.968 64.175 103.048 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[62]

	PIN Q[63]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 104.600 64.175 104.680 ;
			LAYER M2 ;
			RECT 63.927 104.600 64.175 104.680 ;
			LAYER M3 ;
			RECT 63.927 104.600 64.175 104.680 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[63]

	PIN Q[64]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 106.232 64.175 106.312 ;
			LAYER M2 ;
			RECT 63.927 106.232 64.175 106.312 ;
			LAYER M3 ;
			RECT 63.927 106.232 64.175 106.312 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[64]

	PIN Q[65]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 107.864 64.175 107.944 ;
			LAYER M2 ;
			RECT 63.927 107.864 64.175 107.944 ;
			LAYER M3 ;
			RECT 63.927 107.864 64.175 107.944 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[65]

	PIN Q[66]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 109.496 64.175 109.576 ;
			LAYER M2 ;
			RECT 63.927 109.496 64.175 109.576 ;
			LAYER M3 ;
			RECT 63.927 109.496 64.175 109.576 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[66]

	PIN Q[67]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 111.128 64.175 111.208 ;
			LAYER M2 ;
			RECT 63.927 111.128 64.175 111.208 ;
			LAYER M3 ;
			RECT 63.927 111.128 64.175 111.208 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[67]

	PIN Q[68]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 112.760 64.175 112.840 ;
			LAYER M2 ;
			RECT 63.927 112.760 64.175 112.840 ;
			LAYER M3 ;
			RECT 63.927 112.760 64.175 112.840 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[68]

	PIN Q[69]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 114.392 64.175 114.472 ;
			LAYER M2 ;
			RECT 63.927 114.392 64.175 114.472 ;
			LAYER M3 ;
			RECT 63.927 114.392 64.175 114.472 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[69]

	PIN Q[70]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 116.024 64.175 116.104 ;
			LAYER M2 ;
			RECT 63.927 116.024 64.175 116.104 ;
			LAYER M3 ;
			RECT 63.927 116.024 64.175 116.104 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[70]

	PIN Q[71]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 117.656 64.175 117.736 ;
			LAYER M2 ;
			RECT 63.927 117.656 64.175 117.736 ;
			LAYER M3 ;
			RECT 63.927 117.656 64.175 117.736 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[71]

	PIN Q[72]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 132.152 64.175 132.232 ;
			LAYER M2 ;
			RECT 63.927 132.152 64.175 132.232 ;
			LAYER M3 ;
			RECT 63.927 132.152 64.175 132.232 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[72]

	PIN Q[73]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 133.784 64.175 133.864 ;
			LAYER M2 ;
			RECT 63.927 133.784 64.175 133.864 ;
			LAYER M3 ;
			RECT 63.927 133.784 64.175 133.864 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[73]

	PIN Q[74]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 135.416 64.175 135.496 ;
			LAYER M2 ;
			RECT 63.927 135.416 64.175 135.496 ;
			LAYER M3 ;
			RECT 63.927 135.416 64.175 135.496 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[74]

	PIN Q[75]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 137.048 64.175 137.128 ;
			LAYER M2 ;
			RECT 63.927 137.048 64.175 137.128 ;
			LAYER M3 ;
			RECT 63.927 137.048 64.175 137.128 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[75]

	PIN Q[76]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 138.680 64.175 138.760 ;
			LAYER M2 ;
			RECT 63.927 138.680 64.175 138.760 ;
			LAYER M3 ;
			RECT 63.927 138.680 64.175 138.760 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[76]

	PIN Q[77]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 140.312 64.175 140.392 ;
			LAYER M2 ;
			RECT 63.927 140.312 64.175 140.392 ;
			LAYER M3 ;
			RECT 63.927 140.312 64.175 140.392 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[77]

	PIN Q[78]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 141.944 64.175 142.024 ;
			LAYER M2 ;
			RECT 63.927 141.944 64.175 142.024 ;
			LAYER M3 ;
			RECT 63.927 141.944 64.175 142.024 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[78]

	PIN Q[79]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 143.576 64.175 143.656 ;
			LAYER M2 ;
			RECT 63.927 143.576 64.175 143.656 ;
			LAYER M3 ;
			RECT 63.927 143.576 64.175 143.656 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[79]

	PIN Q[80]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 145.208 64.175 145.288 ;
			LAYER M2 ;
			RECT 63.927 145.208 64.175 145.288 ;
			LAYER M3 ;
			RECT 63.927 145.208 64.175 145.288 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[80]

	PIN Q[81]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 146.840 64.175 146.920 ;
			LAYER M2 ;
			RECT 63.927 146.840 64.175 146.920 ;
			LAYER M3 ;
			RECT 63.927 146.840 64.175 146.920 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[81]

	PIN Q[82]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 148.472 64.175 148.552 ;
			LAYER M2 ;
			RECT 63.927 148.472 64.175 148.552 ;
			LAYER M3 ;
			RECT 63.927 148.472 64.175 148.552 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[82]

	PIN Q[83]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 150.104 64.175 150.184 ;
			LAYER M2 ;
			RECT 63.927 150.104 64.175 150.184 ;
			LAYER M3 ;
			RECT 63.927 150.104 64.175 150.184 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[83]

	PIN Q[84]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 151.736 64.175 151.816 ;
			LAYER M2 ;
			RECT 63.927 151.736 64.175 151.816 ;
			LAYER M3 ;
			RECT 63.927 151.736 64.175 151.816 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[84]

	PIN Q[85]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 153.368 64.175 153.448 ;
			LAYER M2 ;
			RECT 63.927 153.368 64.175 153.448 ;
			LAYER M3 ;
			RECT 63.927 153.368 64.175 153.448 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[85]

	PIN Q[86]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 155.000 64.175 155.080 ;
			LAYER M2 ;
			RECT 63.927 155.000 64.175 155.080 ;
			LAYER M3 ;
			RECT 63.927 155.000 64.175 155.080 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[86]

	PIN Q[87]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 156.632 64.175 156.712 ;
			LAYER M2 ;
			RECT 63.927 156.632 64.175 156.712 ;
			LAYER M3 ;
			RECT 63.927 156.632 64.175 156.712 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[87]

	PIN Q[88]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 158.264 64.175 158.344 ;
			LAYER M2 ;
			RECT 63.927 158.264 64.175 158.344 ;
			LAYER M3 ;
			RECT 63.927 158.264 64.175 158.344 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[88]

	PIN Q[89]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 159.896 64.175 159.976 ;
			LAYER M2 ;
			RECT 63.927 159.896 64.175 159.976 ;
			LAYER M3 ;
			RECT 63.927 159.896 64.175 159.976 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[89]

	PIN Q[90]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 161.528 64.175 161.608 ;
			LAYER M2 ;
			RECT 63.927 161.528 64.175 161.608 ;
			LAYER M3 ;
			RECT 63.927 161.528 64.175 161.608 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[90]

	PIN Q[91]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 163.160 64.175 163.240 ;
			LAYER M2 ;
			RECT 63.927 163.160 64.175 163.240 ;
			LAYER M3 ;
			RECT 63.927 163.160 64.175 163.240 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[91]

	PIN Q[92]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 164.792 64.175 164.872 ;
			LAYER M2 ;
			RECT 63.927 164.792 64.175 164.872 ;
			LAYER M3 ;
			RECT 63.927 164.792 64.175 164.872 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[92]

	PIN Q[93]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 166.424 64.175 166.504 ;
			LAYER M2 ;
			RECT 63.927 166.424 64.175 166.504 ;
			LAYER M3 ;
			RECT 63.927 166.424 64.175 166.504 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[93]

	PIN Q[94]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 168.056 64.175 168.136 ;
			LAYER M2 ;
			RECT 63.927 168.056 64.175 168.136 ;
			LAYER M3 ;
			RECT 63.927 168.056 64.175 168.136 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[94]

	PIN Q[95]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 169.688 64.175 169.768 ;
			LAYER M2 ;
			RECT 63.927 169.688 64.175 169.768 ;
			LAYER M3 ;
			RECT 63.927 169.688 64.175 169.768 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[95]

	PIN Q[96]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 171.320 64.175 171.400 ;
			LAYER M2 ;
			RECT 63.927 171.320 64.175 171.400 ;
			LAYER M3 ;
			RECT 63.927 171.320 64.175 171.400 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[96]

	PIN Q[97]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 172.952 64.175 173.032 ;
			LAYER M2 ;
			RECT 63.927 172.952 64.175 173.032 ;
			LAYER M3 ;
			RECT 63.927 172.952 64.175 173.032 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[97]

	PIN Q[98]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 174.584 64.175 174.664 ;
			LAYER M2 ;
			RECT 63.927 174.584 64.175 174.664 ;
			LAYER M3 ;
			RECT 63.927 174.584 64.175 174.664 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[98]

	PIN Q[99]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 176.216 64.175 176.296 ;
			LAYER M2 ;
			RECT 63.927 176.216 64.175 176.296 ;
			LAYER M3 ;
			RECT 63.927 176.216 64.175 176.296 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[99]

	PIN Q[100]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 177.848 64.175 177.928 ;
			LAYER M2 ;
			RECT 63.927 177.848 64.175 177.928 ;
			LAYER M3 ;
			RECT 63.927 177.848 64.175 177.928 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[100]

	PIN Q[101]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 179.480 64.175 179.560 ;
			LAYER M2 ;
			RECT 63.927 179.480 64.175 179.560 ;
			LAYER M3 ;
			RECT 63.927 179.480 64.175 179.560 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[101]

	PIN Q[102]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 181.112 64.175 181.192 ;
			LAYER M2 ;
			RECT 63.927 181.112 64.175 181.192 ;
			LAYER M3 ;
			RECT 63.927 181.112 64.175 181.192 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[102]

	PIN Q[103]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 182.744 64.175 182.824 ;
			LAYER M2 ;
			RECT 63.927 182.744 64.175 182.824 ;
			LAYER M3 ;
			RECT 63.927 182.744 64.175 182.824 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[103]

	PIN Q[104]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 184.376 64.175 184.456 ;
			LAYER M2 ;
			RECT 63.927 184.376 64.175 184.456 ;
			LAYER M3 ;
			RECT 63.927 184.376 64.175 184.456 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[104]

	PIN Q[105]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 186.008 64.175 186.088 ;
			LAYER M2 ;
			RECT 63.927 186.008 64.175 186.088 ;
			LAYER M3 ;
			RECT 63.927 186.008 64.175 186.088 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[105]

	PIN Q[106]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 187.640 64.175 187.720 ;
			LAYER M2 ;
			RECT 63.927 187.640 64.175 187.720 ;
			LAYER M3 ;
			RECT 63.927 187.640 64.175 187.720 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[106]

	PIN Q[107]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 189.272 64.175 189.352 ;
			LAYER M2 ;
			RECT 63.927 189.272 64.175 189.352 ;
			LAYER M3 ;
			RECT 63.927 189.272 64.175 189.352 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[107]

	PIN Q[108]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 190.904 64.175 190.984 ;
			LAYER M2 ;
			RECT 63.927 190.904 64.175 190.984 ;
			LAYER M3 ;
			RECT 63.927 190.904 64.175 190.984 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[108]

	PIN Q[109]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 192.536 64.175 192.616 ;
			LAYER M2 ;
			RECT 63.927 192.536 64.175 192.616 ;
			LAYER M3 ;
			RECT 63.927 192.536 64.175 192.616 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[109]

	PIN Q[110]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 194.168 64.175 194.248 ;
			LAYER M2 ;
			RECT 63.927 194.168 64.175 194.248 ;
			LAYER M3 ;
			RECT 63.927 194.168 64.175 194.248 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[110]

	PIN Q[111]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 195.800 64.175 195.880 ;
			LAYER M2 ;
			RECT 63.927 195.800 64.175 195.880 ;
			LAYER M3 ;
			RECT 63.927 195.800 64.175 195.880 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[111]

	PIN Q[112]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 197.432 64.175 197.512 ;
			LAYER M2 ;
			RECT 63.927 197.432 64.175 197.512 ;
			LAYER M3 ;
			RECT 63.927 197.432 64.175 197.512 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[112]

	PIN Q[113]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 199.064 64.175 199.144 ;
			LAYER M2 ;
			RECT 63.927 199.064 64.175 199.144 ;
			LAYER M3 ;
			RECT 63.927 199.064 64.175 199.144 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[113]

	PIN Q[114]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 200.696 64.175 200.776 ;
			LAYER M2 ;
			RECT 63.927 200.696 64.175 200.776 ;
			LAYER M3 ;
			RECT 63.927 200.696 64.175 200.776 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[114]

	PIN Q[115]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 202.328 64.175 202.408 ;
			LAYER M2 ;
			RECT 63.927 202.328 64.175 202.408 ;
			LAYER M3 ;
			RECT 63.927 202.328 64.175 202.408 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[115]

	PIN Q[116]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 203.960 64.175 204.040 ;
			LAYER M2 ;
			RECT 63.927 203.960 64.175 204.040 ;
			LAYER M3 ;
			RECT 63.927 203.960 64.175 204.040 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[116]

	PIN Q[117]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 205.592 64.175 205.672 ;
			LAYER M2 ;
			RECT 63.927 205.592 64.175 205.672 ;
			LAYER M3 ;
			RECT 63.927 205.592 64.175 205.672 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[117]

	PIN Q[118]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 207.224 64.175 207.304 ;
			LAYER M2 ;
			RECT 63.927 207.224 64.175 207.304 ;
			LAYER M3 ;
			RECT 63.927 207.224 64.175 207.304 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[118]

	PIN Q[119]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 208.856 64.175 208.936 ;
			LAYER M2 ;
			RECT 63.927 208.856 64.175 208.936 ;
			LAYER M3 ;
			RECT 63.927 208.856 64.175 208.936 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[119]

	PIN Q[120]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 210.488 64.175 210.568 ;
			LAYER M2 ;
			RECT 63.927 210.488 64.175 210.568 ;
			LAYER M3 ;
			RECT 63.927 210.488 64.175 210.568 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[120]

	PIN Q[121]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 212.120 64.175 212.200 ;
			LAYER M2 ;
			RECT 63.927 212.120 64.175 212.200 ;
			LAYER M3 ;
			RECT 63.927 212.120 64.175 212.200 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[121]

	PIN Q[122]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 213.752 64.175 213.832 ;
			LAYER M2 ;
			RECT 63.927 213.752 64.175 213.832 ;
			LAYER M3 ;
			RECT 63.927 213.752 64.175 213.832 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[122]

	PIN Q[123]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 215.384 64.175 215.464 ;
			LAYER M2 ;
			RECT 63.927 215.384 64.175 215.464 ;
			LAYER M3 ;
			RECT 63.927 215.384 64.175 215.464 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[123]

	PIN Q[124]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 217.016 64.175 217.096 ;
			LAYER M2 ;
			RECT 63.927 217.016 64.175 217.096 ;
			LAYER M3 ;
			RECT 63.927 217.016 64.175 217.096 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[124]

	PIN Q[125]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 218.648 64.175 218.728 ;
			LAYER M2 ;
			RECT 63.927 218.648 64.175 218.728 ;
			LAYER M3 ;
			RECT 63.927 218.648 64.175 218.728 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[125]

	PIN Q[126]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 220.280 64.175 220.360 ;
			LAYER M2 ;
			RECT 63.927 220.280 64.175 220.360 ;
			LAYER M3 ;
			RECT 63.927 220.280 64.175 220.360 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[126]

	PIN Q[127]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 221.912 64.175 221.992 ;
			LAYER M2 ;
			RECT 63.927 221.912 64.175 221.992 ;
			LAYER M3 ;
			RECT 63.927 221.912 64.175 221.992 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[127]

	PIN Q[128]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 223.544 64.175 223.624 ;
			LAYER M2 ;
			RECT 63.927 223.544 64.175 223.624 ;
			LAYER M3 ;
			RECT 63.927 223.544 64.175 223.624 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[128]

	PIN Q[129]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 225.176 64.175 225.256 ;
			LAYER M2 ;
			RECT 63.927 225.176 64.175 225.256 ;
			LAYER M3 ;
			RECT 63.927 225.176 64.175 225.256 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[129]

	PIN Q[130]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 226.808 64.175 226.888 ;
			LAYER M2 ;
			RECT 63.927 226.808 64.175 226.888 ;
			LAYER M3 ;
			RECT 63.927 226.808 64.175 226.888 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[130]

	PIN Q[131]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 228.440 64.175 228.520 ;
			LAYER M2 ;
			RECT 63.927 228.440 64.175 228.520 ;
			LAYER M3 ;
			RECT 63.927 228.440 64.175 228.520 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[131]

	PIN Q[132]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 230.072 64.175 230.152 ;
			LAYER M2 ;
			RECT 63.927 230.072 64.175 230.152 ;
			LAYER M3 ;
			RECT 63.927 230.072 64.175 230.152 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[132]

	PIN Q[133]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 231.704 64.175 231.784 ;
			LAYER M2 ;
			RECT 63.927 231.704 64.175 231.784 ;
			LAYER M3 ;
			RECT 63.927 231.704 64.175 231.784 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[133]

	PIN Q[134]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 233.336 64.175 233.416 ;
			LAYER M2 ;
			RECT 63.927 233.336 64.175 233.416 ;
			LAYER M3 ;
			RECT 63.927 233.336 64.175 233.416 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[134]

	PIN Q[135]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 234.968 64.175 235.048 ;
			LAYER M2 ;
			RECT 63.927 234.968 64.175 235.048 ;
			LAYER M3 ;
			RECT 63.927 234.968 64.175 235.048 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[135]

	PIN Q[136]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 236.600 64.175 236.680 ;
			LAYER M2 ;
			RECT 63.927 236.600 64.175 236.680 ;
			LAYER M3 ;
			RECT 63.927 236.600 64.175 236.680 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[136]

	PIN Q[137]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 238.232 64.175 238.312 ;
			LAYER M2 ;
			RECT 63.927 238.232 64.175 238.312 ;
			LAYER M3 ;
			RECT 63.927 238.232 64.175 238.312 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[137]

	PIN Q[138]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 239.864 64.175 239.944 ;
			LAYER M2 ;
			RECT 63.927 239.864 64.175 239.944 ;
			LAYER M3 ;
			RECT 63.927 239.864 64.175 239.944 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[138]

	PIN Q[139]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 241.496 64.175 241.576 ;
			LAYER M2 ;
			RECT 63.927 241.496 64.175 241.576 ;
			LAYER M3 ;
			RECT 63.927 241.496 64.175 241.576 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[139]

	PIN Q[140]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 243.128 64.175 243.208 ;
			LAYER M2 ;
			RECT 63.927 243.128 64.175 243.208 ;
			LAYER M3 ;
			RECT 63.927 243.128 64.175 243.208 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[140]

	PIN Q[141]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 244.760 64.175 244.840 ;
			LAYER M2 ;
			RECT 63.927 244.760 64.175 244.840 ;
			LAYER M3 ;
			RECT 63.927 244.760 64.175 244.840 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[141]

	PIN Q[142]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 246.392 64.175 246.472 ;
			LAYER M2 ;
			RECT 63.927 246.392 64.175 246.472 ;
			LAYER M3 ;
			RECT 63.927 246.392 64.175 246.472 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[142]

	PIN Q[143]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 248.024 64.175 248.104 ;
			LAYER M2 ;
			RECT 63.927 248.024 64.175 248.104 ;
			LAYER M3 ;
			RECT 63.927 248.024 64.175 248.104 ;
		END
		ANTENNADIFFAREA 0.034480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.205200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.015960 LAYER VIA1 ;
		ANTENNADIFFAREA 0.034480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.283320 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNADIFFAREA 0.034480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.554520 LAYER M3 ;
	END Q[143]

	PIN RTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 130.184 64.175 130.264 ;
			LAYER M2 ;
			RECT 63.927 130.184 64.175 130.264 ;
			LAYER M3 ;
			RECT 63.927 130.184 64.175 130.264 ;
		END
		ANTENNAGATEAREA 0.003360 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.077400 LAYER M1 ;
		ANTENNAMAXAREACAR 9.919800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.289800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.003360 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.091080 LAYER M2 ;
		ANTENNAMAXAREACAR 12.849000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.579600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.003360 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.055280 LAYER M3 ;
		ANTENNAMAXAREACAR 261.708000 LAYER M3 ;
	END RTSEL[0]

	PIN RTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 130.376 64.175 130.456 ;
			LAYER M2 ;
			RECT 63.927 130.376 64.175 130.456 ;
			LAYER M3 ;
			RECT 63.927 130.376 64.175 130.456 ;
		END
		ANTENNAGATEAREA 0.003360 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.077400 LAYER M1 ;
		ANTENNAMAXAREACAR 9.919800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.289800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.003360 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.091080 LAYER M2 ;
		ANTENNAMAXAREACAR 12.849000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.579600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.003360 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.055280 LAYER M3 ;
		ANTENNAMAXAREACAR 261.708000 LAYER M3 ;
	END RTSEL[1]

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.120 0.904 64.055 1.064 ;
			LAYER M4 ;
			RECT 0.120 2.536 64.055 2.696 ;
			LAYER M4 ;
			RECT 0.120 4.168 64.055 4.328 ;
			LAYER M4 ;
			RECT 0.120 5.800 64.055 5.960 ;
			LAYER M4 ;
			RECT 0.120 7.432 64.055 7.592 ;
			LAYER M4 ;
			RECT 0.120 9.064 64.055 9.224 ;
			LAYER M4 ;
			RECT 0.120 10.696 64.055 10.856 ;
			LAYER M4 ;
			RECT 0.120 12.328 64.055 12.488 ;
			LAYER M4 ;
			RECT 0.120 13.960 64.055 14.120 ;
			LAYER M4 ;
			RECT 0.120 15.592 64.055 15.752 ;
			LAYER M4 ;
			RECT 0.120 17.224 64.055 17.384 ;
			LAYER M4 ;
			RECT 0.120 18.856 64.055 19.016 ;
			LAYER M4 ;
			RECT 0.120 20.488 64.055 20.648 ;
			LAYER M4 ;
			RECT 0.120 22.120 64.055 22.280 ;
			LAYER M4 ;
			RECT 0.120 23.752 64.055 23.912 ;
			LAYER M4 ;
			RECT 0.120 25.384 64.055 25.544 ;
			LAYER M4 ;
			RECT 0.120 27.016 64.055 27.176 ;
			LAYER M4 ;
			RECT 0.120 28.648 64.055 28.808 ;
			LAYER M4 ;
			RECT 0.120 30.280 64.055 30.440 ;
			LAYER M4 ;
			RECT 0.120 31.912 64.055 32.072 ;
			LAYER M4 ;
			RECT 0.120 33.544 64.055 33.704 ;
			LAYER M4 ;
			RECT 0.120 35.176 64.055 35.336 ;
			LAYER M4 ;
			RECT 0.120 36.808 64.055 36.968 ;
			LAYER M4 ;
			RECT 0.120 38.440 64.055 38.600 ;
			LAYER M4 ;
			RECT 0.120 40.072 64.055 40.232 ;
			LAYER M4 ;
			RECT 0.120 41.704 64.055 41.864 ;
			LAYER M4 ;
			RECT 0.120 43.336 64.055 43.496 ;
			LAYER M4 ;
			RECT 0.120 44.968 64.055 45.128 ;
			LAYER M4 ;
			RECT 0.120 46.600 64.055 46.760 ;
			LAYER M4 ;
			RECT 0.120 48.232 64.055 48.392 ;
			LAYER M4 ;
			RECT 0.120 49.864 64.055 50.024 ;
			LAYER M4 ;
			RECT 0.120 51.496 64.055 51.656 ;
			LAYER M4 ;
			RECT 0.120 53.128 64.055 53.288 ;
			LAYER M4 ;
			RECT 0.120 54.760 64.055 54.920 ;
			LAYER M4 ;
			RECT 0.120 56.392 64.055 56.552 ;
			LAYER M4 ;
			RECT 0.120 58.024 64.055 58.184 ;
			LAYER M4 ;
			RECT 0.120 59.656 64.055 59.816 ;
			LAYER M4 ;
			RECT 0.120 61.288 64.055 61.448 ;
			LAYER M4 ;
			RECT 0.120 62.920 64.055 63.080 ;
			LAYER M4 ;
			RECT 0.120 64.552 64.055 64.712 ;
			LAYER M4 ;
			RECT 0.120 66.184 64.055 66.344 ;
			LAYER M4 ;
			RECT 0.120 67.816 64.055 67.976 ;
			LAYER M4 ;
			RECT 0.120 69.448 64.055 69.608 ;
			LAYER M4 ;
			RECT 0.120 71.080 64.055 71.240 ;
			LAYER M4 ;
			RECT 0.120 72.712 64.055 72.872 ;
			LAYER M4 ;
			RECT 0.120 74.344 64.055 74.504 ;
			LAYER M4 ;
			RECT 0.120 75.976 64.055 76.136 ;
			LAYER M4 ;
			RECT 0.120 77.608 64.055 77.768 ;
			LAYER M4 ;
			RECT 0.120 79.240 64.055 79.400 ;
			LAYER M4 ;
			RECT 0.120 80.872 64.055 81.032 ;
			LAYER M4 ;
			RECT 0.120 82.504 64.055 82.664 ;
			LAYER M4 ;
			RECT 0.120 84.136 64.055 84.296 ;
			LAYER M4 ;
			RECT 0.120 85.768 64.055 85.928 ;
			LAYER M4 ;
			RECT 0.120 87.400 64.055 87.560 ;
			LAYER M4 ;
			RECT 0.120 89.032 64.055 89.192 ;
			LAYER M4 ;
			RECT 0.120 90.664 64.055 90.824 ;
			LAYER M4 ;
			RECT 0.120 92.296 64.055 92.456 ;
			LAYER M4 ;
			RECT 0.120 93.928 64.055 94.088 ;
			LAYER M4 ;
			RECT 0.120 95.560 64.055 95.720 ;
			LAYER M4 ;
			RECT 0.120 97.192 64.055 97.352 ;
			LAYER M4 ;
			RECT 0.120 98.824 64.055 98.984 ;
			LAYER M4 ;
			RECT 0.120 100.456 64.055 100.616 ;
			LAYER M4 ;
			RECT 0.120 102.088 64.055 102.248 ;
			LAYER M4 ;
			RECT 0.120 103.720 64.055 103.880 ;
			LAYER M4 ;
			RECT 0.120 105.352 64.055 105.512 ;
			LAYER M4 ;
			RECT 0.120 106.984 64.055 107.144 ;
			LAYER M4 ;
			RECT 0.120 108.616 64.055 108.776 ;
			LAYER M4 ;
			RECT 0.120 110.248 64.055 110.408 ;
			LAYER M4 ;
			RECT 0.120 111.880 64.055 112.040 ;
			LAYER M4 ;
			RECT 0.120 113.512 64.055 113.672 ;
			LAYER M4 ;
			RECT 0.120 115.144 64.055 115.304 ;
			LAYER M4 ;
			RECT 0.120 116.776 64.055 116.936 ;
			LAYER M4 ;
			RECT 0.120 118.408 64.055 118.568 ;
			LAYER M4 ;
			RECT 0.120 118.948 64.055 119.068 ;
			LAYER M4 ;
			RECT 0.120 119.572 64.055 119.692 ;
			LAYER M4 ;
			RECT 0.120 119.978 64.055 120.098 ;
			LAYER M4 ;
			RECT 0.120 120.438 64.055 120.558 ;
			LAYER M4 ;
			RECT 0.120 120.898 64.055 121.018 ;
			LAYER M4 ;
			RECT 0.120 121.358 64.055 121.478 ;
			LAYER M4 ;
			RECT 0.120 121.588 64.055 121.708 ;
			LAYER M4 ;
			RECT 0.120 121.980 64.055 122.100 ;
			LAYER M4 ;
			RECT 0.120 123.130 64.055 123.250 ;
			LAYER M4 ;
			RECT 0.120 123.812 64.055 123.932 ;
			LAYER M4 ;
			RECT 0.120 124.724 64.055 124.844 ;
			LAYER M4 ;
			RECT 0.120 125.903 64.055 126.023 ;
			LAYER M4 ;
			RECT 0.120 126.592 64.055 126.712 ;
			LAYER M4 ;
			RECT 0.120 127.052 64.055 127.172 ;
			LAYER M4 ;
			RECT 0.120 127.928 64.055 128.048 ;
			LAYER M4 ;
			RECT 0.120 128.388 64.055 128.508 ;
			LAYER M4 ;
			RECT 0.120 129.256 64.055 129.376 ;
			LAYER M4 ;
			RECT 0.120 129.690 64.055 129.810 ;
			LAYER M4 ;
			RECT 0.120 130.150 64.055 130.270 ;
			LAYER M4 ;
			RECT 0.120 130.564 64.055 130.684 ;
			LAYER M4 ;
			RECT 0.120 131.024 64.055 131.144 ;
			LAYER M4 ;
			RECT 0.120 131.272 64.055 131.432 ;
			LAYER M4 ;
			RECT 0.120 132.904 64.055 133.064 ;
			LAYER M4 ;
			RECT 0.120 134.536 64.055 134.696 ;
			LAYER M4 ;
			RECT 0.120 136.168 64.055 136.328 ;
			LAYER M4 ;
			RECT 0.120 137.800 64.055 137.960 ;
			LAYER M4 ;
			RECT 0.120 139.432 64.055 139.592 ;
			LAYER M4 ;
			RECT 0.120 141.064 64.055 141.224 ;
			LAYER M4 ;
			RECT 0.120 142.696 64.055 142.856 ;
			LAYER M4 ;
			RECT 0.120 144.328 64.055 144.488 ;
			LAYER M4 ;
			RECT 0.120 145.960 64.055 146.120 ;
			LAYER M4 ;
			RECT 0.120 147.592 64.055 147.752 ;
			LAYER M4 ;
			RECT 0.120 149.224 64.055 149.384 ;
			LAYER M4 ;
			RECT 0.120 150.856 64.055 151.016 ;
			LAYER M4 ;
			RECT 0.120 152.488 64.055 152.648 ;
			LAYER M4 ;
			RECT 0.120 154.120 64.055 154.280 ;
			LAYER M4 ;
			RECT 0.120 155.752 64.055 155.912 ;
			LAYER M4 ;
			RECT 0.120 157.384 64.055 157.544 ;
			LAYER M4 ;
			RECT 0.120 159.016 64.055 159.176 ;
			LAYER M4 ;
			RECT 0.120 160.648 64.055 160.808 ;
			LAYER M4 ;
			RECT 0.120 162.280 64.055 162.440 ;
			LAYER M4 ;
			RECT 0.120 163.912 64.055 164.072 ;
			LAYER M4 ;
			RECT 0.120 165.544 64.055 165.704 ;
			LAYER M4 ;
			RECT 0.120 167.176 64.055 167.336 ;
			LAYER M4 ;
			RECT 0.120 168.808 64.055 168.968 ;
			LAYER M4 ;
			RECT 0.120 170.440 64.055 170.600 ;
			LAYER M4 ;
			RECT 0.120 172.072 64.055 172.232 ;
			LAYER M4 ;
			RECT 0.120 173.704 64.055 173.864 ;
			LAYER M4 ;
			RECT 0.120 175.336 64.055 175.496 ;
			LAYER M4 ;
			RECT 0.120 176.968 64.055 177.128 ;
			LAYER M4 ;
			RECT 0.120 178.600 64.055 178.760 ;
			LAYER M4 ;
			RECT 0.120 180.232 64.055 180.392 ;
			LAYER M4 ;
			RECT 0.120 181.864 64.055 182.024 ;
			LAYER M4 ;
			RECT 0.120 183.496 64.055 183.656 ;
			LAYER M4 ;
			RECT 0.120 185.128 64.055 185.288 ;
			LAYER M4 ;
			RECT 0.120 186.760 64.055 186.920 ;
			LAYER M4 ;
			RECT 0.120 188.392 64.055 188.552 ;
			LAYER M4 ;
			RECT 0.120 190.024 64.055 190.184 ;
			LAYER M4 ;
			RECT 0.120 191.656 64.055 191.816 ;
			LAYER M4 ;
			RECT 0.120 193.288 64.055 193.448 ;
			LAYER M4 ;
			RECT 0.120 194.920 64.055 195.080 ;
			LAYER M4 ;
			RECT 0.120 196.552 64.055 196.712 ;
			LAYER M4 ;
			RECT 0.120 198.184 64.055 198.344 ;
			LAYER M4 ;
			RECT 0.120 199.816 64.055 199.976 ;
			LAYER M4 ;
			RECT 0.120 201.448 64.055 201.608 ;
			LAYER M4 ;
			RECT 0.120 203.080 64.055 203.240 ;
			LAYER M4 ;
			RECT 0.120 204.712 64.055 204.872 ;
			LAYER M4 ;
			RECT 0.120 206.344 64.055 206.504 ;
			LAYER M4 ;
			RECT 0.120 207.976 64.055 208.136 ;
			LAYER M4 ;
			RECT 0.120 209.608 64.055 209.768 ;
			LAYER M4 ;
			RECT 0.120 211.240 64.055 211.400 ;
			LAYER M4 ;
			RECT 0.120 212.872 64.055 213.032 ;
			LAYER M4 ;
			RECT 0.120 214.504 64.055 214.664 ;
			LAYER M4 ;
			RECT 0.120 216.136 64.055 216.296 ;
			LAYER M4 ;
			RECT 0.120 217.768 64.055 217.928 ;
			LAYER M4 ;
			RECT 0.120 219.400 64.055 219.560 ;
			LAYER M4 ;
			RECT 0.120 221.032 64.055 221.192 ;
			LAYER M4 ;
			RECT 0.120 222.664 64.055 222.824 ;
			LAYER M4 ;
			RECT 0.120 224.296 64.055 224.456 ;
			LAYER M4 ;
			RECT 0.120 225.928 64.055 226.088 ;
			LAYER M4 ;
			RECT 0.120 227.560 64.055 227.720 ;
			LAYER M4 ;
			RECT 0.120 229.192 64.055 229.352 ;
			LAYER M4 ;
			RECT 0.120 230.824 64.055 230.984 ;
			LAYER M4 ;
			RECT 0.120 232.456 64.055 232.616 ;
			LAYER M4 ;
			RECT 0.120 234.088 64.055 234.248 ;
			LAYER M4 ;
			RECT 0.120 235.720 64.055 235.880 ;
			LAYER M4 ;
			RECT 0.120 237.352 64.055 237.512 ;
			LAYER M4 ;
			RECT 0.120 238.984 64.055 239.144 ;
			LAYER M4 ;
			RECT 0.120 240.616 64.055 240.776 ;
			LAYER M4 ;
			RECT 0.120 242.248 64.055 242.408 ;
			LAYER M4 ;
			RECT 0.120 243.880 64.055 244.040 ;
			LAYER M4 ;
			RECT 0.120 245.512 64.055 245.672 ;
			LAYER M4 ;
			RECT 0.120 247.144 64.055 247.304 ;
			LAYER M4 ;
			RECT 0.120 248.776 64.055 248.936 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 0.120 1.312 64.055 1.472 ;
			LAYER M4 ;
			RECT 0.120 2.128 64.055 2.288 ;
			LAYER M4 ;
			RECT 0.120 2.944 64.055 3.104 ;
			LAYER M4 ;
			RECT 0.120 3.760 64.055 3.920 ;
			LAYER M4 ;
			RECT 0.120 4.576 64.055 4.736 ;
			LAYER M4 ;
			RECT 0.120 5.392 64.055 5.552 ;
			LAYER M4 ;
			RECT 0.120 6.208 64.055 6.368 ;
			LAYER M4 ;
			RECT 0.120 7.024 64.055 7.184 ;
			LAYER M4 ;
			RECT 0.120 7.840 64.055 8.000 ;
			LAYER M4 ;
			RECT 0.120 8.656 64.055 8.816 ;
			LAYER M4 ;
			RECT 0.120 9.472 64.055 9.632 ;
			LAYER M4 ;
			RECT 0.120 10.288 64.055 10.448 ;
			LAYER M4 ;
			RECT 0.120 11.104 64.055 11.264 ;
			LAYER M4 ;
			RECT 0.120 11.920 64.055 12.080 ;
			LAYER M4 ;
			RECT 0.120 12.736 64.055 12.896 ;
			LAYER M4 ;
			RECT 0.120 13.552 64.055 13.712 ;
			LAYER M4 ;
			RECT 0.120 14.368 64.055 14.528 ;
			LAYER M4 ;
			RECT 0.120 15.184 64.055 15.344 ;
			LAYER M4 ;
			RECT 0.120 16.000 64.055 16.160 ;
			LAYER M4 ;
			RECT 0.120 16.816 64.055 16.976 ;
			LAYER M4 ;
			RECT 0.120 17.632 64.055 17.792 ;
			LAYER M4 ;
			RECT 0.120 18.448 64.055 18.608 ;
			LAYER M4 ;
			RECT 0.120 19.264 64.055 19.424 ;
			LAYER M4 ;
			RECT 0.120 20.080 64.055 20.240 ;
			LAYER M4 ;
			RECT 0.120 20.896 64.055 21.056 ;
			LAYER M4 ;
			RECT 0.120 21.712 64.055 21.872 ;
			LAYER M4 ;
			RECT 0.120 22.528 64.055 22.688 ;
			LAYER M4 ;
			RECT 0.120 23.344 64.055 23.504 ;
			LAYER M4 ;
			RECT 0.120 24.160 64.055 24.320 ;
			LAYER M4 ;
			RECT 0.120 24.976 64.055 25.136 ;
			LAYER M4 ;
			RECT 0.120 25.792 64.055 25.952 ;
			LAYER M4 ;
			RECT 0.120 26.608 64.055 26.768 ;
			LAYER M4 ;
			RECT 0.120 27.424 64.055 27.584 ;
			LAYER M4 ;
			RECT 0.120 28.240 64.055 28.400 ;
			LAYER M4 ;
			RECT 0.120 29.056 64.055 29.216 ;
			LAYER M4 ;
			RECT 0.120 29.872 64.055 30.032 ;
			LAYER M4 ;
			RECT 0.120 30.688 64.055 30.848 ;
			LAYER M4 ;
			RECT 0.120 31.504 64.055 31.664 ;
			LAYER M4 ;
			RECT 0.120 32.320 64.055 32.480 ;
			LAYER M4 ;
			RECT 0.120 33.136 64.055 33.296 ;
			LAYER M4 ;
			RECT 0.120 33.952 64.055 34.112 ;
			LAYER M4 ;
			RECT 0.120 34.768 64.055 34.928 ;
			LAYER M4 ;
			RECT 0.120 35.584 64.055 35.744 ;
			LAYER M4 ;
			RECT 0.120 36.400 64.055 36.560 ;
			LAYER M4 ;
			RECT 0.120 37.216 64.055 37.376 ;
			LAYER M4 ;
			RECT 0.120 38.032 64.055 38.192 ;
			LAYER M4 ;
			RECT 0.120 38.848 64.055 39.008 ;
			LAYER M4 ;
			RECT 0.120 39.664 64.055 39.824 ;
			LAYER M4 ;
			RECT 0.120 40.480 64.055 40.640 ;
			LAYER M4 ;
			RECT 0.120 41.296 64.055 41.456 ;
			LAYER M4 ;
			RECT 0.120 42.112 64.055 42.272 ;
			LAYER M4 ;
			RECT 0.120 42.928 64.055 43.088 ;
			LAYER M4 ;
			RECT 0.120 43.744 64.055 43.904 ;
			LAYER M4 ;
			RECT 0.120 44.560 64.055 44.720 ;
			LAYER M4 ;
			RECT 0.120 45.376 64.055 45.536 ;
			LAYER M4 ;
			RECT 0.120 46.192 64.055 46.352 ;
			LAYER M4 ;
			RECT 0.120 47.008 64.055 47.168 ;
			LAYER M4 ;
			RECT 0.120 47.824 64.055 47.984 ;
			LAYER M4 ;
			RECT 0.120 48.640 64.055 48.800 ;
			LAYER M4 ;
			RECT 0.120 49.456 64.055 49.616 ;
			LAYER M4 ;
			RECT 0.120 50.272 64.055 50.432 ;
			LAYER M4 ;
			RECT 0.120 51.088 64.055 51.248 ;
			LAYER M4 ;
			RECT 0.120 51.904 64.055 52.064 ;
			LAYER M4 ;
			RECT 0.120 52.720 64.055 52.880 ;
			LAYER M4 ;
			RECT 0.120 53.536 64.055 53.696 ;
			LAYER M4 ;
			RECT 0.120 54.352 64.055 54.512 ;
			LAYER M4 ;
			RECT 0.120 55.168 64.055 55.328 ;
			LAYER M4 ;
			RECT 0.120 55.984 64.055 56.144 ;
			LAYER M4 ;
			RECT 0.120 56.800 64.055 56.960 ;
			LAYER M4 ;
			RECT 0.120 57.616 64.055 57.776 ;
			LAYER M4 ;
			RECT 0.120 58.432 64.055 58.592 ;
			LAYER M4 ;
			RECT 0.120 59.248 64.055 59.408 ;
			LAYER M4 ;
			RECT 0.120 60.064 64.055 60.224 ;
			LAYER M4 ;
			RECT 0.120 60.880 64.055 61.040 ;
			LAYER M4 ;
			RECT 0.120 61.696 64.055 61.856 ;
			LAYER M4 ;
			RECT 0.120 62.512 64.055 62.672 ;
			LAYER M4 ;
			RECT 0.120 63.328 64.055 63.488 ;
			LAYER M4 ;
			RECT 0.120 64.144 64.055 64.304 ;
			LAYER M4 ;
			RECT 0.120 64.960 64.055 65.120 ;
			LAYER M4 ;
			RECT 0.120 65.776 64.055 65.936 ;
			LAYER M4 ;
			RECT 0.120 66.592 64.055 66.752 ;
			LAYER M4 ;
			RECT 0.120 67.408 64.055 67.568 ;
			LAYER M4 ;
			RECT 0.120 68.224 64.055 68.384 ;
			LAYER M4 ;
			RECT 0.120 69.040 64.055 69.200 ;
			LAYER M4 ;
			RECT 0.120 69.856 64.055 70.016 ;
			LAYER M4 ;
			RECT 0.120 70.672 64.055 70.832 ;
			LAYER M4 ;
			RECT 0.120 71.488 64.055 71.648 ;
			LAYER M4 ;
			RECT 0.120 72.304 64.055 72.464 ;
			LAYER M4 ;
			RECT 0.120 73.120 64.055 73.280 ;
			LAYER M4 ;
			RECT 0.120 73.936 64.055 74.096 ;
			LAYER M4 ;
			RECT 0.120 74.752 64.055 74.912 ;
			LAYER M4 ;
			RECT 0.120 75.568 64.055 75.728 ;
			LAYER M4 ;
			RECT 0.120 76.384 64.055 76.544 ;
			LAYER M4 ;
			RECT 0.120 77.200 64.055 77.360 ;
			LAYER M4 ;
			RECT 0.120 78.016 64.055 78.176 ;
			LAYER M4 ;
			RECT 0.120 78.832 64.055 78.992 ;
			LAYER M4 ;
			RECT 0.120 79.648 64.055 79.808 ;
			LAYER M4 ;
			RECT 0.120 80.464 64.055 80.624 ;
			LAYER M4 ;
			RECT 0.120 81.280 64.055 81.440 ;
			LAYER M4 ;
			RECT 0.120 82.096 64.055 82.256 ;
			LAYER M4 ;
			RECT 0.120 82.912 64.055 83.072 ;
			LAYER M4 ;
			RECT 0.120 83.728 64.055 83.888 ;
			LAYER M4 ;
			RECT 0.120 84.544 64.055 84.704 ;
			LAYER M4 ;
			RECT 0.120 85.360 64.055 85.520 ;
			LAYER M4 ;
			RECT 0.120 86.176 64.055 86.336 ;
			LAYER M4 ;
			RECT 0.120 86.992 64.055 87.152 ;
			LAYER M4 ;
			RECT 0.120 87.808 64.055 87.968 ;
			LAYER M4 ;
			RECT 0.120 88.624 64.055 88.784 ;
			LAYER M4 ;
			RECT 0.120 89.440 64.055 89.600 ;
			LAYER M4 ;
			RECT 0.120 90.256 64.055 90.416 ;
			LAYER M4 ;
			RECT 0.120 91.072 64.055 91.232 ;
			LAYER M4 ;
			RECT 0.120 91.888 64.055 92.048 ;
			LAYER M4 ;
			RECT 0.120 92.704 64.055 92.864 ;
			LAYER M4 ;
			RECT 0.120 93.520 64.055 93.680 ;
			LAYER M4 ;
			RECT 0.120 94.336 64.055 94.496 ;
			LAYER M4 ;
			RECT 0.120 95.152 64.055 95.312 ;
			LAYER M4 ;
			RECT 0.120 95.968 64.055 96.128 ;
			LAYER M4 ;
			RECT 0.120 96.784 64.055 96.944 ;
			LAYER M4 ;
			RECT 0.120 97.600 64.055 97.760 ;
			LAYER M4 ;
			RECT 0.120 98.416 64.055 98.576 ;
			LAYER M4 ;
			RECT 0.120 99.232 64.055 99.392 ;
			LAYER M4 ;
			RECT 0.120 100.048 64.055 100.208 ;
			LAYER M4 ;
			RECT 0.120 100.864 64.055 101.024 ;
			LAYER M4 ;
			RECT 0.120 101.680 64.055 101.840 ;
			LAYER M4 ;
			RECT 0.120 102.496 64.055 102.656 ;
			LAYER M4 ;
			RECT 0.120 103.312 64.055 103.472 ;
			LAYER M4 ;
			RECT 0.120 104.128 64.055 104.288 ;
			LAYER M4 ;
			RECT 0.120 104.944 64.055 105.104 ;
			LAYER M4 ;
			RECT 0.120 105.760 64.055 105.920 ;
			LAYER M4 ;
			RECT 0.120 106.576 64.055 106.736 ;
			LAYER M4 ;
			RECT 0.120 107.392 64.055 107.552 ;
			LAYER M4 ;
			RECT 0.120 108.208 64.055 108.368 ;
			LAYER M4 ;
			RECT 0.120 109.024 64.055 109.184 ;
			LAYER M4 ;
			RECT 0.120 109.840 64.055 110.000 ;
			LAYER M4 ;
			RECT 0.120 110.656 64.055 110.816 ;
			LAYER M4 ;
			RECT 0.120 111.472 64.055 111.632 ;
			LAYER M4 ;
			RECT 0.120 112.288 64.055 112.448 ;
			LAYER M4 ;
			RECT 0.120 113.104 64.055 113.264 ;
			LAYER M4 ;
			RECT 0.120 113.920 64.055 114.080 ;
			LAYER M4 ;
			RECT 0.120 114.736 64.055 114.896 ;
			LAYER M4 ;
			RECT 0.120 115.552 64.055 115.712 ;
			LAYER M4 ;
			RECT 0.120 116.368 64.055 116.528 ;
			LAYER M4 ;
			RECT 0.120 117.184 64.055 117.344 ;
			LAYER M4 ;
			RECT 0.120 118.000 64.055 118.160 ;
			LAYER M4 ;
			RECT 0.120 119.342 64.055 119.462 ;
			LAYER M4 ;
			RECT 0.120 120.208 64.055 120.328 ;
			LAYER M4 ;
			RECT 0.120 120.668 64.055 120.788 ;
			LAYER M4 ;
			RECT 0.120 121.128 64.055 121.248 ;
			LAYER M4 ;
			RECT 0.120 122.210 64.055 122.330 ;
			LAYER M4 ;
			RECT 0.120 122.900 64.055 123.020 ;
			LAYER M4 ;
			RECT 0.120 124.042 64.055 124.162 ;
			LAYER M4 ;
			RECT 0.120 124.954 64.055 125.074 ;
			LAYER M4 ;
			RECT 0.120 125.673 64.055 125.793 ;
			LAYER M4 ;
			RECT 0.120 126.822 64.055 126.942 ;
			LAYER M4 ;
			RECT 0.120 127.282 64.055 127.402 ;
			LAYER M4 ;
			RECT 0.120 127.698 64.055 127.818 ;
			LAYER M4 ;
			RECT 0.120 128.158 64.055 128.278 ;
			LAYER M4 ;
			RECT 0.120 128.618 64.055 128.738 ;
			LAYER M4 ;
			RECT 0.120 129.026 64.055 129.146 ;
			LAYER M4 ;
			RECT 0.120 129.920 64.055 130.040 ;
			LAYER M4 ;
			RECT 0.120 130.794 64.055 130.914 ;
			LAYER M4 ;
			RECT 0.120 131.680 64.055 131.840 ;
			LAYER M4 ;
			RECT 0.120 132.496 64.055 132.656 ;
			LAYER M4 ;
			RECT 0.120 133.312 64.055 133.472 ;
			LAYER M4 ;
			RECT 0.120 134.128 64.055 134.288 ;
			LAYER M4 ;
			RECT 0.120 134.944 64.055 135.104 ;
			LAYER M4 ;
			RECT 0.120 135.760 64.055 135.920 ;
			LAYER M4 ;
			RECT 0.120 136.576 64.055 136.736 ;
			LAYER M4 ;
			RECT 0.120 137.392 64.055 137.552 ;
			LAYER M4 ;
			RECT 0.120 138.208 64.055 138.368 ;
			LAYER M4 ;
			RECT 0.120 139.024 64.055 139.184 ;
			LAYER M4 ;
			RECT 0.120 139.840 64.055 140.000 ;
			LAYER M4 ;
			RECT 0.120 140.656 64.055 140.816 ;
			LAYER M4 ;
			RECT 0.120 141.472 64.055 141.632 ;
			LAYER M4 ;
			RECT 0.120 142.288 64.055 142.448 ;
			LAYER M4 ;
			RECT 0.120 143.104 64.055 143.264 ;
			LAYER M4 ;
			RECT 0.120 143.920 64.055 144.080 ;
			LAYER M4 ;
			RECT 0.120 144.736 64.055 144.896 ;
			LAYER M4 ;
			RECT 0.120 145.552 64.055 145.712 ;
			LAYER M4 ;
			RECT 0.120 146.368 64.055 146.528 ;
			LAYER M4 ;
			RECT 0.120 147.184 64.055 147.344 ;
			LAYER M4 ;
			RECT 0.120 148.000 64.055 148.160 ;
			LAYER M4 ;
			RECT 0.120 148.816 64.055 148.976 ;
			LAYER M4 ;
			RECT 0.120 149.632 64.055 149.792 ;
			LAYER M4 ;
			RECT 0.120 150.448 64.055 150.608 ;
			LAYER M4 ;
			RECT 0.120 151.264 64.055 151.424 ;
			LAYER M4 ;
			RECT 0.120 152.080 64.055 152.240 ;
			LAYER M4 ;
			RECT 0.120 152.896 64.055 153.056 ;
			LAYER M4 ;
			RECT 0.120 153.712 64.055 153.872 ;
			LAYER M4 ;
			RECT 0.120 154.528 64.055 154.688 ;
			LAYER M4 ;
			RECT 0.120 155.344 64.055 155.504 ;
			LAYER M4 ;
			RECT 0.120 156.160 64.055 156.320 ;
			LAYER M4 ;
			RECT 0.120 156.976 64.055 157.136 ;
			LAYER M4 ;
			RECT 0.120 157.792 64.055 157.952 ;
			LAYER M4 ;
			RECT 0.120 158.608 64.055 158.768 ;
			LAYER M4 ;
			RECT 0.120 159.424 64.055 159.584 ;
			LAYER M4 ;
			RECT 0.120 160.240 64.055 160.400 ;
			LAYER M4 ;
			RECT 0.120 161.056 64.055 161.216 ;
			LAYER M4 ;
			RECT 0.120 161.872 64.055 162.032 ;
			LAYER M4 ;
			RECT 0.120 162.688 64.055 162.848 ;
			LAYER M4 ;
			RECT 0.120 163.504 64.055 163.664 ;
			LAYER M4 ;
			RECT 0.120 164.320 64.055 164.480 ;
			LAYER M4 ;
			RECT 0.120 165.136 64.055 165.296 ;
			LAYER M4 ;
			RECT 0.120 165.952 64.055 166.112 ;
			LAYER M4 ;
			RECT 0.120 166.768 64.055 166.928 ;
			LAYER M4 ;
			RECT 0.120 167.584 64.055 167.744 ;
			LAYER M4 ;
			RECT 0.120 168.400 64.055 168.560 ;
			LAYER M4 ;
			RECT 0.120 169.216 64.055 169.376 ;
			LAYER M4 ;
			RECT 0.120 170.032 64.055 170.192 ;
			LAYER M4 ;
			RECT 0.120 170.848 64.055 171.008 ;
			LAYER M4 ;
			RECT 0.120 171.664 64.055 171.824 ;
			LAYER M4 ;
			RECT 0.120 172.480 64.055 172.640 ;
			LAYER M4 ;
			RECT 0.120 173.296 64.055 173.456 ;
			LAYER M4 ;
			RECT 0.120 174.112 64.055 174.272 ;
			LAYER M4 ;
			RECT 0.120 174.928 64.055 175.088 ;
			LAYER M4 ;
			RECT 0.120 175.744 64.055 175.904 ;
			LAYER M4 ;
			RECT 0.120 176.560 64.055 176.720 ;
			LAYER M4 ;
			RECT 0.120 177.376 64.055 177.536 ;
			LAYER M4 ;
			RECT 0.120 178.192 64.055 178.352 ;
			LAYER M4 ;
			RECT 0.120 179.008 64.055 179.168 ;
			LAYER M4 ;
			RECT 0.120 179.824 64.055 179.984 ;
			LAYER M4 ;
			RECT 0.120 180.640 64.055 180.800 ;
			LAYER M4 ;
			RECT 0.120 181.456 64.055 181.616 ;
			LAYER M4 ;
			RECT 0.120 182.272 64.055 182.432 ;
			LAYER M4 ;
			RECT 0.120 183.088 64.055 183.248 ;
			LAYER M4 ;
			RECT 0.120 183.904 64.055 184.064 ;
			LAYER M4 ;
			RECT 0.120 184.720 64.055 184.880 ;
			LAYER M4 ;
			RECT 0.120 185.536 64.055 185.696 ;
			LAYER M4 ;
			RECT 0.120 186.352 64.055 186.512 ;
			LAYER M4 ;
			RECT 0.120 187.168 64.055 187.328 ;
			LAYER M4 ;
			RECT 0.120 187.984 64.055 188.144 ;
			LAYER M4 ;
			RECT 0.120 188.800 64.055 188.960 ;
			LAYER M4 ;
			RECT 0.120 189.616 64.055 189.776 ;
			LAYER M4 ;
			RECT 0.120 190.432 64.055 190.592 ;
			LAYER M4 ;
			RECT 0.120 191.248 64.055 191.408 ;
			LAYER M4 ;
			RECT 0.120 192.064 64.055 192.224 ;
			LAYER M4 ;
			RECT 0.120 192.880 64.055 193.040 ;
			LAYER M4 ;
			RECT 0.120 193.696 64.055 193.856 ;
			LAYER M4 ;
			RECT 0.120 194.512 64.055 194.672 ;
			LAYER M4 ;
			RECT 0.120 195.328 64.055 195.488 ;
			LAYER M4 ;
			RECT 0.120 196.144 64.055 196.304 ;
			LAYER M4 ;
			RECT 0.120 196.960 64.055 197.120 ;
			LAYER M4 ;
			RECT 0.120 197.776 64.055 197.936 ;
			LAYER M4 ;
			RECT 0.120 198.592 64.055 198.752 ;
			LAYER M4 ;
			RECT 0.120 199.408 64.055 199.568 ;
			LAYER M4 ;
			RECT 0.120 200.224 64.055 200.384 ;
			LAYER M4 ;
			RECT 0.120 201.040 64.055 201.200 ;
			LAYER M4 ;
			RECT 0.120 201.856 64.055 202.016 ;
			LAYER M4 ;
			RECT 0.120 202.672 64.055 202.832 ;
			LAYER M4 ;
			RECT 0.120 203.488 64.055 203.648 ;
			LAYER M4 ;
			RECT 0.120 204.304 64.055 204.464 ;
			LAYER M4 ;
			RECT 0.120 205.120 64.055 205.280 ;
			LAYER M4 ;
			RECT 0.120 205.936 64.055 206.096 ;
			LAYER M4 ;
			RECT 0.120 206.752 64.055 206.912 ;
			LAYER M4 ;
			RECT 0.120 207.568 64.055 207.728 ;
			LAYER M4 ;
			RECT 0.120 208.384 64.055 208.544 ;
			LAYER M4 ;
			RECT 0.120 209.200 64.055 209.360 ;
			LAYER M4 ;
			RECT 0.120 210.016 64.055 210.176 ;
			LAYER M4 ;
			RECT 0.120 210.832 64.055 210.992 ;
			LAYER M4 ;
			RECT 0.120 211.648 64.055 211.808 ;
			LAYER M4 ;
			RECT 0.120 212.464 64.055 212.624 ;
			LAYER M4 ;
			RECT 0.120 213.280 64.055 213.440 ;
			LAYER M4 ;
			RECT 0.120 214.096 64.055 214.256 ;
			LAYER M4 ;
			RECT 0.120 214.912 64.055 215.072 ;
			LAYER M4 ;
			RECT 0.120 215.728 64.055 215.888 ;
			LAYER M4 ;
			RECT 0.120 216.544 64.055 216.704 ;
			LAYER M4 ;
			RECT 0.120 217.360 64.055 217.520 ;
			LAYER M4 ;
			RECT 0.120 218.176 64.055 218.336 ;
			LAYER M4 ;
			RECT 0.120 218.992 64.055 219.152 ;
			LAYER M4 ;
			RECT 0.120 219.808 64.055 219.968 ;
			LAYER M4 ;
			RECT 0.120 220.624 64.055 220.784 ;
			LAYER M4 ;
			RECT 0.120 221.440 64.055 221.600 ;
			LAYER M4 ;
			RECT 0.120 222.256 64.055 222.416 ;
			LAYER M4 ;
			RECT 0.120 223.072 64.055 223.232 ;
			LAYER M4 ;
			RECT 0.120 223.888 64.055 224.048 ;
			LAYER M4 ;
			RECT 0.120 224.704 64.055 224.864 ;
			LAYER M4 ;
			RECT 0.120 225.520 64.055 225.680 ;
			LAYER M4 ;
			RECT 0.120 226.336 64.055 226.496 ;
			LAYER M4 ;
			RECT 0.120 227.152 64.055 227.312 ;
			LAYER M4 ;
			RECT 0.120 227.968 64.055 228.128 ;
			LAYER M4 ;
			RECT 0.120 228.784 64.055 228.944 ;
			LAYER M4 ;
			RECT 0.120 229.600 64.055 229.760 ;
			LAYER M4 ;
			RECT 0.120 230.416 64.055 230.576 ;
			LAYER M4 ;
			RECT 0.120 231.232 64.055 231.392 ;
			LAYER M4 ;
			RECT 0.120 232.048 64.055 232.208 ;
			LAYER M4 ;
			RECT 0.120 232.864 64.055 233.024 ;
			LAYER M4 ;
			RECT 0.120 233.680 64.055 233.840 ;
			LAYER M4 ;
			RECT 0.120 234.496 64.055 234.656 ;
			LAYER M4 ;
			RECT 0.120 235.312 64.055 235.472 ;
			LAYER M4 ;
			RECT 0.120 236.128 64.055 236.288 ;
			LAYER M4 ;
			RECT 0.120 236.944 64.055 237.104 ;
			LAYER M4 ;
			RECT 0.120 237.760 64.055 237.920 ;
			LAYER M4 ;
			RECT 0.120 238.576 64.055 238.736 ;
			LAYER M4 ;
			RECT 0.120 239.392 64.055 239.552 ;
			LAYER M4 ;
			RECT 0.120 240.208 64.055 240.368 ;
			LAYER M4 ;
			RECT 0.120 241.024 64.055 241.184 ;
			LAYER M4 ;
			RECT 0.120 241.840 64.055 242.000 ;
			LAYER M4 ;
			RECT 0.120 242.656 64.055 242.816 ;
			LAYER M4 ;
			RECT 0.120 243.472 64.055 243.632 ;
			LAYER M4 ;
			RECT 0.120 244.288 64.055 244.448 ;
			LAYER M4 ;
			RECT 0.120 245.104 64.055 245.264 ;
			LAYER M4 ;
			RECT 0.120 245.920 64.055 246.080 ;
			LAYER M4 ;
			RECT 0.120 246.736 64.055 246.896 ;
			LAYER M4 ;
			RECT 0.120 247.552 64.055 247.712 ;
			LAYER M4 ;
			RECT 0.120 248.368 64.055 248.528 ;
		END
	END VSS

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 123.080 64.175 123.160 ;
			LAYER M2 ;
			RECT 63.927 123.080 64.175 123.160 ;
			LAYER M3 ;
			RECT 63.927 123.080 64.175 123.160 ;
		END
		ANTENNAGATEAREA 0.006480 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.067800 LAYER M1 ;
		ANTENNAMAXAREACAR 4.009920 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.152040 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006480 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.082320 LAYER M2 ;
		ANTENNAMAXAREACAR 7.834200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.304200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006480 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.113520 LAYER M3 ;
		ANTENNAMAXAREACAR 21.891100 LAYER M3 ;
	END WEB

	PIN WTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 122.888 64.175 122.968 ;
			LAYER M2 ;
			RECT 63.927 122.888 64.175 122.968 ;
			LAYER M3 ;
			RECT 63.927 122.888 64.175 122.968 ;
		END
		ANTENNAGATEAREA 0.003360 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.060360 LAYER M1 ;
		ANTENNAMAXAREACAR 5.886840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.289800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.003360 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.138360 LAYER M2 ;
		ANTENNAMAXAREACAR 27.863200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.579600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.003360 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.810960 LAYER M3 ;
		ANTENNAMAXAREACAR 199.728000 LAYER M3 ;
	END WTSEL[0]

	PIN WTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.927 124.040 64.175 124.120 ;
			LAYER M2 ;
			RECT 63.927 124.040 64.175 124.120 ;
			LAYER M3 ;
			RECT 63.927 124.040 64.175 124.120 ;
		END
		ANTENNAGATEAREA 0.003360 LAYER M1 ;
		ANTENNADIFFAREA 0.006480 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.060360 LAYER M1 ;
		ANTENNAMAXAREACAR 5.886840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.289800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.003360 LAYER M2 ;
		ANTENNADIFFAREA 0.006480 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.138360 LAYER M2 ;
		ANTENNAMAXAREACAR 27.863200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.579600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.003360 LAYER M3 ;
		ANTENNADIFFAREA 0.006480 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.810960 LAYER M3 ;
		ANTENNAMAXAREACAR 199.728000 LAYER M3 ;
	END WTSEL[1]

	OBS
		LAYER M1 SPACING 0.000 ;
		RECT 0.000 0.000 64.175 249.840 ;
		LAYER M2 SPACING 0.000 ;
		RECT 0.000 0.000 64.175 249.840 ;
		LAYER M3 SPACING 0.000 ;
		RECT 0.000 0.000 64.175 249.840 ;
		LAYER M4 ;
		RECT 0.400 0.431 63.775 0.551 ;
		LAYER M4 ;
		RECT 0.400 249.289 63.775 249.409 ;
		LAYER M4 ;
		RECT 0.783 130.360 58.953 130.437 ;
		LAYER M4 ;
		RECT 1.218 123.317 58.953 123.415 ;
		LAYER M4 ;
		RECT 1.218 123.497 58.953 123.595 ;
		LAYER M4 ;
		RECT 1.218 123.677 58.953 123.775 ;
		LAYER M4 ;
		RECT 1.218 124.229 58.953 124.327 ;
		LAYER M4 ;
		RECT 1.218 124.409 58.953 124.507 ;
		LAYER M4 ;
		RECT 1.218 124.589 58.953 124.687 ;
		LAYER M4 ;
		RECT 1.218 125.175 58.953 125.273 ;
		LAYER M4 ;
		RECT 1.218 125.355 58.953 125.453 ;
		LAYER M4 ;
		RECT 1.218 125.535 58.953 125.633 ;
		LAYER M4 ;
		RECT 1.218 126.087 58.953 126.185 ;
		LAYER M4 ;
		RECT 1.218 126.267 58.953 126.365 ;
		LAYER M4 ;
		RECT 1.218 126.447 58.953 126.545 ;
		LAYER M4 ;
		RECT 1.627 122.365 58.953 122.463 ;
		LAYER M4 ;
		RECT 1.627 122.545 58.953 122.643 ;
		LAYER M4 ;
		RECT 1.627 122.725 58.953 122.823 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 64.175 249.840 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 64.175 249.840 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 64.175 249.840 ;
	END
END TS1N16FFCLLSBLVTC1024X144M4SW

END LIBRARY
