should try this pipcleaner during this weekend(3rd/Apr/2021)
