magic
tech sky130A
timestamp 1619949044
<< dnwell >>
rect 759 5481 877 5599
rect 534 4966 652 5084
rect 776 5003 894 5121
rect 1012 4985 1130 5103
rect 1255 4965 1373 5083
rect 1441 4969 1559 5087
rect 1631 4976 1749 5094
<< metal3 >>
rect 2939 -652 4545 66
<< via4 >>
rect 88 5407 206 5525
rect 526 5420 644 5538
rect 759 5481 877 5599
rect 534 4966 652 5084
rect 776 5003 894 5121
rect 1012 4985 1130 5103
rect 1255 4965 1373 5083
rect 1441 4969 1559 5087
rect 1631 4976 1749 5094
<< metal5 >>
rect 2908 19715 4514 20433
rect -1030 19099 -467 19126
rect -1030 17920 1759 19099
rect -1030 6258 -467 17920
rect 2882 15120 4488 15838
rect 7922 7728 8606 7782
rect 6951 7213 8606 7728
rect 0 6744 427 7130
rect -1408 5525 468 6258
rect -1408 5407 88 5525
rect 206 5407 468 5525
rect -1408 3981 468 5407
rect -1408 3890 541 3981
rect -1408 2597 468 3890
rect 7922 2383 8606 7213
rect 385 319 1347 2349
rect 7206 2042 8606 2383
rect 7206 2035 8539 2042
use test  test_0
timestamp 1619945680
transform 1 0 0 0 1 0
box 0 0 7500 20000
<< labels >>
flabel metal5 385 319 1347 2349 1 FreeSans 3200 0 0 0 VDD
port 3 n
flabel metal3 2939 -652 4545 66 1 FreeSans 3200 0 0 0 in
port 1 n
flabel metal5 2882 15120 4488 15838 1 FreeSans 3200 0 0 0 out
port 2 n
flabel metal5 2908 19715 4514 20433 1 FreeSans 3200 0 0 0 GND
port 4 n
<< end >>
