magic
tech sky130A
magscale 1 2
timestamp 1619862920
<< checkpaint >>
rect -1288 -1260 1388 1323
use sky130_fd_pr__hvdfl1sd__example_55959141808280  sky130_fd_pr__hvdfl1sd__example_55959141808280_0
timestamp 1619862920
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808510  sky130_fd_pr__dfl1sd__example_55959141808510_0
timestamp 1619862920
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 128 63 128 63 0 FreeSans 300 0 0 0 D
flabel comment s -28 63 -28 63 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 48196018
string GDS_START 48195094
<< end >>
