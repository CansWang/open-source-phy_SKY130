magic
tech sky130A
magscale 1 2
timestamp 1619341889
<< nwell >>
rect -111 263 1134 584
<< pwell >>
rect 19 -15 53 19
rect 434 -15 468 19
rect 849 -15 883 19
<< scnmos >>
rect 110 49 140 179
rect 525 49 555 179
rect 940 49 970 179
<< scpmoshvt >>
rect 110 299 140 499
rect 525 299 555 499
rect 940 299 970 499
<< ndiff >>
rect 58 167 110 179
rect 58 133 66 167
rect 100 133 110 167
rect 58 99 110 133
rect 58 65 66 99
rect 100 65 110 99
rect 58 49 110 65
rect 140 167 192 179
rect 140 133 150 167
rect 184 133 192 167
rect 140 99 192 133
rect 140 65 150 99
rect 184 65 192 99
rect 140 49 192 65
rect 473 167 525 179
rect 473 133 481 167
rect 515 133 525 167
rect 473 99 525 133
rect 473 65 481 99
rect 515 65 525 99
rect 473 49 525 65
rect 555 167 607 179
rect 555 133 565 167
rect 599 133 607 167
rect 555 99 607 133
rect 555 65 565 99
rect 599 65 607 99
rect 555 49 607 65
rect 888 167 940 179
rect 888 133 896 167
rect 930 133 940 167
rect 888 99 940 133
rect 888 65 896 99
rect 930 65 940 99
rect 888 49 940 65
rect 970 167 1022 179
rect 970 133 980 167
rect 1014 133 1022 167
rect 970 99 1022 133
rect 970 65 980 99
rect 1014 65 1022 99
rect 970 49 1022 65
<< pdiff >>
rect 58 487 110 499
rect 58 453 66 487
rect 100 453 110 487
rect 58 419 110 453
rect 58 385 66 419
rect 100 385 110 419
rect 58 351 110 385
rect 58 317 66 351
rect 100 317 110 351
rect 58 299 110 317
rect 140 487 192 499
rect 140 453 150 487
rect 184 453 192 487
rect 473 487 525 499
rect 140 419 192 453
rect 140 385 150 419
rect 184 385 192 419
rect 140 351 192 385
rect 140 317 150 351
rect 184 317 192 351
rect 473 453 481 487
rect 515 453 525 487
rect 473 419 525 453
rect 473 385 481 419
rect 515 385 525 419
rect 473 351 525 385
rect 140 299 192 317
rect 473 317 481 351
rect 515 317 525 351
rect 473 299 525 317
rect 555 487 607 499
rect 555 453 565 487
rect 599 453 607 487
rect 888 487 940 499
rect 555 419 607 453
rect 555 385 565 419
rect 599 385 607 419
rect 555 351 607 385
rect 555 317 565 351
rect 599 317 607 351
rect 888 453 896 487
rect 930 453 940 487
rect 888 419 940 453
rect 888 385 896 419
rect 930 385 940 419
rect 888 351 940 385
rect 555 299 607 317
rect 888 317 896 351
rect 930 317 940 351
rect 888 299 940 317
rect 970 487 1022 499
rect 970 453 980 487
rect 1014 453 1022 487
rect 970 419 1022 453
rect 970 385 980 419
rect 1014 385 1022 419
rect 970 351 1022 385
rect 970 317 980 351
rect 1014 317 1022 351
rect 970 299 1022 317
<< ndiffc >>
rect 66 133 100 167
rect 66 65 100 99
rect 150 133 184 167
rect 150 65 184 99
rect 481 133 515 167
rect 481 65 515 99
rect 565 133 599 167
rect 565 65 599 99
rect 896 133 930 167
rect 896 65 930 99
rect 980 133 1014 167
rect 980 65 1014 99
<< pdiffc >>
rect 66 453 100 487
rect 66 385 100 419
rect 66 317 100 351
rect 150 453 184 487
rect 150 385 184 419
rect 150 317 184 351
rect 481 453 515 487
rect 481 385 515 419
rect 481 317 515 351
rect 565 453 599 487
rect 565 385 599 419
rect 565 317 599 351
rect 896 453 930 487
rect 896 385 930 419
rect 896 317 930 351
rect 980 453 1014 487
rect 980 385 1014 419
rect 980 317 1014 351
<< psubdiff >>
rect -74 162 4 192
rect -74 83 -61 162
rect -9 83 4 162
rect -74 57 4 83
rect 341 162 419 192
rect 341 83 354 162
rect 406 83 419 162
rect 341 57 419 83
rect 756 162 834 192
rect 756 83 769 162
rect 821 83 834 162
rect 756 57 834 83
<< nsubdiff >>
rect -74 450 4 481
rect -74 387 -61 450
rect -7 387 4 450
rect -74 338 4 387
rect 341 450 419 481
rect 341 387 354 450
rect 408 387 419 450
rect 341 338 419 387
rect 756 450 834 481
rect 756 387 769 450
rect 823 387 834 450
rect 756 338 834 387
<< psubdiffcont >>
rect -61 83 -9 162
rect 354 83 406 162
rect 769 83 821 162
<< nsubdiffcont >>
rect -61 387 -7 450
rect 354 387 408 450
rect 769 387 823 450
<< poly >>
rect 110 499 140 525
rect 525 499 555 525
rect 940 499 970 525
rect 110 267 140 299
rect 525 267 555 299
rect 940 267 970 299
rect 54 251 140 267
rect 54 217 70 251
rect 104 217 140 251
rect 54 201 140 217
rect 469 251 555 267
rect 469 217 485 251
rect 519 217 555 251
rect 469 201 555 217
rect 884 251 970 267
rect 884 217 900 251
rect 934 217 970 251
rect 884 201 970 217
rect 110 179 140 201
rect 525 179 555 201
rect 940 179 970 201
rect 110 23 140 49
rect 525 23 555 49
rect 940 23 970 49
<< polycont >>
rect 70 217 104 251
rect 485 217 519 251
rect 900 217 934 251
<< locali >>
rect -10 529 19 563
rect 53 529 111 563
rect 145 529 203 563
rect 237 529 266 563
rect 405 529 434 563
rect 468 529 526 563
rect 560 529 618 563
rect 652 529 681 563
rect 820 529 849 563
rect 883 529 941 563
rect 975 529 1033 563
rect 1067 529 1096 563
rect 58 487 100 529
rect 58 468 66 487
rect -74 453 66 468
rect -74 450 100 453
rect -74 387 -61 450
rect -7 419 100 450
rect -7 387 66 419
rect -74 385 66 387
rect -74 361 100 385
rect 58 351 100 361
rect 58 317 66 351
rect 58 301 100 317
rect 134 487 200 495
rect 134 453 150 487
rect 184 453 200 487
rect 473 487 515 529
rect 473 468 481 487
rect 134 419 200 453
rect 134 385 150 419
rect 184 385 200 419
rect 134 351 200 385
rect 341 453 481 468
rect 341 450 515 453
rect 341 387 354 450
rect 408 419 515 450
rect 408 387 481 419
rect 341 385 481 387
rect 341 361 515 385
rect 134 317 150 351
rect 184 317 200 351
rect 134 299 200 317
rect 473 351 515 361
rect 473 317 481 351
rect 473 301 515 317
rect 549 487 615 495
rect 549 453 565 487
rect 599 453 615 487
rect 888 487 930 529
rect 888 468 896 487
rect 549 419 615 453
rect 549 385 565 419
rect 599 385 615 419
rect 549 351 615 385
rect 756 453 896 468
rect 756 450 930 453
rect 756 387 769 450
rect 823 419 930 450
rect 823 387 896 419
rect 756 385 896 387
rect 756 361 930 385
rect 549 317 565 351
rect 599 317 615 351
rect 549 299 615 317
rect 888 351 930 361
rect 888 317 896 351
rect 888 301 930 317
rect 964 487 1030 495
rect 964 453 980 487
rect 1014 453 1030 487
rect 964 419 1030 453
rect 964 385 980 419
rect 1014 385 1030 419
rect 964 351 1030 385
rect 964 317 980 351
rect 1014 317 1030 351
rect 964 299 1030 317
rect -324 265 -68 298
rect 154 265 200 299
rect 569 265 615 299
rect 984 265 1030 299
rect -324 251 120 265
rect -324 218 70 251
rect -324 -80 -176 218
rect -111 217 70 218
rect 104 217 120 251
rect 154 251 535 265
rect 154 217 485 251
rect 519 217 535 251
rect 569 251 950 265
rect 569 217 900 251
rect 934 217 950 251
rect 984 264 1134 265
rect 984 218 1296 264
rect 984 217 1134 218
rect -74 167 100 183
rect 154 179 200 217
rect -74 162 66 167
rect -74 83 -61 162
rect -9 133 66 162
rect -9 99 100 133
rect -9 83 66 99
rect -74 65 66 83
rect -74 64 100 65
rect 54 19 100 64
rect 134 167 200 179
rect 134 133 150 167
rect 184 133 200 167
rect 134 99 200 133
rect 134 65 150 99
rect 184 65 200 99
rect 134 53 200 65
rect 341 167 515 183
rect 569 179 615 217
rect 341 162 481 167
rect 341 83 354 162
rect 406 133 481 162
rect 406 99 515 133
rect 406 83 481 99
rect 341 65 481 83
rect 341 64 515 65
rect 469 19 515 64
rect 549 167 615 179
rect 549 133 565 167
rect 599 133 615 167
rect 549 99 615 133
rect 549 65 565 99
rect 599 65 615 99
rect 549 53 615 65
rect 756 167 930 183
rect 984 179 1030 217
rect 756 162 896 167
rect 756 83 769 162
rect 821 133 896 162
rect 821 99 930 133
rect 821 83 896 99
rect 756 65 896 83
rect 756 64 930 65
rect 884 19 930 64
rect 964 167 1030 179
rect 964 133 980 167
rect 1014 133 1030 167
rect 964 99 1030 133
rect 964 65 980 99
rect 1014 65 1030 99
rect 964 53 1030 65
rect -10 -15 19 19
rect 53 -15 111 19
rect 145 -15 203 19
rect 237 -15 266 19
rect 405 -15 434 19
rect 468 -15 526 19
rect 560 -15 618 19
rect 652 -15 681 19
rect 820 -15 849 19
rect 883 -15 941 19
rect 975 -15 1033 19
rect 1067 -15 1096 19
rect 1230 -80 1294 218
rect -324 -176 1294 -80
<< viali >>
rect 19 529 53 563
rect 111 529 145 563
rect 203 529 237 563
rect 434 529 468 563
rect 526 529 560 563
rect 618 529 652 563
rect 849 529 883 563
rect 941 529 975 563
rect 1033 529 1067 563
rect 19 -15 53 19
rect 111 -15 145 19
rect 203 -15 237 19
rect 434 -15 468 19
rect 526 -15 560 19
rect 618 -15 652 19
rect 849 -15 883 19
rect 941 -15 975 19
rect 1033 -15 1067 19
<< metal1 >>
rect 662 594 896 680
rect -111 563 1134 594
rect -111 529 19 563
rect 53 529 111 563
rect 145 529 203 563
rect 237 529 434 563
rect 468 529 526 563
rect 560 529 618 563
rect 652 529 849 563
rect 883 529 941 563
rect 975 529 1033 563
rect 1067 529 1134 563
rect -111 498 1134 529
rect 662 50 722 84
rect -111 19 1134 50
rect -111 -15 19 19
rect 53 -15 111 19
rect 145 -15 203 19
rect 237 -15 434 19
rect 468 -15 526 19
rect 560 -15 618 19
rect 652 -15 849 19
rect 883 -15 941 19
rect 975 -15 1033 19
rect 1067 -15 1134 19
rect -111 -46 1134 -15
<< labels >>
flabel locali 1150 224 1252 256 1 FreeSans 800 0 0 0 out
port 1 n
flabel space 694 226 796 258 1 FreeSans 800 0 0 0 n2
flabel space 280 230 382 262 1 FreeSans 800 0 0 0 n1
flabel metal1 662 588 896 680 1 FreeSans 800 0 0 0 VDD
port 2 n
flabel metal1 662 40 722 84 1 FreeSans 800 0 0 0 GND
port 3 n
flabel locali 62 223 96 257 0 FreeSans 340 0 0 0 inv1_0[0]/A
flabel locali 154 291 188 325 0 FreeSans 340 0 0 0 inv1_0[0]/Y
flabel metal1 19 529 53 563 0 FreeSans 200 0 0 0 inv1_0[0]/VPWR
flabel metal1 19 -15 53 19 0 FreeSans 200 0 0 0 inv1_0[0]/VGND
rlabel comment -10 2 -10 2 4 inv1_0[0]/inv_1
flabel locali 477 223 511 257 0 FreeSans 340 0 0 0 inv1_0[1]/A
flabel locali 569 291 603 325 0 FreeSans 340 0 0 0 inv1_0[1]/Y
flabel metal1 434 529 468 563 0 FreeSans 200 0 0 0 inv1_0[1]/VPWR
flabel metal1 434 -15 468 19 0 FreeSans 200 0 0 0 inv1_0[1]/VGND
rlabel comment 405 2 405 2 4 inv1_0[1]/inv_1
flabel locali 892 223 926 257 0 FreeSans 340 0 0 0 inv1_0[2]/A
flabel locali 984 291 1018 325 0 FreeSans 340 0 0 0 inv1_0[2]/Y
flabel metal1 849 529 883 563 0 FreeSans 200 0 0 0 inv1_0[2]/VPWR
flabel metal1 849 -15 883 19 0 FreeSans 200 0 0 0 inv1_0[2]/VGND
rlabel comment 820 2 820 2 4 inv1_0[2]/inv_1
<< end >>
