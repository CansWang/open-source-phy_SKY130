* NGSPICE file created from pad_con_psub.ext - technology: sky130A

.subckt sky130_fd_io__pad_esd VSUBS m4_960_20297# m5_1334_20520# m5_1354_20528#
R0 m4_960_20297# m5_1354_20528# sky130_fd_pr__res_generic_m5 w=2.5296e+08u l=100000u
C0 m5_1334_20520# m4_960_20297# 1.87fF
C1 m5_1354_20528# m4_960_20297# 23.34fF
C2 m5_1354_20528# VSUBS 24.78fF
C3 m5_1334_20520# VSUBS -0.02fF
C4 m4_960_20297# VSUBS 34.99fF
.ends

.subckt sky130_fd_io__com_busses_esd sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_bus_hookup_0/VSSA
+ sky130_fd_io__com_bus_hookup_0/VDDIO_Q sky130_fd_io__com_bus_hookup_0/VSSIO_Q sky130_fd_io__com_bus_hookup_0/VSSIO
+ sky130_fd_io__com_bus_hookup_0/VSWITCH sky130_fd_io__com_bus_hookup_0/AMUXBUS_B
+ sky130_fd_io__com_bus_hookup_0/VCCD sky130_fd_io__com_bus_hookup_0/VDDIO sky130_fd_io__com_bus_hookup_0/AMUXBUS_A
+ sky130_fd_io__pad_esd_0/m5_1334_20520# sky130_fd_io__com_bus_hookup_0/VSSD sky130_fd_io__pad_esd_0/m5_1354_20528#
+ sky130_fd_io__pad_esd_0/m4_960_20297# sky130_fd_io__com_bus_hookup_0/VCCHIB
Xsky130_fd_io__pad_esd_0 VSUBS sky130_fd_io__pad_esd_0/m4_960_20297# sky130_fd_io__pad_esd_0/m5_1334_20520#
+ sky130_fd_io__pad_esd_0/m5_1354_20528# sky130_fd_io__pad_esd
C0 sky130_fd_io__com_bus_hookup_0/VSSD sky130_fd_io__com_bus_hookup_0/VSSA 18.85fF
C1 sky130_fd_io__com_bus_hookup_0/AMUXBUS_A sky130_fd_io__com_bus_hookup_0/VSSA 54.96fF
C2 sky130_fd_io__com_bus_hookup_0/VSSIO_Q sky130_fd_io__com_bus_hookup_0/VDDIO_Q 9.54fF
C3 sky130_fd_io__com_bus_hookup_0/VCCHIB sky130_fd_io__com_bus_hookup_0/VCCD 6.60fF
C4 sky130_fd_io__com_bus_hookup_0/VSSIO_Q sky130_fd_io__com_bus_hookup_0/VSSA 9.30fF
C5 sky130_fd_io__com_bus_hookup_0/VDDIO sky130_fd_io__com_bus_hookup_0/VSSIO 9.54fF
C6 sky130_fd_io__com_bus_hookup_0/VSSA sky130_fd_io__com_bus_hookup_0/VSWITCH 4.15fF
C7 sky130_fd_io__com_bus_hookup_0/AMUXBUS_A sky130_fd_io__com_bus_hookup_0/AMUXBUS_B 2.82fF
C8 sky130_fd_io__com_bus_hookup_0/VSSIO sky130_fd_io__com_bus_hookup_0/VSWITCH 5.74fF
C9 sky130_fd_io__com_bus_hookup_0/VSSA sky130_fd_io__com_bus_hookup_0/AMUXBUS_B 53.92fF
C10 sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_bus_hookup_0/VCCD 9.54fF
C11 sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_bus_hookup_0/VDDIO 9.54fF
C12 sky130_fd_io__com_bus_hookup_0/VDDIO sky130_fd_io__com_bus_hookup_0/VDDIO_Q 9.30fF
C13 sky130_fd_io__pad_esd_0/m5_1354_20528# VSUBS 24.78fF
C14 sky130_fd_io__pad_esd_0/m5_1334_20520# VSUBS -0.02fF
C15 sky130_fd_io__pad_esd_0/m4_960_20297# VSUBS 34.99fF
C16 sky130_fd_io__com_bus_hookup_0/VCCHIB VSUBS 22.19fF
C17 sky130_fd_io__com_bus_hookup_0/VCCD VSUBS 4.99fF
C18 sky130_fd_io__com_bus_hookup_0/VDDA VSUBS 2.34fF
C19 sky130_fd_io__com_bus_hookup_0/VDDIO VSUBS 70.89fF
C20 sky130_fd_io__com_bus_hookup_0/VSSIO VSUBS 72.21fF
C21 sky130_fd_io__com_bus_hookup_0/VSWITCH VSUBS 2.44fF
C22 sky130_fd_io__com_bus_hookup_0/VSSA VSUBS 40.31fF
C23 sky130_fd_io__com_bus_hookup_0/VSSD VSUBS 19.12fF
C24 sky130_fd_io__com_bus_hookup_0/AMUXBUS_B VSUBS 11.34fF
C25 sky130_fd_io__com_bus_hookup_0/AMUXBUS_A VSUBS 11.34fF
C26 sky130_fd_io__com_bus_hookup_0/VSSIO_Q VSUBS 4.60fF
C27 sky130_fd_io__com_bus_hookup_0/VDDIO_Q VSUBS 4.66fF
.ends

.subckt sky130_fd_io__simple_pad_and_busses VSUBS sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCHIB sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO
+ m3_99_16575# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1354_20528# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD
+ w_818_9944# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD
Xsky130_fd_io__com_busses_esd_0 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1334_20520#
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1354_20528#
+ m3_99_16575# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCHIB
+ sky130_fd_io__com_busses_esd
C0 m3_99_16575# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO 66.40fF
C1 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA 17.81fF
C2 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCHIB sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD 6.60fF
C3 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA 4.15fF
C4 m3_99_16575# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A 9.95fF
C5 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA 18.85fF
C6 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A 0.46fF
C7 m3_99_16575# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO 8.93fF
C8 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q 9.54fF
C9 m3_99_16575# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B 9.95fF
C10 m3_99_16575# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q 12.05fF
C11 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO 2.54fF
C12 m3_99_16575# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCHIB 9.48fF
C13 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B 2.52fF
C14 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q 0.80fF
C15 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA 54.96fF
C16 m3_99_16575# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD 10.55fF
C17 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD 9.54fF
C18 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO 5.74fF
C19 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA 53.92fF
C20 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA 9.30fF
C21 sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1354_20528# m3_99_16575# -63.86fF
C22 m3_99_16575# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q 15.51fF
C23 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO 9.54fF
C24 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA 0.80fF
C25 m3_99_16575# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA 19.12fF
C26 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A 2.82fF
C27 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH m3_99_16575# 7.24fF
C28 m3_99_16575# sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1334_20520# -1.24fF
C29 m3_99_16575# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD 9.93fF
C30 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA 4.25fF
C31 m3_99_16575# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA 23.82fF
C32 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD 5.84fF
C33 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA 4.78fF
C34 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO 9.30fF
C35 sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1354_20528# VSUBS 24.78fF
C36 sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1334_20520# VSUBS -0.02fF
C37 m3_99_16575# VSUBS -54.33fF
C38 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCHIB VSUBS 22.19fF
C39 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD VSUBS 4.99fF
C40 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA VSUBS -87.59fF
C41 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO VSUBS 70.89fF
C42 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO VSUBS 72.21fF
C43 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH VSUBS 2.44fF
C44 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA VSUBS 40.31fF
C45 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD VSUBS 19.12fF
C46 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B VSUBS 11.34fF
C47 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A VSUBS 11.34fF
C48 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q VSUBS 4.60fF
C49 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q VSUBS 4.66fF
.ends

.subckt test VSSA AMUXBUS_B VCCHIB sky130_fd_io__simple_pad_and_busses_0/VSUBS VCCD
+ P_PAD VSSIO_Q VDDIO_Q AMUXBUS_A P_CORE VSSIO VDDA VSSD VDDIO VSWITCH
Xsky130_fd_io__simple_pad_and_busses_0 sky130_fd_io__simple_pad_and_busses_0/VSUBS
+ VSSA VSWITCH AMUXBUS_A VDDA VSSIO VCCHIB VDDIO P_CORE VSSIO_Q P_PAD AMUXBUS_B VDDIO_Q
+ VSSD sky130_fd_io__simple_pad_and_busses_0/VSUBS VCCD sky130_fd_io__simple_pad_and_busses
C0 VSSA VSSD 18.71fF
C1 VDDIO VDDIO_Q 9.30fF
C2 VSSA VSSIO_Q 9.30fF
C3 VSWITCH VSSIO 5.74fF
C4 VDDIO VSSIO 9.54fF
C5 VSSA AMUXBUS_B 53.71fF
C6 VCCHIB VCCD 6.47fF
C7 VSSA VSWITCH 4.02fF
C8 VDDA VDDIO 9.54fF
C9 VDDIO_Q VSSIO_Q 9.54fF
C10 VSSA AMUXBUS_A 54.63fF
C11 VDDA VCCD 9.54fF
C12 AMUXBUS_A AMUXBUS_B 2.82fF
C13 P_PAD sky130_fd_io__simple_pad_and_busses_0/VSUBS 23.94fF
C14 sky130_fd_io__simple_pad_and_busses_0/sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1334_20520# sky130_fd_io__simple_pad_and_busses_0/VSUBS -0.02fF
C15 P_CORE sky130_fd_io__simple_pad_and_busses_0/VSUBS -53.74fF
C16 VCCHIB sky130_fd_io__simple_pad_and_busses_0/VSUBS 24.12fF
C17 VCCD sky130_fd_io__simple_pad_and_busses_0/VSUBS 4.81fF
C18 VDDA sky130_fd_io__simple_pad_and_busses_0/VSUBS -87.99fF
C19 VDDIO sky130_fd_io__simple_pad_and_busses_0/VSUBS 66.88fF
C20 VSSIO sky130_fd_io__simple_pad_and_busses_0/VSUBS 69.78fF
C21 VSWITCH sky130_fd_io__simple_pad_and_busses_0/VSUBS 3.72fF
C22 VSSA sky130_fd_io__simple_pad_and_busses_0/VSUBS 40.32fF
C23 VSSD sky130_fd_io__simple_pad_and_busses_0/VSUBS 19.60fF
C24 AMUXBUS_B sky130_fd_io__simple_pad_and_busses_0/VSUBS 11.05fF
C25 AMUXBUS_A sky130_fd_io__simple_pad_and_busses_0/VSUBS 11.96fF
C26 VSSIO_Q sky130_fd_io__simple_pad_and_busses_0/VSUBS 6.20fF
C27 VDDIO_Q sky130_fd_io__simple_pad_and_busses_0/VSUBS 4.06fF
.ends

.subckt pad_con_psub in out VDD GND
Xtest_0 GND GND VDD GND VDD out GND VDD GND in GND VDD GND VDD GND test
C0 out GND 22.02fF
C1 test_0/sky130_fd_io__simple_pad_and_busses_0/sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1334_20520# GND -0.02fF
C2 in GND -52.72fF
C3 VDD GND 6.53fF
.ends

