* NGSPICE file created from sky130_ef_io__analog_pad.ext - technology: sky130A

.subckt sky130_fd_io__pad_esd VSUBS m4_960_20297# m5_1354_20528#
R0 m4_960_20297# m5_1354_20528# sky130_fd_pr__res_generic_m5 w=2.5284e+08u l=100000u
.ends

.subckt sky130_fd_io__com_busses_esd VSUBS sky130_fd_io__com_bus_hookup_0/VCCD sky130_fd_io__com_bus_hookup_0/VSWITCH
+ sky130_fd_io__com_bus_hookup_0/AMUXBUS_A sky130_fd_io__com_bus_hookup_0/VSSIO sky130_fd_io__com_bus_hookup_0/AMUXBUS_B
+ sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_bus_hookup_0/VDDIO sky130_fd_io__com_bus_hookup_0/VSSIO_Q
+ sky130_fd_io__pad_esd_0/m5_1354_20528# sky130_fd_io__pad_esd_0/m4_960_20297# sky130_fd_io__com_bus_hookup_0/VDDIO_Q
+ sky130_fd_io__com_bus_hookup_0/VSSA sky130_fd_io__com_bus_hookup_0/VSSD sky130_fd_io__com_bus_hookup_0/VCCHIB
Xsky130_fd_io__pad_esd_0 VSUBS sky130_fd_io__pad_esd_0/m4_960_20297# sky130_fd_io__pad_esd_0/m5_1354_20528#
+ sky130_fd_io__pad_esd
.ends

.subckt sky130_fd_io__simple_pad_and_busses VSUBS sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCHIB sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO
+ m3_99_16575# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1354_20528#
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD
+ w_818_9944# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD
Xsky130_fd_io__com_busses_esd_0 VSUBS sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1354_20528#
+ m3_99_16575# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCHIB sky130_fd_io__com_busses_esd
.ends

.subckt sky130_ef_io__analog_pad P_CORE VSSA VSSD AMUXBUS_B AMUXBUS_A VDDIO_Q VDDIO
+ VSWITCH VSSIO VDDA VCCD VCCHIB VSSIO_Q P_PAD
Xsky130_fd_io__simple_pad_and_busses_0 sky130_fd_io__simple_pad_and_busses_0/VSUBS
+ VSWITCH VDDA VSSIO VCCHIB VDDIO P_CORE VSSIO_Q AMUXBUS_A P_PAD AMUXBUS_B VSSA VDDIO_Q
+ VSSD sky130_fd_io__simple_pad_and_busses_0/VSUBS VCCD sky130_fd_io__simple_pad_and_busses
.ends


* Wrapper for pad goes here
.subckt pad_example in out VDD GND

Xanalog_pad in GND GND GND GND VDD VDD GND GND VDD VDD VDD GND out sky130_ef_io__analog_pad

.ends




