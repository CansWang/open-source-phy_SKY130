* NGSPICE file created from pad_test.ext - technology: sky130A

.subckt sky130_fd_io__com_busses_esd VSUBS sky130_fd_io__com_bus_hookup_0/VCCD sky130_fd_io__com_bus_hookup_0/VSWITCH
+ sky130_fd_io__pad_esd_0/sky130_fd_pr__padplhp__example_559591418080_0/m5_n540_766#
+ sky130_fd_io__com_bus_hookup_0/AMUXBUS_A sky130_fd_io__com_bus_hookup_0/VSSIO sky130_fd_io__com_bus_hookup_0/AMUXBUS_B
+ sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_bus_hookup_0/VDDIO sky130_fd_io__com_bus_hookup_0/VSSIO_Q
+ sky130_fd_io__com_bus_hookup_0/VDDIO_Q sky130_fd_io__com_bus_hookup_0/VSSA sky130_fd_io__com_bus_hookup_0/VSSD
+ sky130_fd_io__com_bus_hookup_0/VCCHIB
.ends

.subckt sky130_fd_io__simple_pad_and_busses VSUBS sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCHIB sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO
+ m3_99_16575# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD
Xsky130_fd_io__com_busses_esd_0 VSUBS sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH m3_99_16575#
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCHIB
+ sky130_fd_io__com_busses_esd
.ends

.subckt test VSSA VSUBS VSSD VCCHIB VSSIO_Q VCCD P_PAD VDDIO_Q VSSIO VDDA VDDIO VSWITCH
Xsky130_fd_io__simple_pad_and_busses_0 VSUBS VSWITCH VDDA VSSIO VCCHIB VDDIO P_PAD
+ VSSIO_Q AMUXBUS_A AMUXBUS_B VSSA VDDIO_Q VSSD VCCD sky130_fd_io__simple_pad_and_busses
.ends

.subckt pad_test out VDD GND
Xtest_0 GND VSUBS GND VDD GND VDD out VDD GND VDD VDD GND test
.ends

