* Include SKY130 libraries
.lib "/afs/ir.stanford.edu/class/ee272/skywater-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice" tt

.ic V(1)=0 V(sw1)=3.3
*+V(in_dut)=0


* NAND2_8 
.subckt sky130_fd_sc_hs__nand2_8 A B VGND VNB VPB VPWR Y
X0 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X3 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X9 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X14 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X16 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X20 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X22 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__nand2_4 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X8 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X9 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X11 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
X0 Y A1 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 a_114_85# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VGND a_1030_268# a_475_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR a_1030_268# a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X4 a_475_85# A0 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_114_85# S VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_116_368# a_1030_268# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X7 Y A1 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X8 a_475_85# a_1030_268# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 Y A0 a_475_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_478_368# S VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X11 VPWR S a_478_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X12 a_475_85# A0 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_1030_268# S VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X14 Y A1 a_114_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 Y A0 a_475_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_478_368# A0 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X17 a_116_368# a_1030_268# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X18 a_116_368# A1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X19 Y A1 a_114_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 Y A0 a_478_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X21 a_116_368# A1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X22 a_114_85# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 a_475_85# a_1030_268# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 VPWR S a_478_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X25 VGND S a_114_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 VGND S a_1030_268# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 VGND a_1030_268# a_475_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 a_478_368# S VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X29 VPWR S a_1030_268# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X30 VGND S a_114_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 Y A0 a_478_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X32 a_478_368# A0 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X33 VPWR a_1030_268# a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X34 a_114_85# S VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends


.subckt sky130_fd_sc_hs__inv_4 A VGND VNB VPB VPWR Y
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

.subckt cc cin en VDD VGND
X0 cin en VGND VGND VDD VDD z1 sky130_fd_sc_hs__nand2_4 m=1
.ends

.subckt cc1 cin en VDD VGND
X1 VGND cin en VGND VGND VDD VDD z1 sky130_fd_sc_hs__mux2i_4 m=1
.ends


.subckt fc cin en VGND VGND VDD VDD VGND
* inv input buffer
X1 cin VGND VGND VDD VDD Y1 sky130_fd_sc_hs__inv_4
X0 Y1 en VGND VGND VDD VDD z1 sky130_fd_sc_hs__nand2_8
.ends

* Switching signal
Vpump sw1 0 DC 0 PWL(0 1.8 2NS 0 10NS 0)
Vdut sw2 0 DC 0 PWL(0 0 3NS 1.8 10NS 1.8)
Vc out 0 DC 1.8V
Vsup VDD 0 1.8v

* XC bias generation
* XINV1 in_dut 0 0 VDD VDD 2 sky130_fd_sc_hs__inv_4
* XINV2 2 0 0 VDD VDD in_dut sky130_fd_sc_hs__inv_4


.model switch_charge sw vt=1.65 vh=0.01 ron=100 roff=1e12

*Reference cap 
C1 1 0 10fF
R1 1 0 1e10

*DUT cap cell
XC1 in_dut VDD VDD 0 cc
*XC1 in_dut VDD VDD 0 cc1
*XFC1 in_dut VDD 0 0 VDD VDD 0 fc

spump out 1 sw1 0 switch_charge ON
sdut 1 in_dut sw2 0 switch_charge OFF


* specify simulation duration, with "uic"
* indicating "use initial conditions"
.tran 10e-12 12e-09 1e-09 uic CHGTOL=1e-16 TRTOL=1

* ngspice control commands
.control
save all
run
write
display
*plot V(in_dut)
.endc

* end of the testbench


.end

