magic
tech sky130A
magscale 1 2
timestamp 1620043962
<< error_s >>
rect 5548 39000 5557 39003
rect 9506 39000 9518 39006
rect 5542 38994 9524 39000
rect 5536 38988 9530 38994
rect 5536 38982 5554 38988
rect 5548 37779 5554 38982
rect 5539 37776 5554 37779
rect 9512 38982 9530 38988
rect 9512 37779 9524 38982
rect 9512 37776 9527 37779
rect 5539 37770 9527 37776
rect 5548 37761 5557 37770
rect 9506 37764 9524 37770
rect 9506 37758 9518 37764
<< dnwell >>
rect 1518 10962 1754 11198
rect 1068 9932 1304 10168
rect 1552 10006 1788 10242
rect 2024 9970 2260 10206
rect 2510 9930 2746 10166
rect 2882 9938 3118 10174
rect 3262 9952 3498 10188
<< psubdiff >>
rect 5548 38760 9518 38994
rect 5548 37954 6084 38760
rect 9016 37954 9518 38760
rect 5548 37770 9518 37954
<< psubdiffcont >>
rect 6084 37954 9016 38760
<< viali >>
rect 5548 38760 9518 38994
rect 5548 37954 6084 38760
rect 6084 37954 9016 38760
rect 9016 37954 9518 38760
rect 5548 37770 9518 37954
<< via1 >>
rect 5548 37770 9518 38994
<< via2 >>
rect 5548 37770 9518 38994
<< metal3 >>
rect 5878 -1304 9090 132
<< via3 >>
rect 5548 37770 9518 38994
<< via4 >>
rect 176 10814 412 11050
rect 1052 10840 1288 11076
rect 1518 10962 1754 11198
rect 1068 9932 1304 10168
rect 1552 10006 1788 10242
rect 2024 9970 2260 10206
rect 2510 9930 2746 10166
rect 2882 9938 3118 10174
rect 3262 9952 3498 10188
<< metal5 >>
rect 5816 39430 9028 40866
rect -2060 38198 -934 38252
rect -2060 35840 3518 38198
rect -2060 12516 -934 35840
rect 5764 30240 8976 31676
rect 15844 15456 17212 15564
rect 13902 14426 17212 15456
rect 0 13488 854 14260
rect -2816 11050 936 12516
rect -2816 10814 176 11050
rect 412 10814 936 11050
rect -2816 7962 936 10814
rect -2816 7780 1082 7962
rect -2816 5194 936 7780
rect 15844 4766 17212 14426
rect 770 638 2694 4698
rect 14412 4084 17212 4766
rect 14412 4070 17078 4084
use test  test_0
timestamp 1620043962
transform 1 0 0 0 1 0
box 0 0 15000 40000
<< labels >>
flabel metal5 770 638 2694 4698 1 FreeSans 6400 0 0 0 VDD
port 3 n
flabel metal3 5878 -1304 9090 132 1 FreeSans 6400 0 0 0 in
port 1 n
flabel metal5 5764 30240 8976 31676 1 FreeSans 6400 0 0 0 out
port 2 n
flabel metal5 5816 39430 9028 40866 1 FreeSans 6400 0 0 0 GND
port 4 n
<< end >>
