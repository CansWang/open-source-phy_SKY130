magic
tech sky130A
magscale 1 2
timestamp 1619862920
<< checkpaint >>
rect -1285 -960 1385 1561
<< labels >>
flabel comment s 125 300 125 300 0 FreeSans 300 0 0 0 D
flabel comment s -25 300 -25 300 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 1789530
string GDS_START 1788762
<< end >>
