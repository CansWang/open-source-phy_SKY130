magic
tech sky130A
magscale 1 2
timestamp 1619862920
<< checkpaint >>
rect -1260 -1253 16260 40860
<< metal3 >>
tri 12210 18591 12211 18592 se
rect 12211 18591 14932 18592
rect 119 18527 135 18591
rect 199 18527 217 18591
rect 281 18527 299 18591
rect 363 18527 381 18591
rect 445 18527 463 18591
rect 527 18527 545 18591
rect 609 18527 627 18591
rect 691 18527 709 18591
rect 773 18527 791 18591
rect 855 18527 873 18591
rect 937 18527 955 18591
rect 1019 18527 1037 18591
rect 1101 18527 1119 18591
rect 1183 18527 1201 18591
rect 1265 18527 1283 18591
rect 1347 18527 1365 18591
rect 1429 18527 1447 18591
rect 1511 18527 1529 18591
rect 1593 18527 1611 18591
rect 1675 18527 1693 18591
rect 1757 18527 1775 18591
rect 1839 18527 1857 18591
rect 1921 18527 1939 18591
rect 2003 18527 2021 18591
rect 2085 18527 2103 18591
rect 2167 18527 2185 18591
rect 2249 18527 2267 18591
rect 2331 18527 2349 18591
rect 2413 18527 2431 18591
rect 2495 18527 2513 18591
rect 2577 18527 2594 18591
rect 2658 18527 2675 18591
rect 2739 18527 2756 18591
rect 2820 18527 2841 18591
rect 119 18509 2841 18527
rect 119 18445 135 18509
rect 199 18445 217 18509
rect 281 18445 299 18509
rect 363 18445 381 18509
rect 445 18445 463 18509
rect 527 18445 545 18509
rect 609 18445 627 18509
rect 691 18445 709 18509
rect 773 18445 791 18509
rect 855 18445 873 18509
rect 937 18445 955 18509
rect 1019 18445 1037 18509
rect 1101 18445 1119 18509
rect 1183 18445 1201 18509
rect 1265 18445 1283 18509
rect 1347 18445 1365 18509
rect 1429 18445 1447 18509
rect 1511 18445 1529 18509
rect 1593 18445 1611 18509
rect 1675 18445 1693 18509
rect 1757 18445 1775 18509
rect 1839 18445 1857 18509
rect 1921 18445 1939 18509
rect 2003 18445 2021 18509
rect 2085 18445 2103 18509
rect 2167 18445 2185 18509
rect 2249 18445 2267 18509
rect 2331 18445 2349 18509
rect 2413 18445 2431 18509
rect 2495 18445 2513 18509
rect 2577 18445 2594 18509
rect 2658 18445 2675 18509
rect 2739 18445 2756 18509
rect 2820 18445 2841 18509
rect 119 18427 2841 18445
rect 119 18363 135 18427
rect 199 18363 217 18427
rect 281 18363 299 18427
rect 363 18363 381 18427
rect 445 18363 463 18427
rect 527 18363 545 18427
rect 609 18363 627 18427
rect 691 18363 709 18427
rect 773 18363 791 18427
rect 855 18363 873 18427
rect 937 18363 955 18427
rect 1019 18363 1037 18427
rect 1101 18363 1119 18427
rect 1183 18363 1201 18427
rect 1265 18363 1283 18427
rect 1347 18363 1365 18427
rect 1429 18363 1447 18427
rect 1511 18363 1529 18427
rect 1593 18363 1611 18427
rect 1675 18363 1693 18427
rect 1757 18363 1775 18427
rect 1839 18363 1857 18427
rect 1921 18363 1939 18427
rect 2003 18363 2021 18427
rect 2085 18363 2103 18427
rect 2167 18363 2185 18427
rect 2249 18363 2267 18427
rect 2331 18363 2349 18427
rect 2413 18363 2431 18427
rect 2495 18363 2513 18427
rect 2577 18363 2594 18427
rect 2658 18363 2675 18427
rect 2739 18363 2756 18427
rect 2820 18363 2841 18427
rect 119 18347 2841 18363
tri 2841 18347 3085 18591 sw
tri 11966 18347 12210 18591 se
rect 12210 18527 12231 18591
rect 12295 18527 12312 18591
rect 12376 18527 12393 18591
rect 12457 18527 12474 18591
rect 12538 18527 12556 18591
rect 12620 18527 12638 18591
rect 12702 18527 12720 18591
rect 12784 18527 12802 18591
rect 12866 18527 12884 18591
rect 12948 18527 12966 18591
rect 13030 18527 13048 18591
rect 13112 18527 13130 18591
rect 13194 18527 13212 18591
rect 13276 18527 13294 18591
rect 13358 18527 13376 18591
rect 13440 18527 13458 18591
rect 13522 18527 13540 18591
rect 13604 18527 13622 18591
rect 13686 18527 13704 18591
rect 13768 18527 13786 18591
rect 13850 18527 13868 18591
rect 13932 18527 13950 18591
rect 14014 18527 14032 18591
rect 14096 18527 14114 18591
rect 14178 18527 14196 18591
rect 14260 18527 14278 18591
rect 14342 18527 14360 18591
rect 14424 18527 14442 18591
rect 14506 18527 14524 18591
rect 14588 18527 14606 18591
rect 14670 18527 14688 18591
rect 14752 18527 14770 18591
rect 14834 18527 14852 18591
rect 14916 18527 14932 18591
rect 12210 18509 14932 18527
rect 12210 18445 12231 18509
rect 12295 18445 12312 18509
rect 12376 18445 12393 18509
rect 12457 18445 12474 18509
rect 12538 18445 12556 18509
rect 12620 18445 12638 18509
rect 12702 18445 12720 18509
rect 12784 18445 12802 18509
rect 12866 18445 12884 18509
rect 12948 18445 12966 18509
rect 13030 18445 13048 18509
rect 13112 18445 13130 18509
rect 13194 18445 13212 18509
rect 13276 18445 13294 18509
rect 13358 18445 13376 18509
rect 13440 18445 13458 18509
rect 13522 18445 13540 18509
rect 13604 18445 13622 18509
rect 13686 18445 13704 18509
rect 13768 18445 13786 18509
rect 13850 18445 13868 18509
rect 13932 18445 13950 18509
rect 14014 18445 14032 18509
rect 14096 18445 14114 18509
rect 14178 18445 14196 18509
rect 14260 18445 14278 18509
rect 14342 18445 14360 18509
rect 14424 18445 14442 18509
rect 14506 18445 14524 18509
rect 14588 18445 14606 18509
rect 14670 18445 14688 18509
rect 14752 18445 14770 18509
rect 14834 18445 14852 18509
rect 14916 18445 14932 18509
rect 12210 18427 14932 18445
rect 12210 18363 12231 18427
rect 12295 18363 12312 18427
rect 12376 18363 12393 18427
rect 12457 18363 12474 18427
rect 12538 18363 12556 18427
rect 12620 18363 12638 18427
rect 12702 18363 12720 18427
rect 12784 18363 12802 18427
rect 12866 18363 12884 18427
rect 12948 18363 12966 18427
rect 13030 18363 13048 18427
rect 13112 18363 13130 18427
rect 13194 18363 13212 18427
rect 13276 18363 13294 18427
rect 13358 18363 13376 18427
rect 13440 18363 13458 18427
rect 13522 18363 13540 18427
rect 13604 18363 13622 18427
rect 13686 18363 13704 18427
rect 13768 18363 13786 18427
rect 13850 18363 13868 18427
rect 13932 18363 13950 18427
rect 14014 18363 14032 18427
rect 14096 18363 14114 18427
rect 14178 18363 14196 18427
rect 14260 18363 14278 18427
rect 14342 18363 14360 18427
rect 14424 18363 14442 18427
rect 14506 18363 14524 18427
rect 14588 18363 14606 18427
rect 14670 18363 14688 18427
rect 14752 18363 14770 18427
rect 14834 18363 14852 18427
rect 14916 18363 14932 18427
rect 12210 18347 14932 18363
rect 119 18345 3085 18347
rect 119 18281 135 18345
rect 199 18281 217 18345
rect 281 18281 299 18345
rect 363 18281 381 18345
rect 445 18281 463 18345
rect 527 18281 545 18345
rect 609 18281 627 18345
rect 691 18281 709 18345
rect 773 18281 791 18345
rect 855 18281 873 18345
rect 937 18281 955 18345
rect 1019 18281 1037 18345
rect 1101 18281 1119 18345
rect 1183 18281 1201 18345
rect 1265 18281 1283 18345
rect 1347 18281 1365 18345
rect 1429 18281 1447 18345
rect 1511 18281 1529 18345
rect 1593 18281 1611 18345
rect 1675 18281 1693 18345
rect 1757 18281 1775 18345
rect 1839 18281 1857 18345
rect 1921 18281 1939 18345
rect 2003 18281 2021 18345
rect 2085 18281 2103 18345
rect 2167 18281 2185 18345
rect 2249 18281 2267 18345
rect 2331 18281 2349 18345
rect 2413 18281 2431 18345
rect 2495 18281 2513 18345
rect 2577 18281 2594 18345
rect 2658 18281 2675 18345
rect 2739 18281 2756 18345
rect 2820 18341 3085 18345
rect 2820 18281 2852 18341
rect 119 18277 2852 18281
rect 2916 18277 3008 18341
rect 3072 18277 3085 18341
rect 119 18263 3085 18277
rect 119 18199 135 18263
rect 199 18199 217 18263
rect 281 18199 299 18263
rect 363 18199 381 18263
rect 445 18199 463 18263
rect 527 18199 545 18263
rect 609 18199 627 18263
rect 691 18199 709 18263
rect 773 18199 791 18263
rect 855 18199 873 18263
rect 937 18199 955 18263
rect 1019 18199 1037 18263
rect 1101 18199 1119 18263
rect 1183 18199 1201 18263
rect 1265 18199 1283 18263
rect 1347 18199 1365 18263
rect 1429 18199 1447 18263
rect 1511 18199 1529 18263
rect 1593 18199 1611 18263
rect 1675 18199 1693 18263
rect 1757 18199 1775 18263
rect 1839 18199 1857 18263
rect 1921 18199 1939 18263
rect 2003 18199 2021 18263
rect 2085 18199 2103 18263
rect 2167 18199 2185 18263
rect 2249 18199 2267 18263
rect 2331 18199 2349 18263
rect 2413 18199 2431 18263
rect 2495 18199 2513 18263
rect 2577 18199 2594 18263
rect 2658 18199 2675 18263
rect 2739 18199 2756 18263
rect 2820 18255 3085 18263
rect 2820 18199 2852 18255
rect 119 18191 2852 18199
rect 2916 18191 3008 18255
rect 3072 18191 3085 18255
rect 119 18185 3085 18191
tri 3085 18185 3247 18347 sw
tri 11804 18185 11966 18347 se
rect 11966 18345 14932 18347
rect 11966 18341 12231 18345
rect 11966 18277 11979 18341
rect 12043 18277 12135 18341
rect 12199 18281 12231 18341
rect 12295 18281 12312 18345
rect 12376 18281 12393 18345
rect 12457 18281 12474 18345
rect 12538 18281 12556 18345
rect 12620 18281 12638 18345
rect 12702 18281 12720 18345
rect 12784 18281 12802 18345
rect 12866 18281 12884 18345
rect 12948 18281 12966 18345
rect 13030 18281 13048 18345
rect 13112 18281 13130 18345
rect 13194 18281 13212 18345
rect 13276 18281 13294 18345
rect 13358 18281 13376 18345
rect 13440 18281 13458 18345
rect 13522 18281 13540 18345
rect 13604 18281 13622 18345
rect 13686 18281 13704 18345
rect 13768 18281 13786 18345
rect 13850 18281 13868 18345
rect 13932 18281 13950 18345
rect 14014 18281 14032 18345
rect 14096 18281 14114 18345
rect 14178 18281 14196 18345
rect 14260 18281 14278 18345
rect 14342 18281 14360 18345
rect 14424 18281 14442 18345
rect 14506 18281 14524 18345
rect 14588 18281 14606 18345
rect 14670 18281 14688 18345
rect 14752 18281 14770 18345
rect 14834 18281 14852 18345
rect 14916 18281 14932 18345
rect 12199 18277 14932 18281
rect 11966 18263 14932 18277
rect 11966 18255 12231 18263
rect 11966 18191 11979 18255
rect 12043 18191 12135 18255
rect 12199 18199 12231 18255
rect 12295 18199 12312 18263
rect 12376 18199 12393 18263
rect 12457 18199 12474 18263
rect 12538 18199 12556 18263
rect 12620 18199 12638 18263
rect 12702 18199 12720 18263
rect 12784 18199 12802 18263
rect 12866 18199 12884 18263
rect 12948 18199 12966 18263
rect 13030 18199 13048 18263
rect 13112 18199 13130 18263
rect 13194 18199 13212 18263
rect 13276 18199 13294 18263
rect 13358 18199 13376 18263
rect 13440 18199 13458 18263
rect 13522 18199 13540 18263
rect 13604 18199 13622 18263
rect 13686 18199 13704 18263
rect 13768 18199 13786 18263
rect 13850 18199 13868 18263
rect 13932 18199 13950 18263
rect 14014 18199 14032 18263
rect 14096 18199 14114 18263
rect 14178 18199 14196 18263
rect 14260 18199 14278 18263
rect 14342 18199 14360 18263
rect 14424 18199 14442 18263
rect 14506 18199 14524 18263
rect 14588 18199 14606 18263
rect 14670 18199 14688 18263
rect 14752 18199 14770 18263
rect 14834 18199 14852 18263
rect 14916 18199 14932 18263
rect 12199 18191 14932 18199
rect 11966 18185 14932 18191
rect 119 18181 3247 18185
rect 119 18117 135 18181
rect 199 18117 217 18181
rect 281 18117 299 18181
rect 363 18117 381 18181
rect 445 18117 463 18181
rect 527 18117 545 18181
rect 609 18117 627 18181
rect 691 18117 709 18181
rect 773 18117 791 18181
rect 855 18117 873 18181
rect 937 18117 955 18181
rect 1019 18117 1037 18181
rect 1101 18117 1119 18181
rect 1183 18117 1201 18181
rect 1265 18117 1283 18181
rect 1347 18117 1365 18181
rect 1429 18117 1447 18181
rect 1511 18117 1529 18181
rect 1593 18117 1611 18181
rect 1675 18117 1693 18181
rect 1757 18117 1775 18181
rect 1839 18117 1857 18181
rect 1921 18117 1939 18181
rect 2003 18117 2021 18181
rect 2085 18117 2103 18181
rect 2167 18117 2185 18181
rect 2249 18117 2267 18181
rect 2331 18117 2349 18181
rect 2413 18117 2431 18181
rect 2495 18117 2513 18181
rect 2577 18117 2594 18181
rect 2658 18117 2675 18181
rect 2739 18117 2756 18181
rect 2820 18169 3247 18181
tri 3247 18169 3263 18185 sw
tri 11788 18169 11804 18185 se
rect 11804 18181 14932 18185
rect 11804 18169 12231 18181
rect 2820 18163 3263 18169
rect 2820 18117 2856 18163
rect 119 18099 2856 18117
rect 2920 18099 2938 18163
rect 3002 18099 3020 18163
rect 3084 18099 3102 18163
rect 3166 18099 3184 18163
rect 3248 18099 3263 18163
rect 119 18035 135 18099
rect 199 18035 217 18099
rect 281 18035 299 18099
rect 363 18035 381 18099
rect 445 18035 463 18099
rect 527 18035 545 18099
rect 609 18035 627 18099
rect 691 18035 709 18099
rect 773 18035 791 18099
rect 855 18035 873 18099
rect 937 18035 955 18099
rect 1019 18035 1037 18099
rect 1101 18035 1119 18099
rect 1183 18035 1201 18099
rect 1265 18035 1283 18099
rect 1347 18035 1365 18099
rect 1429 18035 1447 18099
rect 1511 18035 1529 18099
rect 1593 18035 1611 18099
rect 1675 18035 1693 18099
rect 1757 18035 1775 18099
rect 1839 18035 1857 18099
rect 1921 18035 1939 18099
rect 2003 18035 2021 18099
rect 2085 18035 2103 18099
rect 2167 18035 2185 18099
rect 2249 18035 2267 18099
rect 2331 18035 2349 18099
rect 2413 18035 2431 18099
rect 2495 18035 2513 18099
rect 2577 18035 2594 18099
rect 2658 18035 2675 18099
rect 2739 18035 2756 18099
rect 2820 18077 3263 18099
rect 2820 18035 2856 18077
rect 119 18017 2856 18035
rect 119 17953 135 18017
rect 199 17953 217 18017
rect 281 17953 299 18017
rect 363 17953 381 18017
rect 445 17953 463 18017
rect 527 17953 545 18017
rect 609 17953 627 18017
rect 691 17953 709 18017
rect 773 17953 791 18017
rect 855 17953 873 18017
rect 937 17953 955 18017
rect 1019 17953 1037 18017
rect 1101 17953 1119 18017
rect 1183 17953 1201 18017
rect 1265 17953 1283 18017
rect 1347 17953 1365 18017
rect 1429 17953 1447 18017
rect 1511 17953 1529 18017
rect 1593 17953 1611 18017
rect 1675 17953 1693 18017
rect 1757 17953 1775 18017
rect 1839 17953 1857 18017
rect 1921 17953 1939 18017
rect 2003 17953 2021 18017
rect 2085 17953 2103 18017
rect 2167 17953 2185 18017
rect 2249 17953 2267 18017
rect 2331 17953 2349 18017
rect 2413 17953 2431 18017
rect 2495 17953 2513 18017
rect 2577 17953 2594 18017
rect 2658 17953 2675 18017
rect 2739 17953 2756 18017
rect 2820 18013 2856 18017
rect 2920 18013 2938 18077
rect 3002 18013 3020 18077
rect 3084 18013 3102 18077
rect 3166 18013 3184 18077
rect 3248 18013 3263 18077
rect 2820 17991 3263 18013
rect 2820 17953 2856 17991
rect 119 17935 2856 17953
rect 119 17871 135 17935
rect 199 17871 217 17935
rect 281 17871 299 17935
rect 363 17871 381 17935
rect 445 17871 463 17935
rect 527 17871 545 17935
rect 609 17871 627 17935
rect 691 17871 709 17935
rect 773 17871 791 17935
rect 855 17871 873 17935
rect 937 17871 955 17935
rect 1019 17871 1037 17935
rect 1101 17871 1119 17935
rect 1183 17871 1201 17935
rect 1265 17871 1283 17935
rect 1347 17871 1365 17935
rect 1429 17871 1447 17935
rect 1511 17871 1529 17935
rect 1593 17871 1611 17935
rect 1675 17871 1693 17935
rect 1757 17871 1775 17935
rect 1839 17871 1857 17935
rect 1921 17871 1939 17935
rect 2003 17871 2021 17935
rect 2085 17871 2103 17935
rect 2167 17871 2185 17935
rect 2249 17871 2267 17935
rect 2331 17871 2349 17935
rect 2413 17871 2431 17935
rect 2495 17871 2513 17935
rect 2577 17871 2594 17935
rect 2658 17871 2675 17935
rect 2739 17871 2756 17935
rect 2820 17927 2856 17935
rect 2920 17927 2938 17991
rect 3002 17927 3020 17991
rect 3084 17927 3102 17991
rect 3166 17927 3184 17991
rect 3248 17927 3263 17991
rect 2820 17911 3263 17927
tri 3263 17911 3521 18169 sw
tri 11530 17911 11788 18169 se
rect 11788 18163 12231 18169
rect 11788 18099 11803 18163
rect 11867 18099 11885 18163
rect 11949 18099 11967 18163
rect 12031 18099 12049 18163
rect 12113 18099 12131 18163
rect 12195 18117 12231 18163
rect 12295 18117 12312 18181
rect 12376 18117 12393 18181
rect 12457 18117 12474 18181
rect 12538 18117 12556 18181
rect 12620 18117 12638 18181
rect 12702 18117 12720 18181
rect 12784 18117 12802 18181
rect 12866 18117 12884 18181
rect 12948 18117 12966 18181
rect 13030 18117 13048 18181
rect 13112 18117 13130 18181
rect 13194 18117 13212 18181
rect 13276 18117 13294 18181
rect 13358 18117 13376 18181
rect 13440 18117 13458 18181
rect 13522 18117 13540 18181
rect 13604 18117 13622 18181
rect 13686 18117 13704 18181
rect 13768 18117 13786 18181
rect 13850 18117 13868 18181
rect 13932 18117 13950 18181
rect 14014 18117 14032 18181
rect 14096 18117 14114 18181
rect 14178 18117 14196 18181
rect 14260 18117 14278 18181
rect 14342 18117 14360 18181
rect 14424 18117 14442 18181
rect 14506 18117 14524 18181
rect 14588 18117 14606 18181
rect 14670 18117 14688 18181
rect 14752 18117 14770 18181
rect 14834 18117 14852 18181
rect 14916 18117 14932 18181
rect 12195 18099 14932 18117
rect 11788 18077 12231 18099
rect 11788 18013 11803 18077
rect 11867 18013 11885 18077
rect 11949 18013 11967 18077
rect 12031 18013 12049 18077
rect 12113 18013 12131 18077
rect 12195 18035 12231 18077
rect 12295 18035 12312 18099
rect 12376 18035 12393 18099
rect 12457 18035 12474 18099
rect 12538 18035 12556 18099
rect 12620 18035 12638 18099
rect 12702 18035 12720 18099
rect 12784 18035 12802 18099
rect 12866 18035 12884 18099
rect 12948 18035 12966 18099
rect 13030 18035 13048 18099
rect 13112 18035 13130 18099
rect 13194 18035 13212 18099
rect 13276 18035 13294 18099
rect 13358 18035 13376 18099
rect 13440 18035 13458 18099
rect 13522 18035 13540 18099
rect 13604 18035 13622 18099
rect 13686 18035 13704 18099
rect 13768 18035 13786 18099
rect 13850 18035 13868 18099
rect 13932 18035 13950 18099
rect 14014 18035 14032 18099
rect 14096 18035 14114 18099
rect 14178 18035 14196 18099
rect 14260 18035 14278 18099
rect 14342 18035 14360 18099
rect 14424 18035 14442 18099
rect 14506 18035 14524 18099
rect 14588 18035 14606 18099
rect 14670 18035 14688 18099
rect 14752 18035 14770 18099
rect 14834 18035 14852 18099
rect 14916 18035 14932 18099
rect 12195 18017 14932 18035
rect 12195 18013 12231 18017
rect 11788 17991 12231 18013
rect 11788 17927 11803 17991
rect 11867 17927 11885 17991
rect 11949 17927 11967 17991
rect 12031 17927 12049 17991
rect 12113 17927 12131 17991
rect 12195 17953 12231 17991
rect 12295 17953 12312 18017
rect 12376 17953 12393 18017
rect 12457 17953 12474 18017
rect 12538 17953 12556 18017
rect 12620 17953 12638 18017
rect 12702 17953 12720 18017
rect 12784 17953 12802 18017
rect 12866 17953 12884 18017
rect 12948 17953 12966 18017
rect 13030 17953 13048 18017
rect 13112 17953 13130 18017
rect 13194 17953 13212 18017
rect 13276 17953 13294 18017
rect 13358 17953 13376 18017
rect 13440 17953 13458 18017
rect 13522 17953 13540 18017
rect 13604 17953 13622 18017
rect 13686 17953 13704 18017
rect 13768 17953 13786 18017
rect 13850 17953 13868 18017
rect 13932 17953 13950 18017
rect 14014 17953 14032 18017
rect 14096 17953 14114 18017
rect 14178 17953 14196 18017
rect 14260 17953 14278 18017
rect 14342 17953 14360 18017
rect 14424 17953 14442 18017
rect 14506 17953 14524 18017
rect 14588 17953 14606 18017
rect 14670 17953 14688 18017
rect 14752 17953 14770 18017
rect 14834 17953 14852 18017
rect 14916 17953 14932 18017
rect 12195 17935 14932 17953
rect 12195 17927 12231 17935
rect 11788 17911 12231 17927
rect 2820 17905 3521 17911
rect 2820 17871 2856 17905
rect 119 17853 2856 17871
rect 119 17789 135 17853
rect 199 17789 217 17853
rect 281 17789 299 17853
rect 363 17789 381 17853
rect 445 17789 463 17853
rect 527 17789 545 17853
rect 609 17789 627 17853
rect 691 17789 709 17853
rect 773 17789 791 17853
rect 855 17789 873 17853
rect 937 17789 955 17853
rect 1019 17789 1037 17853
rect 1101 17789 1119 17853
rect 1183 17789 1201 17853
rect 1265 17789 1283 17853
rect 1347 17789 1365 17853
rect 1429 17789 1447 17853
rect 1511 17789 1529 17853
rect 1593 17789 1611 17853
rect 1675 17789 1693 17853
rect 1757 17789 1775 17853
rect 1839 17789 1857 17853
rect 1921 17789 1939 17853
rect 2003 17789 2021 17853
rect 2085 17789 2103 17853
rect 2167 17789 2185 17853
rect 2249 17789 2267 17853
rect 2331 17789 2349 17853
rect 2413 17789 2431 17853
rect 2495 17789 2513 17853
rect 2577 17789 2594 17853
rect 2658 17789 2675 17853
rect 2739 17789 2756 17853
rect 2820 17841 2856 17853
rect 2920 17841 2938 17905
rect 3002 17841 3020 17905
rect 3084 17841 3102 17905
rect 3166 17841 3184 17905
rect 3248 17841 3284 17905
rect 3348 17841 3440 17905
rect 3504 17841 3521 17905
rect 2820 17821 3521 17841
rect 2820 17819 3284 17821
rect 2820 17789 2856 17819
rect 119 17771 2856 17789
rect 119 17707 135 17771
rect 199 17707 217 17771
rect 281 17707 299 17771
rect 363 17707 381 17771
rect 445 17707 463 17771
rect 527 17707 545 17771
rect 609 17707 627 17771
rect 691 17707 709 17771
rect 773 17707 791 17771
rect 855 17707 873 17771
rect 937 17707 955 17771
rect 1019 17707 1037 17771
rect 1101 17707 1119 17771
rect 1183 17707 1201 17771
rect 1265 17707 1283 17771
rect 1347 17707 1365 17771
rect 1429 17707 1447 17771
rect 1511 17707 1529 17771
rect 1593 17707 1611 17771
rect 1675 17707 1693 17771
rect 1757 17707 1775 17771
rect 1839 17707 1857 17771
rect 1921 17707 1939 17771
rect 2003 17707 2021 17771
rect 2085 17707 2103 17771
rect 2167 17707 2185 17771
rect 2249 17707 2267 17771
rect 2331 17707 2349 17771
rect 2413 17707 2431 17771
rect 2495 17707 2513 17771
rect 2577 17707 2594 17771
rect 2658 17707 2675 17771
rect 2739 17707 2756 17771
rect 2820 17755 2856 17771
rect 2920 17755 2938 17819
rect 3002 17755 3020 17819
rect 3084 17755 3102 17819
rect 3166 17755 3184 17819
rect 3248 17757 3284 17819
rect 3348 17757 3440 17821
rect 3504 17757 3521 17821
rect 3248 17755 3521 17757
rect 2820 17738 3521 17755
rect 2820 17734 3284 17738
rect 2820 17707 2856 17734
rect 119 17689 2856 17707
rect 119 17625 135 17689
rect 199 17625 217 17689
rect 281 17625 299 17689
rect 363 17625 381 17689
rect 445 17625 463 17689
rect 527 17625 545 17689
rect 609 17625 627 17689
rect 691 17625 709 17689
rect 773 17625 791 17689
rect 855 17625 873 17689
rect 937 17625 955 17689
rect 1019 17625 1037 17689
rect 1101 17625 1119 17689
rect 1183 17625 1201 17689
rect 1265 17625 1283 17689
rect 1347 17625 1365 17689
rect 1429 17625 1447 17689
rect 1511 17625 1529 17689
rect 1593 17625 1611 17689
rect 1675 17625 1693 17689
rect 1757 17625 1775 17689
rect 1839 17625 1857 17689
rect 1921 17625 1939 17689
rect 2003 17625 2021 17689
rect 2085 17625 2103 17689
rect 2167 17625 2185 17689
rect 2249 17625 2267 17689
rect 2331 17625 2349 17689
rect 2413 17625 2431 17689
rect 2495 17625 2513 17689
rect 2577 17625 2594 17689
rect 2658 17625 2675 17689
rect 2739 17625 2756 17689
rect 2820 17670 2856 17689
rect 2920 17670 2938 17734
rect 3002 17670 3020 17734
rect 3084 17670 3102 17734
rect 3166 17670 3184 17734
rect 3248 17674 3284 17734
rect 3348 17674 3440 17738
rect 3504 17674 3521 17738
rect 3248 17670 3521 17674
rect 2820 17668 3521 17670
tri 3521 17668 3764 17911 sw
tri 11287 17668 11530 17911 se
rect 11530 17905 12231 17911
rect 11530 17841 11547 17905
rect 11611 17841 11703 17905
rect 11767 17841 11803 17905
rect 11867 17841 11885 17905
rect 11949 17841 11967 17905
rect 12031 17841 12049 17905
rect 12113 17841 12131 17905
rect 12195 17871 12231 17905
rect 12295 17871 12312 17935
rect 12376 17871 12393 17935
rect 12457 17871 12474 17935
rect 12538 17871 12556 17935
rect 12620 17871 12638 17935
rect 12702 17871 12720 17935
rect 12784 17871 12802 17935
rect 12866 17871 12884 17935
rect 12948 17871 12966 17935
rect 13030 17871 13048 17935
rect 13112 17871 13130 17935
rect 13194 17871 13212 17935
rect 13276 17871 13294 17935
rect 13358 17871 13376 17935
rect 13440 17871 13458 17935
rect 13522 17871 13540 17935
rect 13604 17871 13622 17935
rect 13686 17871 13704 17935
rect 13768 17871 13786 17935
rect 13850 17871 13868 17935
rect 13932 17871 13950 17935
rect 14014 17871 14032 17935
rect 14096 17871 14114 17935
rect 14178 17871 14196 17935
rect 14260 17871 14278 17935
rect 14342 17871 14360 17935
rect 14424 17871 14442 17935
rect 14506 17871 14524 17935
rect 14588 17871 14606 17935
rect 14670 17871 14688 17935
rect 14752 17871 14770 17935
rect 14834 17871 14852 17935
rect 14916 17871 14932 17935
rect 12195 17853 14932 17871
rect 12195 17841 12231 17853
rect 11530 17821 12231 17841
rect 11530 17757 11547 17821
rect 11611 17757 11703 17821
rect 11767 17819 12231 17821
rect 11767 17757 11803 17819
rect 11530 17755 11803 17757
rect 11867 17755 11885 17819
rect 11949 17755 11967 17819
rect 12031 17755 12049 17819
rect 12113 17755 12131 17819
rect 12195 17789 12231 17819
rect 12295 17789 12312 17853
rect 12376 17789 12393 17853
rect 12457 17789 12474 17853
rect 12538 17789 12556 17853
rect 12620 17789 12638 17853
rect 12702 17789 12720 17853
rect 12784 17789 12802 17853
rect 12866 17789 12884 17853
rect 12948 17789 12966 17853
rect 13030 17789 13048 17853
rect 13112 17789 13130 17853
rect 13194 17789 13212 17853
rect 13276 17789 13294 17853
rect 13358 17789 13376 17853
rect 13440 17789 13458 17853
rect 13522 17789 13540 17853
rect 13604 17789 13622 17853
rect 13686 17789 13704 17853
rect 13768 17789 13786 17853
rect 13850 17789 13868 17853
rect 13932 17789 13950 17853
rect 14014 17789 14032 17853
rect 14096 17789 14114 17853
rect 14178 17789 14196 17853
rect 14260 17789 14278 17853
rect 14342 17789 14360 17853
rect 14424 17789 14442 17853
rect 14506 17789 14524 17853
rect 14588 17789 14606 17853
rect 14670 17789 14688 17853
rect 14752 17789 14770 17853
rect 14834 17789 14852 17853
rect 14916 17789 14932 17853
rect 12195 17771 14932 17789
rect 12195 17755 12231 17771
rect 11530 17738 12231 17755
rect 11530 17674 11547 17738
rect 11611 17674 11703 17738
rect 11767 17734 12231 17738
rect 11767 17674 11803 17734
rect 11530 17670 11803 17674
rect 11867 17670 11885 17734
rect 11949 17670 11967 17734
rect 12031 17670 12049 17734
rect 12113 17670 12131 17734
rect 12195 17707 12231 17734
rect 12295 17707 12312 17771
rect 12376 17707 12393 17771
rect 12457 17707 12474 17771
rect 12538 17707 12556 17771
rect 12620 17707 12638 17771
rect 12702 17707 12720 17771
rect 12784 17707 12802 17771
rect 12866 17707 12884 17771
rect 12948 17707 12966 17771
rect 13030 17707 13048 17771
rect 13112 17707 13130 17771
rect 13194 17707 13212 17771
rect 13276 17707 13294 17771
rect 13358 17707 13376 17771
rect 13440 17707 13458 17771
rect 13522 17707 13540 17771
rect 13604 17707 13622 17771
rect 13686 17707 13704 17771
rect 13768 17707 13786 17771
rect 13850 17707 13868 17771
rect 13932 17707 13950 17771
rect 14014 17707 14032 17771
rect 14096 17707 14114 17771
rect 14178 17707 14196 17771
rect 14260 17707 14278 17771
rect 14342 17707 14360 17771
rect 14424 17707 14442 17771
rect 14506 17707 14524 17771
rect 14588 17707 14606 17771
rect 14670 17707 14688 17771
rect 14752 17707 14770 17771
rect 14834 17707 14852 17771
rect 14916 17707 14932 17771
rect 12195 17689 14932 17707
rect 12195 17670 12231 17689
rect 11530 17668 12231 17670
rect 2820 17664 3764 17668
tri 3764 17664 3768 17668 sw
tri 11283 17664 11287 17668 se
rect 11287 17664 12231 17668
rect 2820 17633 3768 17664
tri 3768 17633 3799 17664 sw
tri 11252 17633 11283 17664 se
rect 11283 17633 12231 17664
rect 2820 17627 3799 17633
rect 2820 17625 2881 17627
rect 119 17607 2881 17625
rect 119 17543 135 17607
rect 199 17543 217 17607
rect 281 17543 299 17607
rect 363 17543 381 17607
rect 445 17543 463 17607
rect 527 17543 545 17607
rect 609 17543 627 17607
rect 691 17543 709 17607
rect 773 17543 791 17607
rect 855 17543 873 17607
rect 937 17543 955 17607
rect 1019 17543 1037 17607
rect 1101 17543 1119 17607
rect 1183 17543 1201 17607
rect 1265 17543 1283 17607
rect 1347 17543 1365 17607
rect 1429 17543 1447 17607
rect 1511 17543 1529 17607
rect 1593 17543 1611 17607
rect 1675 17543 1693 17607
rect 1757 17543 1775 17607
rect 1839 17543 1857 17607
rect 1921 17543 1939 17607
rect 2003 17543 2021 17607
rect 2085 17543 2103 17607
rect 2167 17543 2185 17607
rect 2249 17543 2267 17607
rect 2331 17543 2349 17607
rect 2413 17543 2431 17607
rect 2495 17543 2513 17607
rect 2577 17543 2594 17607
rect 2658 17543 2675 17607
rect 2739 17543 2756 17607
rect 2820 17563 2881 17607
rect 2945 17563 2963 17627
rect 3027 17563 3045 17627
rect 3109 17563 3127 17627
rect 3191 17563 3209 17627
rect 3273 17563 3291 17627
rect 3355 17563 3373 17627
rect 3437 17563 3455 17627
rect 3519 17563 3537 17627
rect 3601 17563 3619 17627
rect 3683 17563 3701 17627
rect 3765 17563 3799 17627
rect 2820 17546 3799 17563
rect 2820 17543 2881 17546
rect 119 17525 2881 17543
rect 119 17461 135 17525
rect 199 17461 217 17525
rect 281 17461 299 17525
rect 363 17461 381 17525
rect 445 17461 463 17525
rect 527 17461 545 17525
rect 609 17461 627 17525
rect 691 17461 709 17525
rect 773 17461 791 17525
rect 855 17461 873 17525
rect 937 17461 955 17525
rect 1019 17461 1037 17525
rect 1101 17461 1119 17525
rect 1183 17461 1201 17525
rect 1265 17461 1283 17525
rect 1347 17461 1365 17525
rect 1429 17461 1447 17525
rect 1511 17461 1529 17525
rect 1593 17461 1611 17525
rect 1675 17461 1693 17525
rect 1757 17461 1775 17525
rect 1839 17461 1857 17525
rect 1921 17461 1939 17525
rect 2003 17461 2021 17525
rect 2085 17461 2103 17525
rect 2167 17461 2185 17525
rect 2249 17461 2267 17525
rect 2331 17461 2349 17525
rect 2413 17461 2431 17525
rect 2495 17461 2513 17525
rect 2577 17461 2594 17525
rect 2658 17461 2675 17525
rect 2739 17461 2756 17525
rect 2820 17482 2881 17525
rect 2945 17482 2963 17546
rect 3027 17482 3045 17546
rect 3109 17482 3127 17546
rect 3191 17482 3209 17546
rect 3273 17482 3291 17546
rect 3355 17482 3373 17546
rect 3437 17482 3455 17546
rect 3519 17482 3537 17546
rect 3601 17482 3619 17546
rect 3683 17482 3701 17546
rect 3765 17482 3799 17546
rect 2820 17465 3799 17482
rect 2820 17461 2881 17465
rect 119 17443 2881 17461
rect 119 17379 135 17443
rect 199 17379 217 17443
rect 281 17379 299 17443
rect 363 17379 381 17443
rect 445 17379 463 17443
rect 527 17379 545 17443
rect 609 17379 627 17443
rect 691 17379 709 17443
rect 773 17379 791 17443
rect 855 17379 873 17443
rect 937 17379 955 17443
rect 1019 17379 1037 17443
rect 1101 17379 1119 17443
rect 1183 17379 1201 17443
rect 1265 17379 1283 17443
rect 1347 17379 1365 17443
rect 1429 17379 1447 17443
rect 1511 17379 1529 17443
rect 1593 17379 1611 17443
rect 1675 17379 1693 17443
rect 1757 17379 1775 17443
rect 1839 17379 1857 17443
rect 1921 17379 1939 17443
rect 2003 17379 2021 17443
rect 2085 17379 2103 17443
rect 2167 17379 2185 17443
rect 2249 17379 2267 17443
rect 2331 17379 2349 17443
rect 2413 17379 2431 17443
rect 2495 17379 2513 17443
rect 2577 17379 2594 17443
rect 2658 17379 2675 17443
rect 2739 17379 2756 17443
rect 2820 17401 2881 17443
rect 2945 17401 2963 17465
rect 3027 17401 3045 17465
rect 3109 17401 3127 17465
rect 3191 17401 3209 17465
rect 3273 17401 3291 17465
rect 3355 17401 3373 17465
rect 3437 17401 3455 17465
rect 3519 17401 3537 17465
rect 3601 17401 3619 17465
rect 3683 17401 3701 17465
rect 3765 17408 3799 17465
tri 3799 17408 4024 17633 sw
tri 11027 17408 11252 17633 se
rect 11252 17627 12231 17633
rect 11252 17563 11286 17627
rect 11350 17563 11368 17627
rect 11432 17563 11450 17627
rect 11514 17563 11532 17627
rect 11596 17563 11614 17627
rect 11678 17563 11696 17627
rect 11760 17563 11778 17627
rect 11842 17563 11860 17627
rect 11924 17563 11942 17627
rect 12006 17563 12024 17627
rect 12088 17563 12106 17627
rect 12170 17625 12231 17627
rect 12295 17625 12312 17689
rect 12376 17625 12393 17689
rect 12457 17625 12474 17689
rect 12538 17625 12556 17689
rect 12620 17625 12638 17689
rect 12702 17625 12720 17689
rect 12784 17625 12802 17689
rect 12866 17625 12884 17689
rect 12948 17625 12966 17689
rect 13030 17625 13048 17689
rect 13112 17625 13130 17689
rect 13194 17625 13212 17689
rect 13276 17625 13294 17689
rect 13358 17625 13376 17689
rect 13440 17625 13458 17689
rect 13522 17625 13540 17689
rect 13604 17625 13622 17689
rect 13686 17625 13704 17689
rect 13768 17625 13786 17689
rect 13850 17625 13868 17689
rect 13932 17625 13950 17689
rect 14014 17625 14032 17689
rect 14096 17625 14114 17689
rect 14178 17625 14196 17689
rect 14260 17625 14278 17689
rect 14342 17625 14360 17689
rect 14424 17625 14442 17689
rect 14506 17625 14524 17689
rect 14588 17625 14606 17689
rect 14670 17625 14688 17689
rect 14752 17625 14770 17689
rect 14834 17625 14852 17689
rect 14916 17625 14932 17689
rect 12170 17607 14932 17625
rect 12170 17563 12231 17607
rect 11252 17546 12231 17563
rect 11252 17482 11286 17546
rect 11350 17482 11368 17546
rect 11432 17482 11450 17546
rect 11514 17482 11532 17546
rect 11596 17482 11614 17546
rect 11678 17482 11696 17546
rect 11760 17482 11778 17546
rect 11842 17482 11860 17546
rect 11924 17482 11942 17546
rect 12006 17482 12024 17546
rect 12088 17482 12106 17546
rect 12170 17543 12231 17546
rect 12295 17543 12312 17607
rect 12376 17543 12393 17607
rect 12457 17543 12474 17607
rect 12538 17543 12556 17607
rect 12620 17543 12638 17607
rect 12702 17543 12720 17607
rect 12784 17543 12802 17607
rect 12866 17543 12884 17607
rect 12948 17543 12966 17607
rect 13030 17543 13048 17607
rect 13112 17543 13130 17607
rect 13194 17543 13212 17607
rect 13276 17543 13294 17607
rect 13358 17543 13376 17607
rect 13440 17543 13458 17607
rect 13522 17543 13540 17607
rect 13604 17543 13622 17607
rect 13686 17543 13704 17607
rect 13768 17543 13786 17607
rect 13850 17543 13868 17607
rect 13932 17543 13950 17607
rect 14014 17543 14032 17607
rect 14096 17543 14114 17607
rect 14178 17543 14196 17607
rect 14260 17543 14278 17607
rect 14342 17543 14360 17607
rect 14424 17543 14442 17607
rect 14506 17543 14524 17607
rect 14588 17543 14606 17607
rect 14670 17543 14688 17607
rect 14752 17543 14770 17607
rect 14834 17543 14852 17607
rect 14916 17543 14932 17607
rect 12170 17525 14932 17543
rect 12170 17482 12231 17525
rect 11252 17465 12231 17482
rect 11252 17408 11286 17465
rect 3765 17402 4024 17408
rect 3765 17401 3800 17402
rect 2820 17384 3800 17401
rect 2820 17379 2881 17384
rect 119 17361 2881 17379
rect 119 17297 135 17361
rect 199 17297 217 17361
rect 281 17297 299 17361
rect 363 17297 381 17361
rect 445 17297 463 17361
rect 527 17297 545 17361
rect 609 17297 627 17361
rect 691 17297 709 17361
rect 773 17297 791 17361
rect 855 17297 873 17361
rect 937 17297 955 17361
rect 1019 17297 1037 17361
rect 1101 17297 1119 17361
rect 1183 17297 1201 17361
rect 1265 17297 1283 17361
rect 1347 17297 1365 17361
rect 1429 17297 1447 17361
rect 1511 17297 1529 17361
rect 1593 17297 1611 17361
rect 1675 17297 1693 17361
rect 1757 17297 1775 17361
rect 1839 17297 1857 17361
rect 1921 17297 1939 17361
rect 2003 17297 2021 17361
rect 2085 17297 2103 17361
rect 2167 17297 2185 17361
rect 2249 17297 2267 17361
rect 2331 17297 2349 17361
rect 2413 17297 2431 17361
rect 2495 17297 2513 17361
rect 2577 17297 2594 17361
rect 2658 17297 2675 17361
rect 2739 17297 2756 17361
rect 2820 17320 2881 17361
rect 2945 17320 2963 17384
rect 3027 17320 3045 17384
rect 3109 17320 3127 17384
rect 3191 17320 3209 17384
rect 3273 17320 3291 17384
rect 3355 17320 3373 17384
rect 3437 17320 3455 17384
rect 3519 17320 3537 17384
rect 3601 17320 3619 17384
rect 3683 17320 3701 17384
rect 3765 17338 3800 17384
rect 3864 17338 3948 17402
rect 4012 17338 4024 17402
rect 3765 17320 4024 17338
rect 2820 17314 4024 17320
rect 2820 17303 3800 17314
rect 2820 17297 2881 17303
rect 119 17279 2881 17297
rect 119 17215 135 17279
rect 199 17215 217 17279
rect 281 17215 299 17279
rect 363 17215 381 17279
rect 445 17215 463 17279
rect 527 17215 545 17279
rect 609 17215 627 17279
rect 691 17215 709 17279
rect 773 17215 791 17279
rect 855 17215 873 17279
rect 937 17215 955 17279
rect 1019 17215 1037 17279
rect 1101 17215 1119 17279
rect 1183 17215 1201 17279
rect 1265 17215 1283 17279
rect 1347 17215 1365 17279
rect 1429 17215 1447 17279
rect 1511 17215 1529 17279
rect 1593 17215 1611 17279
rect 1675 17215 1693 17279
rect 1757 17215 1775 17279
rect 1839 17215 1857 17279
rect 1921 17215 1939 17279
rect 2003 17215 2021 17279
rect 2085 17215 2103 17279
rect 2167 17215 2185 17279
rect 2249 17215 2267 17279
rect 2331 17215 2349 17279
rect 2413 17215 2431 17279
rect 2495 17215 2513 17279
rect 2577 17215 2594 17279
rect 2658 17215 2675 17279
rect 2739 17215 2756 17279
rect 2820 17239 2881 17279
rect 2945 17239 2963 17303
rect 3027 17239 3045 17303
rect 3109 17239 3127 17303
rect 3191 17239 3209 17303
rect 3273 17239 3291 17303
rect 3355 17239 3373 17303
rect 3437 17239 3455 17303
rect 3519 17239 3537 17303
rect 3601 17239 3619 17303
rect 3683 17239 3701 17303
rect 3765 17250 3800 17303
rect 3864 17250 3948 17314
rect 4012 17250 4024 17314
rect 3765 17239 4024 17250
rect 2820 17227 4024 17239
rect 2820 17223 3800 17227
rect 2820 17215 2881 17223
rect 119 17197 2881 17215
rect 119 17133 135 17197
rect 199 17133 217 17197
rect 281 17133 299 17197
rect 363 17133 381 17197
rect 445 17133 463 17197
rect 527 17133 545 17197
rect 609 17133 627 17197
rect 691 17133 709 17197
rect 773 17133 791 17197
rect 855 17133 873 17197
rect 937 17133 955 17197
rect 1019 17133 1037 17197
rect 1101 17133 1119 17197
rect 1183 17133 1201 17197
rect 1265 17133 1283 17197
rect 1347 17133 1365 17197
rect 1429 17133 1447 17197
rect 1511 17133 1529 17197
rect 1593 17133 1611 17197
rect 1675 17133 1693 17197
rect 1757 17133 1775 17197
rect 1839 17133 1857 17197
rect 1921 17133 1939 17197
rect 2003 17133 2021 17197
rect 2085 17133 2103 17197
rect 2167 17133 2185 17197
rect 2249 17133 2267 17197
rect 2331 17133 2349 17197
rect 2413 17133 2431 17197
rect 2495 17133 2513 17197
rect 2577 17133 2594 17197
rect 2658 17133 2675 17197
rect 2739 17133 2756 17197
rect 2820 17159 2881 17197
rect 2945 17159 2963 17223
rect 3027 17159 3045 17223
rect 3109 17159 3127 17223
rect 3191 17159 3209 17223
rect 3273 17159 3291 17223
rect 3355 17159 3373 17223
rect 3437 17159 3455 17223
rect 3519 17159 3537 17223
rect 3601 17159 3619 17223
rect 3683 17159 3701 17223
rect 3765 17163 3800 17223
rect 3864 17163 3948 17227
rect 4012 17163 4024 17227
rect 3765 17159 4024 17163
rect 2820 17157 4024 17159
tri 4024 17157 4275 17408 sw
tri 10776 17157 11027 17408 se
rect 11027 17402 11286 17408
rect 11027 17338 11039 17402
rect 11103 17338 11187 17402
rect 11251 17401 11286 17402
rect 11350 17401 11368 17465
rect 11432 17401 11450 17465
rect 11514 17401 11532 17465
rect 11596 17401 11614 17465
rect 11678 17401 11696 17465
rect 11760 17401 11778 17465
rect 11842 17401 11860 17465
rect 11924 17401 11942 17465
rect 12006 17401 12024 17465
rect 12088 17401 12106 17465
rect 12170 17461 12231 17465
rect 12295 17461 12312 17525
rect 12376 17461 12393 17525
rect 12457 17461 12474 17525
rect 12538 17461 12556 17525
rect 12620 17461 12638 17525
rect 12702 17461 12720 17525
rect 12784 17461 12802 17525
rect 12866 17461 12884 17525
rect 12948 17461 12966 17525
rect 13030 17461 13048 17525
rect 13112 17461 13130 17525
rect 13194 17461 13212 17525
rect 13276 17461 13294 17525
rect 13358 17461 13376 17525
rect 13440 17461 13458 17525
rect 13522 17461 13540 17525
rect 13604 17461 13622 17525
rect 13686 17461 13704 17525
rect 13768 17461 13786 17525
rect 13850 17461 13868 17525
rect 13932 17461 13950 17525
rect 14014 17461 14032 17525
rect 14096 17461 14114 17525
rect 14178 17461 14196 17525
rect 14260 17461 14278 17525
rect 14342 17461 14360 17525
rect 14424 17461 14442 17525
rect 14506 17461 14524 17525
rect 14588 17461 14606 17525
rect 14670 17461 14688 17525
rect 14752 17461 14770 17525
rect 14834 17461 14852 17525
rect 14916 17461 14932 17525
rect 12170 17443 14932 17461
rect 12170 17401 12231 17443
rect 11251 17384 12231 17401
rect 11251 17338 11286 17384
rect 11027 17320 11286 17338
rect 11350 17320 11368 17384
rect 11432 17320 11450 17384
rect 11514 17320 11532 17384
rect 11596 17320 11614 17384
rect 11678 17320 11696 17384
rect 11760 17320 11778 17384
rect 11842 17320 11860 17384
rect 11924 17320 11942 17384
rect 12006 17320 12024 17384
rect 12088 17320 12106 17384
rect 12170 17379 12231 17384
rect 12295 17379 12312 17443
rect 12376 17379 12393 17443
rect 12457 17379 12474 17443
rect 12538 17379 12556 17443
rect 12620 17379 12638 17443
rect 12702 17379 12720 17443
rect 12784 17379 12802 17443
rect 12866 17379 12884 17443
rect 12948 17379 12966 17443
rect 13030 17379 13048 17443
rect 13112 17379 13130 17443
rect 13194 17379 13212 17443
rect 13276 17379 13294 17443
rect 13358 17379 13376 17443
rect 13440 17379 13458 17443
rect 13522 17379 13540 17443
rect 13604 17379 13622 17443
rect 13686 17379 13704 17443
rect 13768 17379 13786 17443
rect 13850 17379 13868 17443
rect 13932 17379 13950 17443
rect 14014 17379 14032 17443
rect 14096 17379 14114 17443
rect 14178 17379 14196 17443
rect 14260 17379 14278 17443
rect 14342 17379 14360 17443
rect 14424 17379 14442 17443
rect 14506 17379 14524 17443
rect 14588 17379 14606 17443
rect 14670 17379 14688 17443
rect 14752 17379 14770 17443
rect 14834 17379 14852 17443
rect 14916 17379 14932 17443
rect 12170 17361 14932 17379
rect 12170 17320 12231 17361
rect 11027 17314 12231 17320
rect 11027 17250 11039 17314
rect 11103 17250 11187 17314
rect 11251 17303 12231 17314
rect 11251 17250 11286 17303
rect 11027 17239 11286 17250
rect 11350 17239 11368 17303
rect 11432 17239 11450 17303
rect 11514 17239 11532 17303
rect 11596 17239 11614 17303
rect 11678 17239 11696 17303
rect 11760 17239 11778 17303
rect 11842 17239 11860 17303
rect 11924 17239 11942 17303
rect 12006 17239 12024 17303
rect 12088 17239 12106 17303
rect 12170 17297 12231 17303
rect 12295 17297 12312 17361
rect 12376 17297 12393 17361
rect 12457 17297 12474 17361
rect 12538 17297 12556 17361
rect 12620 17297 12638 17361
rect 12702 17297 12720 17361
rect 12784 17297 12802 17361
rect 12866 17297 12884 17361
rect 12948 17297 12966 17361
rect 13030 17297 13048 17361
rect 13112 17297 13130 17361
rect 13194 17297 13212 17361
rect 13276 17297 13294 17361
rect 13358 17297 13376 17361
rect 13440 17297 13458 17361
rect 13522 17297 13540 17361
rect 13604 17297 13622 17361
rect 13686 17297 13704 17361
rect 13768 17297 13786 17361
rect 13850 17297 13868 17361
rect 13932 17297 13950 17361
rect 14014 17297 14032 17361
rect 14096 17297 14114 17361
rect 14178 17297 14196 17361
rect 14260 17297 14278 17361
rect 14342 17297 14360 17361
rect 14424 17297 14442 17361
rect 14506 17297 14524 17361
rect 14588 17297 14606 17361
rect 14670 17297 14688 17361
rect 14752 17297 14770 17361
rect 14834 17297 14852 17361
rect 14916 17297 14932 17361
rect 12170 17279 14932 17297
rect 12170 17239 12231 17279
rect 11027 17227 12231 17239
rect 11027 17163 11039 17227
rect 11103 17163 11187 17227
rect 11251 17223 12231 17227
rect 11251 17163 11286 17223
rect 11027 17159 11286 17163
rect 11350 17159 11368 17223
rect 11432 17159 11450 17223
rect 11514 17159 11532 17223
rect 11596 17159 11614 17223
rect 11678 17159 11696 17223
rect 11760 17159 11778 17223
rect 11842 17159 11860 17223
rect 11924 17159 11942 17223
rect 12006 17159 12024 17223
rect 12088 17159 12106 17223
rect 12170 17215 12231 17223
rect 12295 17215 12312 17279
rect 12376 17215 12393 17279
rect 12457 17215 12474 17279
rect 12538 17215 12556 17279
rect 12620 17215 12638 17279
rect 12702 17215 12720 17279
rect 12784 17215 12802 17279
rect 12866 17215 12884 17279
rect 12948 17215 12966 17279
rect 13030 17215 13048 17279
rect 13112 17215 13130 17279
rect 13194 17215 13212 17279
rect 13276 17215 13294 17279
rect 13358 17215 13376 17279
rect 13440 17215 13458 17279
rect 13522 17215 13540 17279
rect 13604 17215 13622 17279
rect 13686 17215 13704 17279
rect 13768 17215 13786 17279
rect 13850 17215 13868 17279
rect 13932 17215 13950 17279
rect 14014 17215 14032 17279
rect 14096 17215 14114 17279
rect 14178 17215 14196 17279
rect 14260 17215 14278 17279
rect 14342 17215 14360 17279
rect 14424 17215 14442 17279
rect 14506 17215 14524 17279
rect 14588 17215 14606 17279
rect 14670 17215 14688 17279
rect 14752 17215 14770 17279
rect 14834 17215 14852 17279
rect 14916 17215 14932 17279
rect 12170 17197 14932 17215
rect 12170 17159 12231 17197
rect 11027 17157 12231 17159
rect 2820 17143 4275 17157
rect 2820 17133 2881 17143
rect 119 17115 2881 17133
rect 119 17051 135 17115
rect 199 17051 217 17115
rect 281 17051 299 17115
rect 363 17051 381 17115
rect 445 17051 463 17115
rect 527 17051 545 17115
rect 609 17051 627 17115
rect 691 17051 709 17115
rect 773 17051 791 17115
rect 855 17051 873 17115
rect 937 17051 955 17115
rect 1019 17051 1037 17115
rect 1101 17051 1119 17115
rect 1183 17051 1201 17115
rect 1265 17051 1283 17115
rect 1347 17051 1365 17115
rect 1429 17051 1447 17115
rect 1511 17051 1529 17115
rect 1593 17051 1611 17115
rect 1675 17051 1693 17115
rect 1757 17051 1775 17115
rect 1839 17051 1857 17115
rect 1921 17051 1939 17115
rect 2003 17051 2021 17115
rect 2085 17051 2103 17115
rect 2167 17051 2185 17115
rect 2249 17051 2267 17115
rect 2331 17051 2349 17115
rect 2413 17051 2431 17115
rect 2495 17051 2513 17115
rect 2577 17051 2594 17115
rect 2658 17051 2675 17115
rect 2739 17051 2756 17115
rect 2820 17079 2881 17115
rect 2945 17079 2963 17143
rect 3027 17079 3045 17143
rect 3109 17079 3127 17143
rect 3191 17079 3209 17143
rect 3273 17079 3291 17143
rect 3355 17079 3373 17143
rect 3437 17079 3455 17143
rect 3519 17079 3537 17143
rect 3601 17079 3619 17143
rect 3683 17079 3701 17143
rect 3765 17123 4275 17143
tri 4275 17123 4309 17157 sw
tri 10742 17123 10776 17157 se
rect 10776 17143 12231 17157
rect 10776 17123 11286 17143
rect 3765 17117 4309 17123
rect 3765 17079 3838 17117
rect 2820 17063 3838 17079
rect 2820 17051 2881 17063
rect 119 17033 2881 17051
rect 119 16969 135 17033
rect 199 16969 217 17033
rect 281 16969 299 17033
rect 363 16969 381 17033
rect 445 16969 463 17033
rect 527 16969 545 17033
rect 609 16969 627 17033
rect 691 16969 709 17033
rect 773 16969 791 17033
rect 855 16969 873 17033
rect 937 16969 955 17033
rect 1019 16969 1037 17033
rect 1101 16969 1119 17033
rect 1183 16969 1201 17033
rect 1265 16969 1283 17033
rect 1347 16969 1365 17033
rect 1429 16969 1447 17033
rect 1511 16969 1529 17033
rect 1593 16969 1611 17033
rect 1675 16969 1693 17033
rect 1757 16969 1775 17033
rect 1839 16969 1857 17033
rect 1921 16969 1939 17033
rect 2003 16969 2021 17033
rect 2085 16969 2103 17033
rect 2167 16969 2185 17033
rect 2249 16969 2267 17033
rect 2331 16969 2349 17033
rect 2413 16969 2431 17033
rect 2495 16969 2513 17033
rect 2577 16969 2594 17033
rect 2658 16969 2675 17033
rect 2739 16969 2756 17033
rect 2820 16999 2881 17033
rect 2945 16999 2963 17063
rect 3027 16999 3045 17063
rect 3109 16999 3127 17063
rect 3191 16999 3209 17063
rect 3273 16999 3291 17063
rect 3355 16999 3373 17063
rect 3437 16999 3455 17063
rect 3519 16999 3537 17063
rect 3601 16999 3619 17063
rect 3683 16999 3701 17063
rect 3765 17053 3838 17063
rect 3902 17053 3934 17117
rect 3998 17053 4030 17117
rect 4094 17053 4126 17117
rect 4190 17053 4222 17117
rect 4286 17053 4309 17117
rect 3765 17024 4309 17053
rect 3765 16999 3838 17024
rect 2820 16983 3838 16999
rect 2820 16969 2881 16983
rect 119 16951 2881 16969
rect 119 16887 135 16951
rect 199 16887 217 16951
rect 281 16887 299 16951
rect 363 16887 381 16951
rect 445 16887 463 16951
rect 527 16887 545 16951
rect 609 16887 627 16951
rect 691 16887 709 16951
rect 773 16887 791 16951
rect 855 16887 873 16951
rect 937 16887 955 16951
rect 1019 16887 1037 16951
rect 1101 16887 1119 16951
rect 1183 16887 1201 16951
rect 1265 16887 1283 16951
rect 1347 16887 1365 16951
rect 1429 16887 1447 16951
rect 1511 16887 1529 16951
rect 1593 16887 1611 16951
rect 1675 16887 1693 16951
rect 1757 16887 1775 16951
rect 1839 16887 1857 16951
rect 1921 16887 1939 16951
rect 2003 16887 2021 16951
rect 2085 16887 2103 16951
rect 2167 16887 2185 16951
rect 2249 16887 2267 16951
rect 2331 16887 2349 16951
rect 2413 16887 2431 16951
rect 2495 16887 2513 16951
rect 2577 16887 2594 16951
rect 2658 16887 2675 16951
rect 2739 16887 2756 16951
rect 2820 16919 2881 16951
rect 2945 16919 2963 16983
rect 3027 16919 3045 16983
rect 3109 16919 3127 16983
rect 3191 16919 3209 16983
rect 3273 16919 3291 16983
rect 3355 16919 3373 16983
rect 3437 16919 3455 16983
rect 3519 16919 3537 16983
rect 3601 16919 3619 16983
rect 3683 16919 3701 16983
rect 3765 16960 3838 16983
rect 3902 16960 3934 17024
rect 3998 16960 4030 17024
rect 4094 16960 4126 17024
rect 4190 16960 4222 17024
rect 4286 16960 4309 17024
rect 3765 16931 4309 16960
rect 3765 16919 3838 16931
rect 2820 16903 3838 16919
rect 2820 16887 2881 16903
rect 119 16869 2881 16887
rect 119 16805 135 16869
rect 199 16805 217 16869
rect 281 16805 299 16869
rect 363 16805 381 16869
rect 445 16805 463 16869
rect 527 16805 545 16869
rect 609 16805 627 16869
rect 691 16805 709 16869
rect 773 16805 791 16869
rect 855 16805 873 16869
rect 937 16805 955 16869
rect 1019 16805 1037 16869
rect 1101 16805 1119 16869
rect 1183 16805 1201 16869
rect 1265 16805 1283 16869
rect 1347 16805 1365 16869
rect 1429 16805 1447 16869
rect 1511 16805 1529 16869
rect 1593 16805 1611 16869
rect 1675 16805 1693 16869
rect 1757 16805 1775 16869
rect 1839 16805 1857 16869
rect 1921 16805 1939 16869
rect 2003 16805 2021 16869
rect 2085 16805 2103 16869
rect 2167 16805 2185 16869
rect 2249 16805 2267 16869
rect 2331 16805 2349 16869
rect 2413 16805 2431 16869
rect 2495 16805 2513 16869
rect 2577 16805 2594 16869
rect 2658 16805 2675 16869
rect 2739 16805 2756 16869
rect 2820 16839 2881 16869
rect 2945 16839 2963 16903
rect 3027 16839 3045 16903
rect 3109 16839 3127 16903
rect 3191 16839 3209 16903
rect 3273 16839 3291 16903
rect 3355 16839 3373 16903
rect 3437 16839 3455 16903
rect 3519 16839 3537 16903
rect 3601 16839 3619 16903
rect 3683 16839 3701 16903
rect 3765 16867 3838 16903
rect 3902 16867 3934 16931
rect 3998 16867 4030 16931
rect 4094 16867 4126 16931
rect 4190 16867 4222 16931
rect 4286 16867 4309 16931
rect 3765 16862 4309 16867
tri 4309 16862 4570 17123 sw
tri 10481 16862 10742 17123 se
rect 10742 17117 11286 17123
rect 10742 17053 10765 17117
rect 10829 17053 10861 17117
rect 10925 17053 10957 17117
rect 11021 17053 11053 17117
rect 11117 17053 11149 17117
rect 11213 17079 11286 17117
rect 11350 17079 11368 17143
rect 11432 17079 11450 17143
rect 11514 17079 11532 17143
rect 11596 17079 11614 17143
rect 11678 17079 11696 17143
rect 11760 17079 11778 17143
rect 11842 17079 11860 17143
rect 11924 17079 11942 17143
rect 12006 17079 12024 17143
rect 12088 17079 12106 17143
rect 12170 17133 12231 17143
rect 12295 17133 12312 17197
rect 12376 17133 12393 17197
rect 12457 17133 12474 17197
rect 12538 17133 12556 17197
rect 12620 17133 12638 17197
rect 12702 17133 12720 17197
rect 12784 17133 12802 17197
rect 12866 17133 12884 17197
rect 12948 17133 12966 17197
rect 13030 17133 13048 17197
rect 13112 17133 13130 17197
rect 13194 17133 13212 17197
rect 13276 17133 13294 17197
rect 13358 17133 13376 17197
rect 13440 17133 13458 17197
rect 13522 17133 13540 17197
rect 13604 17133 13622 17197
rect 13686 17133 13704 17197
rect 13768 17133 13786 17197
rect 13850 17133 13868 17197
rect 13932 17133 13950 17197
rect 14014 17133 14032 17197
rect 14096 17133 14114 17197
rect 14178 17133 14196 17197
rect 14260 17133 14278 17197
rect 14342 17133 14360 17197
rect 14424 17133 14442 17197
rect 14506 17133 14524 17197
rect 14588 17133 14606 17197
rect 14670 17133 14688 17197
rect 14752 17133 14770 17197
rect 14834 17133 14852 17197
rect 14916 17133 14932 17197
rect 12170 17115 14932 17133
rect 12170 17079 12231 17115
rect 11213 17063 12231 17079
rect 11213 17053 11286 17063
rect 10742 17024 11286 17053
rect 10742 16960 10765 17024
rect 10829 16960 10861 17024
rect 10925 16960 10957 17024
rect 11021 16960 11053 17024
rect 11117 16960 11149 17024
rect 11213 16999 11286 17024
rect 11350 16999 11368 17063
rect 11432 16999 11450 17063
rect 11514 16999 11532 17063
rect 11596 16999 11614 17063
rect 11678 16999 11696 17063
rect 11760 16999 11778 17063
rect 11842 16999 11860 17063
rect 11924 16999 11942 17063
rect 12006 16999 12024 17063
rect 12088 16999 12106 17063
rect 12170 17051 12231 17063
rect 12295 17051 12312 17115
rect 12376 17051 12393 17115
rect 12457 17051 12474 17115
rect 12538 17051 12556 17115
rect 12620 17051 12638 17115
rect 12702 17051 12720 17115
rect 12784 17051 12802 17115
rect 12866 17051 12884 17115
rect 12948 17051 12966 17115
rect 13030 17051 13048 17115
rect 13112 17051 13130 17115
rect 13194 17051 13212 17115
rect 13276 17051 13294 17115
rect 13358 17051 13376 17115
rect 13440 17051 13458 17115
rect 13522 17051 13540 17115
rect 13604 17051 13622 17115
rect 13686 17051 13704 17115
rect 13768 17051 13786 17115
rect 13850 17051 13868 17115
rect 13932 17051 13950 17115
rect 14014 17051 14032 17115
rect 14096 17051 14114 17115
rect 14178 17051 14196 17115
rect 14260 17051 14278 17115
rect 14342 17051 14360 17115
rect 14424 17051 14442 17115
rect 14506 17051 14524 17115
rect 14588 17051 14606 17115
rect 14670 17051 14688 17115
rect 14752 17051 14770 17115
rect 14834 17051 14852 17115
rect 14916 17051 14932 17115
rect 12170 17033 14932 17051
rect 12170 16999 12231 17033
rect 11213 16983 12231 16999
rect 11213 16960 11286 16983
rect 10742 16931 11286 16960
rect 10742 16867 10765 16931
rect 10829 16867 10861 16931
rect 10925 16867 10957 16931
rect 11021 16867 11053 16931
rect 11117 16867 11149 16931
rect 11213 16919 11286 16931
rect 11350 16919 11368 16983
rect 11432 16919 11450 16983
rect 11514 16919 11532 16983
rect 11596 16919 11614 16983
rect 11678 16919 11696 16983
rect 11760 16919 11778 16983
rect 11842 16919 11860 16983
rect 11924 16919 11942 16983
rect 12006 16919 12024 16983
rect 12088 16919 12106 16983
rect 12170 16969 12231 16983
rect 12295 16969 12312 17033
rect 12376 16969 12393 17033
rect 12457 16969 12474 17033
rect 12538 16969 12556 17033
rect 12620 16969 12638 17033
rect 12702 16969 12720 17033
rect 12784 16969 12802 17033
rect 12866 16969 12884 17033
rect 12948 16969 12966 17033
rect 13030 16969 13048 17033
rect 13112 16969 13130 17033
rect 13194 16969 13212 17033
rect 13276 16969 13294 17033
rect 13358 16969 13376 17033
rect 13440 16969 13458 17033
rect 13522 16969 13540 17033
rect 13604 16969 13622 17033
rect 13686 16969 13704 17033
rect 13768 16969 13786 17033
rect 13850 16969 13868 17033
rect 13932 16969 13950 17033
rect 14014 16969 14032 17033
rect 14096 16969 14114 17033
rect 14178 16969 14196 17033
rect 14260 16969 14278 17033
rect 14342 16969 14360 17033
rect 14424 16969 14442 17033
rect 14506 16969 14524 17033
rect 14588 16969 14606 17033
rect 14670 16969 14688 17033
rect 14752 16969 14770 17033
rect 14834 16969 14852 17033
rect 14916 16969 14932 17033
rect 12170 16951 14932 16969
rect 12170 16919 12231 16951
rect 11213 16903 12231 16919
rect 11213 16867 11286 16903
rect 10742 16862 11286 16867
rect 3765 16856 4570 16862
rect 3765 16839 4331 16856
rect 2820 16838 4331 16839
rect 2820 16823 3838 16838
rect 2820 16805 2881 16823
rect 119 16787 2881 16805
rect 119 16723 135 16787
rect 199 16723 217 16787
rect 281 16723 299 16787
rect 363 16723 381 16787
rect 445 16723 463 16787
rect 527 16723 545 16787
rect 609 16723 627 16787
rect 691 16723 709 16787
rect 773 16723 791 16787
rect 855 16723 873 16787
rect 937 16723 955 16787
rect 1019 16723 1037 16787
rect 1101 16723 1119 16787
rect 1183 16723 1201 16787
rect 1265 16723 1283 16787
rect 1347 16723 1365 16787
rect 1429 16723 1447 16787
rect 1511 16723 1529 16787
rect 1593 16723 1611 16787
rect 1675 16723 1693 16787
rect 1757 16723 1775 16787
rect 1839 16723 1857 16787
rect 1921 16723 1939 16787
rect 2003 16723 2021 16787
rect 2085 16723 2103 16787
rect 2167 16723 2185 16787
rect 2249 16723 2267 16787
rect 2331 16723 2349 16787
rect 2413 16723 2431 16787
rect 2495 16723 2513 16787
rect 2577 16723 2594 16787
rect 2658 16723 2675 16787
rect 2739 16723 2756 16787
rect 2820 16759 2881 16787
rect 2945 16759 2963 16823
rect 3027 16759 3045 16823
rect 3109 16759 3127 16823
rect 3191 16759 3209 16823
rect 3273 16759 3291 16823
rect 3355 16759 3373 16823
rect 3437 16759 3455 16823
rect 3519 16759 3537 16823
rect 3601 16759 3619 16823
rect 3683 16759 3701 16823
rect 3765 16774 3838 16823
rect 3902 16774 3934 16838
rect 3998 16774 4030 16838
rect 4094 16774 4126 16838
rect 4190 16774 4222 16838
rect 4286 16792 4331 16838
rect 4395 16792 4489 16856
rect 4553 16792 4570 16856
rect 4286 16774 4570 16792
rect 3765 16759 4570 16774
rect 2820 16746 4570 16759
rect 2820 16743 3838 16746
rect 2820 16723 2881 16743
rect 119 16705 2881 16723
rect 119 16641 135 16705
rect 199 16641 217 16705
rect 281 16641 299 16705
rect 363 16641 381 16705
rect 445 16641 463 16705
rect 527 16641 545 16705
rect 609 16641 627 16705
rect 691 16641 709 16705
rect 773 16641 791 16705
rect 855 16641 873 16705
rect 937 16641 955 16705
rect 1019 16641 1037 16705
rect 1101 16641 1119 16705
rect 1183 16641 1201 16705
rect 1265 16641 1283 16705
rect 1347 16641 1365 16705
rect 1429 16641 1447 16705
rect 1511 16641 1529 16705
rect 1593 16641 1611 16705
rect 1675 16641 1693 16705
rect 1757 16641 1775 16705
rect 1839 16641 1857 16705
rect 1921 16641 1939 16705
rect 2003 16641 2021 16705
rect 2085 16641 2103 16705
rect 2167 16641 2185 16705
rect 2249 16641 2267 16705
rect 2331 16641 2349 16705
rect 2413 16641 2431 16705
rect 2495 16641 2513 16705
rect 2577 16641 2594 16705
rect 2658 16641 2675 16705
rect 2739 16641 2756 16705
rect 2820 16679 2881 16705
rect 2945 16679 2963 16743
rect 3027 16679 3045 16743
rect 3109 16679 3127 16743
rect 3191 16679 3209 16743
rect 3273 16679 3291 16743
rect 3355 16679 3373 16743
rect 3437 16679 3455 16743
rect 3519 16679 3537 16743
rect 3601 16679 3619 16743
rect 3683 16679 3701 16743
rect 3765 16682 3838 16743
rect 3902 16682 3934 16746
rect 3998 16682 4030 16746
rect 4094 16682 4126 16746
rect 4190 16682 4222 16746
rect 4286 16682 4331 16746
rect 4395 16682 4489 16746
rect 4553 16682 4570 16746
rect 3765 16679 4570 16682
rect 2820 16663 4570 16679
rect 2820 16641 2881 16663
rect 119 16623 2881 16641
rect 119 16559 135 16623
rect 199 16559 217 16623
rect 281 16559 299 16623
rect 363 16559 381 16623
rect 445 16559 463 16623
rect 527 16559 545 16623
rect 609 16559 627 16623
rect 691 16559 709 16623
rect 773 16559 791 16623
rect 855 16559 873 16623
rect 937 16559 955 16623
rect 1019 16559 1037 16623
rect 1101 16559 1119 16623
rect 1183 16559 1201 16623
rect 1265 16559 1283 16623
rect 1347 16559 1365 16623
rect 1429 16559 1447 16623
rect 1511 16559 1529 16623
rect 1593 16559 1611 16623
rect 1675 16559 1693 16623
rect 1757 16559 1775 16623
rect 1839 16559 1857 16623
rect 1921 16559 1939 16623
rect 2003 16559 2021 16623
rect 2085 16559 2103 16623
rect 2167 16559 2185 16623
rect 2249 16559 2267 16623
rect 2331 16559 2349 16623
rect 2413 16559 2431 16623
rect 2495 16559 2513 16623
rect 2577 16559 2594 16623
rect 2658 16559 2675 16623
rect 2739 16559 2756 16623
rect 2820 16599 2881 16623
rect 2945 16599 2963 16663
rect 3027 16599 3045 16663
rect 3109 16599 3127 16663
rect 3191 16599 3209 16663
rect 3273 16599 3291 16663
rect 3355 16599 3373 16663
rect 3437 16599 3455 16663
rect 3519 16599 3537 16663
rect 3601 16599 3619 16663
rect 3683 16599 3701 16663
rect 3765 16654 4570 16663
rect 3765 16599 3838 16654
rect 2820 16590 3838 16599
rect 3902 16590 3934 16654
rect 3998 16590 4030 16654
rect 4094 16590 4126 16654
rect 4190 16590 4222 16654
rect 4286 16636 4570 16654
rect 4286 16590 4331 16636
rect 2820 16572 4331 16590
rect 4395 16572 4489 16636
rect 4553 16572 4570 16636
rect 2820 16566 4570 16572
tri 4570 16566 4866 16862 sw
tri 10185 16566 10481 16862 se
rect 10481 16856 11286 16862
rect 10481 16792 10498 16856
rect 10562 16792 10656 16856
rect 10720 16839 11286 16856
rect 11350 16839 11368 16903
rect 11432 16839 11450 16903
rect 11514 16839 11532 16903
rect 11596 16839 11614 16903
rect 11678 16839 11696 16903
rect 11760 16839 11778 16903
rect 11842 16839 11860 16903
rect 11924 16839 11942 16903
rect 12006 16839 12024 16903
rect 12088 16839 12106 16903
rect 12170 16887 12231 16903
rect 12295 16887 12312 16951
rect 12376 16887 12393 16951
rect 12457 16887 12474 16951
rect 12538 16887 12556 16951
rect 12620 16887 12638 16951
rect 12702 16887 12720 16951
rect 12784 16887 12802 16951
rect 12866 16887 12884 16951
rect 12948 16887 12966 16951
rect 13030 16887 13048 16951
rect 13112 16887 13130 16951
rect 13194 16887 13212 16951
rect 13276 16887 13294 16951
rect 13358 16887 13376 16951
rect 13440 16887 13458 16951
rect 13522 16887 13540 16951
rect 13604 16887 13622 16951
rect 13686 16887 13704 16951
rect 13768 16887 13786 16951
rect 13850 16887 13868 16951
rect 13932 16887 13950 16951
rect 14014 16887 14032 16951
rect 14096 16887 14114 16951
rect 14178 16887 14196 16951
rect 14260 16887 14278 16951
rect 14342 16887 14360 16951
rect 14424 16887 14442 16951
rect 14506 16887 14524 16951
rect 14588 16887 14606 16951
rect 14670 16887 14688 16951
rect 14752 16887 14770 16951
rect 14834 16887 14852 16951
rect 14916 16887 14932 16951
rect 12170 16869 14932 16887
rect 12170 16839 12231 16869
rect 10720 16838 12231 16839
rect 10720 16792 10765 16838
rect 10481 16774 10765 16792
rect 10829 16774 10861 16838
rect 10925 16774 10957 16838
rect 11021 16774 11053 16838
rect 11117 16774 11149 16838
rect 11213 16823 12231 16838
rect 11213 16774 11286 16823
rect 10481 16759 11286 16774
rect 11350 16759 11368 16823
rect 11432 16759 11450 16823
rect 11514 16759 11532 16823
rect 11596 16759 11614 16823
rect 11678 16759 11696 16823
rect 11760 16759 11778 16823
rect 11842 16759 11860 16823
rect 11924 16759 11942 16823
rect 12006 16759 12024 16823
rect 12088 16759 12106 16823
rect 12170 16805 12231 16823
rect 12295 16805 12312 16869
rect 12376 16805 12393 16869
rect 12457 16805 12474 16869
rect 12538 16805 12556 16869
rect 12620 16805 12638 16869
rect 12702 16805 12720 16869
rect 12784 16805 12802 16869
rect 12866 16805 12884 16869
rect 12948 16805 12966 16869
rect 13030 16805 13048 16869
rect 13112 16805 13130 16869
rect 13194 16805 13212 16869
rect 13276 16805 13294 16869
rect 13358 16805 13376 16869
rect 13440 16805 13458 16869
rect 13522 16805 13540 16869
rect 13604 16805 13622 16869
rect 13686 16805 13704 16869
rect 13768 16805 13786 16869
rect 13850 16805 13868 16869
rect 13932 16805 13950 16869
rect 14014 16805 14032 16869
rect 14096 16805 14114 16869
rect 14178 16805 14196 16869
rect 14260 16805 14278 16869
rect 14342 16805 14360 16869
rect 14424 16805 14442 16869
rect 14506 16805 14524 16869
rect 14588 16805 14606 16869
rect 14670 16805 14688 16869
rect 14752 16805 14770 16869
rect 14834 16805 14852 16869
rect 14916 16805 14932 16869
rect 12170 16787 14932 16805
rect 12170 16759 12231 16787
rect 10481 16746 12231 16759
rect 10481 16682 10498 16746
rect 10562 16682 10656 16746
rect 10720 16682 10765 16746
rect 10829 16682 10861 16746
rect 10925 16682 10957 16746
rect 11021 16682 11053 16746
rect 11117 16682 11149 16746
rect 11213 16743 12231 16746
rect 11213 16682 11286 16743
rect 10481 16679 11286 16682
rect 11350 16679 11368 16743
rect 11432 16679 11450 16743
rect 11514 16679 11532 16743
rect 11596 16679 11614 16743
rect 11678 16679 11696 16743
rect 11760 16679 11778 16743
rect 11842 16679 11860 16743
rect 11924 16679 11942 16743
rect 12006 16679 12024 16743
rect 12088 16679 12106 16743
rect 12170 16723 12231 16743
rect 12295 16723 12312 16787
rect 12376 16723 12393 16787
rect 12457 16723 12474 16787
rect 12538 16723 12556 16787
rect 12620 16723 12638 16787
rect 12702 16723 12720 16787
rect 12784 16723 12802 16787
rect 12866 16723 12884 16787
rect 12948 16723 12966 16787
rect 13030 16723 13048 16787
rect 13112 16723 13130 16787
rect 13194 16723 13212 16787
rect 13276 16723 13294 16787
rect 13358 16723 13376 16787
rect 13440 16723 13458 16787
rect 13522 16723 13540 16787
rect 13604 16723 13622 16787
rect 13686 16723 13704 16787
rect 13768 16723 13786 16787
rect 13850 16723 13868 16787
rect 13932 16723 13950 16787
rect 14014 16723 14032 16787
rect 14096 16723 14114 16787
rect 14178 16723 14196 16787
rect 14260 16723 14278 16787
rect 14342 16723 14360 16787
rect 14424 16723 14442 16787
rect 14506 16723 14524 16787
rect 14588 16723 14606 16787
rect 14670 16723 14688 16787
rect 14752 16723 14770 16787
rect 14834 16723 14852 16787
rect 14916 16723 14932 16787
rect 12170 16705 14932 16723
rect 12170 16679 12231 16705
rect 10481 16663 12231 16679
rect 10481 16654 11286 16663
rect 10481 16636 10765 16654
rect 10481 16572 10498 16636
rect 10562 16572 10656 16636
rect 10720 16590 10765 16636
rect 10829 16590 10861 16654
rect 10925 16590 10957 16654
rect 11021 16590 11053 16654
rect 11117 16590 11149 16654
rect 11213 16599 11286 16654
rect 11350 16599 11368 16663
rect 11432 16599 11450 16663
rect 11514 16599 11532 16663
rect 11596 16599 11614 16663
rect 11678 16599 11696 16663
rect 11760 16599 11778 16663
rect 11842 16599 11860 16663
rect 11924 16599 11942 16663
rect 12006 16599 12024 16663
rect 12088 16599 12106 16663
rect 12170 16641 12231 16663
rect 12295 16641 12312 16705
rect 12376 16641 12393 16705
rect 12457 16641 12474 16705
rect 12538 16641 12556 16705
rect 12620 16641 12638 16705
rect 12702 16641 12720 16705
rect 12784 16641 12802 16705
rect 12866 16641 12884 16705
rect 12948 16641 12966 16705
rect 13030 16641 13048 16705
rect 13112 16641 13130 16705
rect 13194 16641 13212 16705
rect 13276 16641 13294 16705
rect 13358 16641 13376 16705
rect 13440 16641 13458 16705
rect 13522 16641 13540 16705
rect 13604 16641 13622 16705
rect 13686 16641 13704 16705
rect 13768 16641 13786 16705
rect 13850 16641 13868 16705
rect 13932 16641 13950 16705
rect 14014 16641 14032 16705
rect 14096 16641 14114 16705
rect 14178 16641 14196 16705
rect 14260 16641 14278 16705
rect 14342 16641 14360 16705
rect 14424 16641 14442 16705
rect 14506 16641 14524 16705
rect 14588 16641 14606 16705
rect 14670 16641 14688 16705
rect 14752 16641 14770 16705
rect 14834 16641 14852 16705
rect 14916 16641 14932 16705
rect 12170 16623 14932 16641
rect 12170 16599 12231 16623
rect 11213 16590 12231 16599
rect 10720 16572 12231 16590
rect 10481 16566 12231 16572
rect 2820 16559 4866 16566
tri 4866 16559 4873 16566 sw
tri 10178 16559 10185 16566 se
rect 10185 16559 12231 16566
rect 12295 16559 12312 16623
rect 12376 16559 12393 16623
rect 12457 16559 12474 16623
rect 12538 16559 12556 16623
rect 12620 16559 12638 16623
rect 12702 16559 12720 16623
rect 12784 16559 12802 16623
rect 12866 16559 12884 16623
rect 12948 16559 12966 16623
rect 13030 16559 13048 16623
rect 13112 16559 13130 16623
rect 13194 16559 13212 16623
rect 13276 16559 13294 16623
rect 13358 16559 13376 16623
rect 13440 16559 13458 16623
rect 13522 16559 13540 16623
rect 13604 16559 13622 16623
rect 13686 16559 13704 16623
rect 13768 16559 13786 16623
rect 13850 16559 13868 16623
rect 13932 16559 13950 16623
rect 14014 16559 14032 16623
rect 14096 16559 14114 16623
rect 14178 16559 14196 16623
rect 14260 16559 14278 16623
rect 14342 16559 14360 16623
rect 14424 16559 14442 16623
rect 14506 16559 14524 16623
rect 14588 16559 14606 16623
rect 14670 16559 14688 16623
rect 14752 16559 14770 16623
rect 14834 16559 14852 16623
rect 14916 16559 14932 16623
rect 119 16533 4873 16559
tri 4873 16533 4899 16559 sw
tri 10177 16558 10178 16559 se
rect 10178 16558 14932 16559
rect 119 16524 4899 16533
rect 119 16460 157 16524
rect 221 16460 237 16524
rect 301 16460 317 16524
rect 381 16460 397 16524
rect 461 16460 477 16524
rect 541 16460 557 16524
rect 621 16460 637 16524
rect 701 16460 717 16524
rect 781 16460 797 16524
rect 861 16460 877 16524
rect 941 16460 957 16524
rect 1021 16460 1037 16524
rect 1101 16460 1117 16524
rect 1181 16460 1197 16524
rect 1261 16460 1277 16524
rect 1341 16460 1357 16524
rect 1421 16460 1437 16524
rect 1501 16460 1517 16524
rect 1581 16460 1597 16524
rect 1661 16460 1677 16524
rect 1741 16460 1757 16524
rect 1821 16460 1837 16524
rect 1901 16460 1917 16524
rect 1981 16460 1997 16524
rect 2061 16460 2077 16524
rect 2141 16460 2157 16524
rect 2221 16460 2237 16524
rect 2301 16460 2317 16524
rect 2381 16460 2397 16524
rect 2461 16460 2477 16524
rect 2541 16460 2557 16524
rect 2621 16460 2637 16524
rect 2701 16460 2717 16524
rect 2781 16460 2797 16524
rect 2861 16460 2877 16524
rect 2941 16460 2957 16524
rect 3021 16460 3037 16524
rect 3101 16460 3117 16524
rect 3181 16460 3197 16524
rect 3261 16460 3277 16524
rect 3341 16460 3357 16524
rect 3421 16460 3437 16524
rect 3501 16460 3517 16524
rect 3581 16460 3597 16524
rect 3661 16460 3677 16524
rect 3741 16460 3757 16524
rect 3821 16460 3837 16524
rect 3901 16460 3917 16524
rect 3981 16460 3997 16524
rect 4061 16460 4077 16524
rect 4141 16460 4157 16524
rect 4221 16460 4237 16524
rect 4301 16460 4317 16524
rect 4381 16460 4397 16524
rect 4461 16460 4477 16524
rect 4541 16460 4557 16524
rect 4621 16460 4637 16524
rect 4701 16460 4717 16524
rect 4781 16460 4797 16524
rect 4861 16460 4899 16524
rect 119 16443 4899 16460
rect 119 16379 157 16443
rect 221 16379 237 16443
rect 301 16379 317 16443
rect 381 16379 397 16443
rect 461 16379 477 16443
rect 541 16379 557 16443
rect 621 16379 637 16443
rect 701 16379 717 16443
rect 781 16379 797 16443
rect 861 16379 877 16443
rect 941 16379 957 16443
rect 1021 16379 1037 16443
rect 1101 16379 1117 16443
rect 1181 16379 1197 16443
rect 1261 16379 1277 16443
rect 1341 16379 1357 16443
rect 1421 16379 1437 16443
rect 1501 16379 1517 16443
rect 1581 16379 1597 16443
rect 1661 16379 1677 16443
rect 1741 16379 1757 16443
rect 1821 16379 1837 16443
rect 1901 16379 1917 16443
rect 1981 16379 1997 16443
rect 2061 16379 2077 16443
rect 2141 16379 2157 16443
rect 2221 16379 2237 16443
rect 2301 16379 2317 16443
rect 2381 16379 2397 16443
rect 2461 16379 2477 16443
rect 2541 16379 2557 16443
rect 2621 16379 2637 16443
rect 2701 16379 2717 16443
rect 2781 16379 2797 16443
rect 2861 16379 2877 16443
rect 2941 16379 2957 16443
rect 3021 16379 3037 16443
rect 3101 16379 3117 16443
rect 3181 16379 3197 16443
rect 3261 16379 3277 16443
rect 3341 16379 3357 16443
rect 3421 16379 3437 16443
rect 3501 16379 3517 16443
rect 3581 16379 3597 16443
rect 3661 16379 3677 16443
rect 3741 16379 3757 16443
rect 3821 16379 3837 16443
rect 3901 16379 3917 16443
rect 3981 16379 3997 16443
rect 4061 16379 4077 16443
rect 4141 16379 4157 16443
rect 4221 16379 4237 16443
rect 4301 16379 4317 16443
rect 4381 16379 4397 16443
rect 4461 16379 4477 16443
rect 4541 16379 4557 16443
rect 4621 16379 4637 16443
rect 4701 16379 4717 16443
rect 4781 16379 4797 16443
rect 4861 16379 4899 16443
rect 119 16362 4899 16379
rect 119 16298 157 16362
rect 221 16298 237 16362
rect 301 16298 317 16362
rect 381 16298 397 16362
rect 461 16298 477 16362
rect 541 16298 557 16362
rect 621 16298 637 16362
rect 701 16298 717 16362
rect 781 16298 797 16362
rect 861 16298 877 16362
rect 941 16298 957 16362
rect 1021 16298 1037 16362
rect 1101 16298 1117 16362
rect 1181 16298 1197 16362
rect 1261 16298 1277 16362
rect 1341 16298 1357 16362
rect 1421 16298 1437 16362
rect 1501 16298 1517 16362
rect 1581 16298 1597 16362
rect 1661 16298 1677 16362
rect 1741 16298 1757 16362
rect 1821 16298 1837 16362
rect 1901 16298 1917 16362
rect 1981 16298 1997 16362
rect 2061 16298 2077 16362
rect 2141 16298 2157 16362
rect 2221 16298 2237 16362
rect 2301 16298 2317 16362
rect 2381 16298 2397 16362
rect 2461 16298 2477 16362
rect 2541 16298 2557 16362
rect 2621 16298 2637 16362
rect 2701 16298 2717 16362
rect 2781 16298 2797 16362
rect 2861 16298 2877 16362
rect 2941 16298 2957 16362
rect 3021 16298 3037 16362
rect 3101 16298 3117 16362
rect 3181 16298 3197 16362
rect 3261 16298 3277 16362
rect 3341 16298 3357 16362
rect 3421 16298 3437 16362
rect 3501 16298 3517 16362
rect 3581 16298 3597 16362
rect 3661 16298 3677 16362
rect 3741 16298 3757 16362
rect 3821 16298 3837 16362
rect 3901 16298 3917 16362
rect 3981 16298 3997 16362
rect 4061 16298 4077 16362
rect 4141 16298 4157 16362
rect 4221 16298 4237 16362
rect 4301 16298 4317 16362
rect 4381 16298 4397 16362
rect 4461 16298 4477 16362
rect 4541 16298 4557 16362
rect 4621 16298 4637 16362
rect 4701 16298 4717 16362
rect 4781 16298 4797 16362
rect 4861 16298 4899 16362
rect 119 16281 4899 16298
rect 119 16217 157 16281
rect 221 16217 237 16281
rect 301 16217 317 16281
rect 381 16217 397 16281
rect 461 16217 477 16281
rect 541 16217 557 16281
rect 621 16217 637 16281
rect 701 16217 717 16281
rect 781 16217 797 16281
rect 861 16217 877 16281
rect 941 16217 957 16281
rect 1021 16217 1037 16281
rect 1101 16217 1117 16281
rect 1181 16217 1197 16281
rect 1261 16217 1277 16281
rect 1341 16217 1357 16281
rect 1421 16217 1437 16281
rect 1501 16217 1517 16281
rect 1581 16217 1597 16281
rect 1661 16217 1677 16281
rect 1741 16217 1757 16281
rect 1821 16217 1837 16281
rect 1901 16217 1917 16281
rect 1981 16217 1997 16281
rect 2061 16217 2077 16281
rect 2141 16217 2157 16281
rect 2221 16217 2237 16281
rect 2301 16217 2317 16281
rect 2381 16217 2397 16281
rect 2461 16217 2477 16281
rect 2541 16217 2557 16281
rect 2621 16217 2637 16281
rect 2701 16217 2717 16281
rect 2781 16217 2797 16281
rect 2861 16217 2877 16281
rect 2941 16217 2957 16281
rect 3021 16217 3037 16281
rect 3101 16217 3117 16281
rect 3181 16217 3197 16281
rect 3261 16217 3277 16281
rect 3341 16217 3357 16281
rect 3421 16217 3437 16281
rect 3501 16217 3517 16281
rect 3581 16217 3597 16281
rect 3661 16217 3677 16281
rect 3741 16217 3757 16281
rect 3821 16217 3837 16281
rect 3901 16217 3917 16281
rect 3981 16217 3997 16281
rect 4061 16217 4077 16281
rect 4141 16217 4157 16281
rect 4221 16217 4237 16281
rect 4301 16217 4317 16281
rect 4381 16217 4397 16281
rect 4461 16217 4477 16281
rect 4541 16217 4557 16281
rect 4621 16217 4637 16281
rect 4701 16217 4717 16281
rect 4781 16217 4797 16281
rect 4861 16217 4899 16281
rect 119 16200 4899 16217
rect 119 16136 157 16200
rect 221 16136 237 16200
rect 301 16136 317 16200
rect 381 16136 397 16200
rect 461 16136 477 16200
rect 541 16136 557 16200
rect 621 16136 637 16200
rect 701 16136 717 16200
rect 781 16136 797 16200
rect 861 16136 877 16200
rect 941 16136 957 16200
rect 1021 16136 1037 16200
rect 1101 16136 1117 16200
rect 1181 16136 1197 16200
rect 1261 16136 1277 16200
rect 1341 16136 1357 16200
rect 1421 16136 1437 16200
rect 1501 16136 1517 16200
rect 1581 16136 1597 16200
rect 1661 16136 1677 16200
rect 1741 16136 1757 16200
rect 1821 16136 1837 16200
rect 1901 16136 1917 16200
rect 1981 16136 1997 16200
rect 2061 16136 2077 16200
rect 2141 16136 2157 16200
rect 2221 16136 2237 16200
rect 2301 16136 2317 16200
rect 2381 16136 2397 16200
rect 2461 16136 2477 16200
rect 2541 16136 2557 16200
rect 2621 16136 2637 16200
rect 2701 16136 2717 16200
rect 2781 16136 2797 16200
rect 2861 16136 2877 16200
rect 2941 16136 2957 16200
rect 3021 16136 3037 16200
rect 3101 16136 3117 16200
rect 3181 16136 3197 16200
rect 3261 16136 3277 16200
rect 3341 16136 3357 16200
rect 3421 16136 3437 16200
rect 3501 16136 3517 16200
rect 3581 16136 3597 16200
rect 3661 16136 3677 16200
rect 3741 16136 3757 16200
rect 3821 16136 3837 16200
rect 3901 16136 3917 16200
rect 3981 16136 3997 16200
rect 4061 16136 4077 16200
rect 4141 16136 4157 16200
rect 4221 16136 4237 16200
rect 4301 16136 4317 16200
rect 4381 16136 4397 16200
rect 4461 16136 4477 16200
rect 4541 16136 4557 16200
rect 4621 16136 4637 16200
rect 4701 16136 4717 16200
rect 4781 16136 4797 16200
rect 4861 16136 4899 16200
rect 119 16119 4899 16136
rect 119 16055 157 16119
rect 221 16055 237 16119
rect 301 16055 317 16119
rect 381 16055 397 16119
rect 461 16055 477 16119
rect 541 16055 557 16119
rect 621 16055 637 16119
rect 701 16055 717 16119
rect 781 16055 797 16119
rect 861 16055 877 16119
rect 941 16055 957 16119
rect 1021 16055 1037 16119
rect 1101 16055 1117 16119
rect 1181 16055 1197 16119
rect 1261 16055 1277 16119
rect 1341 16055 1357 16119
rect 1421 16055 1437 16119
rect 1501 16055 1517 16119
rect 1581 16055 1597 16119
rect 1661 16055 1677 16119
rect 1741 16055 1757 16119
rect 1821 16055 1837 16119
rect 1901 16055 1917 16119
rect 1981 16055 1997 16119
rect 2061 16055 2077 16119
rect 2141 16055 2157 16119
rect 2221 16055 2237 16119
rect 2301 16055 2317 16119
rect 2381 16055 2397 16119
rect 2461 16055 2477 16119
rect 2541 16055 2557 16119
rect 2621 16055 2637 16119
rect 2701 16055 2717 16119
rect 2781 16055 2797 16119
rect 2861 16055 2877 16119
rect 2941 16055 2957 16119
rect 3021 16055 3037 16119
rect 3101 16055 3117 16119
rect 3181 16055 3197 16119
rect 3261 16055 3277 16119
rect 3341 16055 3357 16119
rect 3421 16055 3437 16119
rect 3501 16055 3517 16119
rect 3581 16055 3597 16119
rect 3661 16055 3677 16119
rect 3741 16055 3757 16119
rect 3821 16055 3837 16119
rect 3901 16055 3917 16119
rect 3981 16055 3997 16119
rect 4061 16055 4077 16119
rect 4141 16055 4157 16119
rect 4221 16055 4237 16119
rect 4301 16055 4317 16119
rect 4381 16055 4397 16119
rect 4461 16055 4477 16119
rect 4541 16055 4557 16119
rect 4621 16055 4637 16119
rect 4701 16055 4717 16119
rect 4781 16055 4797 16119
rect 4861 16055 4899 16119
rect 119 16038 4899 16055
rect 119 15974 157 16038
rect 221 15974 237 16038
rect 301 15974 317 16038
rect 381 15974 397 16038
rect 461 15974 477 16038
rect 541 15974 557 16038
rect 621 15974 637 16038
rect 701 15974 717 16038
rect 781 15974 797 16038
rect 861 15974 877 16038
rect 941 15974 957 16038
rect 1021 15974 1037 16038
rect 1101 15974 1117 16038
rect 1181 15974 1197 16038
rect 1261 15974 1277 16038
rect 1341 15974 1357 16038
rect 1421 15974 1437 16038
rect 1501 15974 1517 16038
rect 1581 15974 1597 16038
rect 1661 15974 1677 16038
rect 1741 15974 1757 16038
rect 1821 15974 1837 16038
rect 1901 15974 1917 16038
rect 1981 15974 1997 16038
rect 2061 15974 2077 16038
rect 2141 15974 2157 16038
rect 2221 15974 2237 16038
rect 2301 15974 2317 16038
rect 2381 15974 2397 16038
rect 2461 15974 2477 16038
rect 2541 15974 2557 16038
rect 2621 15974 2637 16038
rect 2701 15974 2717 16038
rect 2781 15974 2797 16038
rect 2861 15974 2877 16038
rect 2941 15974 2957 16038
rect 3021 15974 3037 16038
rect 3101 15974 3117 16038
rect 3181 15974 3197 16038
rect 3261 15974 3277 16038
rect 3341 15974 3357 16038
rect 3421 15974 3437 16038
rect 3501 15974 3517 16038
rect 3581 15974 3597 16038
rect 3661 15974 3677 16038
rect 3741 15974 3757 16038
rect 3821 15974 3837 16038
rect 3901 15974 3917 16038
rect 3981 15974 3997 16038
rect 4061 15974 4077 16038
rect 4141 15974 4157 16038
rect 4221 15974 4237 16038
rect 4301 15974 4317 16038
rect 4381 15974 4397 16038
rect 4461 15974 4477 16038
rect 4541 15974 4557 16038
rect 4621 15974 4637 16038
rect 4701 15974 4717 16038
rect 4781 15974 4797 16038
rect 4861 15974 4899 16038
rect 119 15957 4899 15974
rect 119 15893 157 15957
rect 221 15893 237 15957
rect 301 15893 317 15957
rect 381 15893 397 15957
rect 461 15893 477 15957
rect 541 15893 557 15957
rect 621 15893 637 15957
rect 701 15893 717 15957
rect 781 15893 797 15957
rect 861 15893 877 15957
rect 941 15893 957 15957
rect 1021 15893 1037 15957
rect 1101 15893 1117 15957
rect 1181 15893 1197 15957
rect 1261 15893 1277 15957
rect 1341 15893 1357 15957
rect 1421 15893 1437 15957
rect 1501 15893 1517 15957
rect 1581 15893 1597 15957
rect 1661 15893 1677 15957
rect 1741 15893 1757 15957
rect 1821 15893 1837 15957
rect 1901 15893 1917 15957
rect 1981 15893 1997 15957
rect 2061 15893 2077 15957
rect 2141 15893 2157 15957
rect 2221 15893 2237 15957
rect 2301 15893 2317 15957
rect 2381 15893 2397 15957
rect 2461 15893 2477 15957
rect 2541 15893 2557 15957
rect 2621 15893 2637 15957
rect 2701 15893 2717 15957
rect 2781 15893 2797 15957
rect 2861 15893 2877 15957
rect 2941 15893 2957 15957
rect 3021 15893 3037 15957
rect 3101 15893 3117 15957
rect 3181 15893 3197 15957
rect 3261 15893 3277 15957
rect 3341 15893 3357 15957
rect 3421 15893 3437 15957
rect 3501 15893 3517 15957
rect 3581 15893 3597 15957
rect 3661 15893 3677 15957
rect 3741 15893 3757 15957
rect 3821 15893 3837 15957
rect 3901 15893 3917 15957
rect 3981 15893 3997 15957
rect 4061 15893 4077 15957
rect 4141 15893 4157 15957
rect 4221 15893 4237 15957
rect 4301 15893 4317 15957
rect 4381 15893 4397 15957
rect 4461 15893 4477 15957
rect 4541 15893 4557 15957
rect 4621 15893 4637 15957
rect 4701 15893 4717 15957
rect 4781 15893 4797 15957
rect 4861 15893 4899 15957
rect 119 15876 4899 15893
rect 119 15812 157 15876
rect 221 15812 237 15876
rect 301 15812 317 15876
rect 381 15812 397 15876
rect 461 15812 477 15876
rect 541 15812 557 15876
rect 621 15812 637 15876
rect 701 15812 717 15876
rect 781 15812 797 15876
rect 861 15812 877 15876
rect 941 15812 957 15876
rect 1021 15812 1037 15876
rect 1101 15812 1117 15876
rect 1181 15812 1197 15876
rect 1261 15812 1277 15876
rect 1341 15812 1357 15876
rect 1421 15812 1437 15876
rect 1501 15812 1517 15876
rect 1581 15812 1597 15876
rect 1661 15812 1677 15876
rect 1741 15812 1757 15876
rect 1821 15812 1837 15876
rect 1901 15812 1917 15876
rect 1981 15812 1997 15876
rect 2061 15812 2077 15876
rect 2141 15812 2157 15876
rect 2221 15812 2237 15876
rect 2301 15812 2317 15876
rect 2381 15812 2397 15876
rect 2461 15812 2477 15876
rect 2541 15812 2557 15876
rect 2621 15812 2637 15876
rect 2701 15812 2717 15876
rect 2781 15812 2797 15876
rect 2861 15812 2877 15876
rect 2941 15812 2957 15876
rect 3021 15812 3037 15876
rect 3101 15812 3117 15876
rect 3181 15812 3197 15876
rect 3261 15812 3277 15876
rect 3341 15812 3357 15876
rect 3421 15812 3437 15876
rect 3501 15812 3517 15876
rect 3581 15812 3597 15876
rect 3661 15812 3677 15876
rect 3741 15812 3757 15876
rect 3821 15812 3837 15876
rect 3901 15812 3917 15876
rect 3981 15812 3997 15876
rect 4061 15812 4077 15876
rect 4141 15812 4157 15876
rect 4221 15812 4237 15876
rect 4301 15812 4317 15876
rect 4381 15812 4397 15876
rect 4461 15812 4477 15876
rect 4541 15812 4557 15876
rect 4621 15812 4637 15876
rect 4701 15812 4717 15876
rect 4781 15812 4797 15876
rect 4861 15812 4899 15876
rect 119 15795 4899 15812
rect 119 15731 157 15795
rect 221 15731 237 15795
rect 301 15731 317 15795
rect 381 15731 397 15795
rect 461 15731 477 15795
rect 541 15731 557 15795
rect 621 15731 637 15795
rect 701 15731 717 15795
rect 781 15731 797 15795
rect 861 15731 877 15795
rect 941 15731 957 15795
rect 1021 15731 1037 15795
rect 1101 15731 1117 15795
rect 1181 15731 1197 15795
rect 1261 15731 1277 15795
rect 1341 15731 1357 15795
rect 1421 15731 1437 15795
rect 1501 15731 1517 15795
rect 1581 15731 1597 15795
rect 1661 15731 1677 15795
rect 1741 15731 1757 15795
rect 1821 15731 1837 15795
rect 1901 15731 1917 15795
rect 1981 15731 1997 15795
rect 2061 15731 2077 15795
rect 2141 15731 2157 15795
rect 2221 15731 2237 15795
rect 2301 15731 2317 15795
rect 2381 15731 2397 15795
rect 2461 15731 2477 15795
rect 2541 15731 2557 15795
rect 2621 15731 2637 15795
rect 2701 15731 2717 15795
rect 2781 15731 2797 15795
rect 2861 15731 2877 15795
rect 2941 15731 2957 15795
rect 3021 15731 3037 15795
rect 3101 15731 3117 15795
rect 3181 15731 3197 15795
rect 3261 15731 3277 15795
rect 3341 15731 3357 15795
rect 3421 15731 3437 15795
rect 3501 15731 3517 15795
rect 3581 15731 3597 15795
rect 3661 15731 3677 15795
rect 3741 15731 3757 15795
rect 3821 15731 3837 15795
rect 3901 15731 3917 15795
rect 3981 15731 3997 15795
rect 4061 15731 4077 15795
rect 4141 15731 4157 15795
rect 4221 15731 4237 15795
rect 4301 15731 4317 15795
rect 4381 15731 4397 15795
rect 4461 15731 4477 15795
rect 4541 15731 4557 15795
rect 4621 15731 4637 15795
rect 4701 15731 4717 15795
rect 4781 15731 4797 15795
rect 4861 15731 4899 15795
rect 119 15714 4899 15731
rect 119 15650 157 15714
rect 221 15650 237 15714
rect 301 15650 317 15714
rect 381 15650 397 15714
rect 461 15650 477 15714
rect 541 15650 557 15714
rect 621 15650 637 15714
rect 701 15650 717 15714
rect 781 15650 797 15714
rect 861 15650 877 15714
rect 941 15650 957 15714
rect 1021 15650 1037 15714
rect 1101 15650 1117 15714
rect 1181 15650 1197 15714
rect 1261 15650 1277 15714
rect 1341 15650 1357 15714
rect 1421 15650 1437 15714
rect 1501 15650 1517 15714
rect 1581 15650 1597 15714
rect 1661 15650 1677 15714
rect 1741 15650 1757 15714
rect 1821 15650 1837 15714
rect 1901 15650 1917 15714
rect 1981 15650 1997 15714
rect 2061 15650 2077 15714
rect 2141 15650 2157 15714
rect 2221 15650 2237 15714
rect 2301 15650 2317 15714
rect 2381 15650 2397 15714
rect 2461 15650 2477 15714
rect 2541 15650 2557 15714
rect 2621 15650 2637 15714
rect 2701 15650 2717 15714
rect 2781 15650 2797 15714
rect 2861 15650 2877 15714
rect 2941 15650 2957 15714
rect 3021 15650 3037 15714
rect 3101 15650 3117 15714
rect 3181 15650 3197 15714
rect 3261 15650 3277 15714
rect 3341 15650 3357 15714
rect 3421 15650 3437 15714
rect 3501 15650 3517 15714
rect 3581 15650 3597 15714
rect 3661 15650 3677 15714
rect 3741 15650 3757 15714
rect 3821 15650 3837 15714
rect 3901 15650 3917 15714
rect 3981 15650 3997 15714
rect 4061 15650 4077 15714
rect 4141 15650 4157 15714
rect 4221 15650 4237 15714
rect 4301 15650 4317 15714
rect 4381 15650 4397 15714
rect 4461 15650 4477 15714
rect 4541 15650 4557 15714
rect 4621 15650 4637 15714
rect 4701 15650 4717 15714
rect 4781 15650 4797 15714
rect 4861 15650 4899 15714
rect 119 15633 4899 15650
rect 119 15569 157 15633
rect 221 15569 237 15633
rect 301 15569 317 15633
rect 381 15569 397 15633
rect 461 15569 477 15633
rect 541 15569 557 15633
rect 621 15569 637 15633
rect 701 15569 717 15633
rect 781 15569 797 15633
rect 861 15569 877 15633
rect 941 15569 957 15633
rect 1021 15569 1037 15633
rect 1101 15569 1117 15633
rect 1181 15569 1197 15633
rect 1261 15569 1277 15633
rect 1341 15569 1357 15633
rect 1421 15569 1437 15633
rect 1501 15569 1517 15633
rect 1581 15569 1597 15633
rect 1661 15569 1677 15633
rect 1741 15569 1757 15633
rect 1821 15569 1837 15633
rect 1901 15569 1917 15633
rect 1981 15569 1997 15633
rect 2061 15569 2077 15633
rect 2141 15569 2157 15633
rect 2221 15569 2237 15633
rect 2301 15569 2317 15633
rect 2381 15569 2397 15633
rect 2461 15569 2477 15633
rect 2541 15569 2557 15633
rect 2621 15569 2637 15633
rect 2701 15569 2717 15633
rect 2781 15569 2797 15633
rect 2861 15569 2877 15633
rect 2941 15569 2957 15633
rect 3021 15569 3037 15633
rect 3101 15569 3117 15633
rect 3181 15569 3197 15633
rect 3261 15569 3277 15633
rect 3341 15569 3357 15633
rect 3421 15569 3437 15633
rect 3501 15569 3517 15633
rect 3581 15569 3597 15633
rect 3661 15569 3677 15633
rect 3741 15569 3757 15633
rect 3821 15569 3837 15633
rect 3901 15569 3917 15633
rect 3981 15569 3997 15633
rect 4061 15569 4077 15633
rect 4141 15569 4157 15633
rect 4221 15569 4237 15633
rect 4301 15569 4317 15633
rect 4381 15569 4397 15633
rect 4461 15569 4477 15633
rect 4541 15569 4557 15633
rect 4621 15569 4637 15633
rect 4701 15569 4717 15633
rect 4781 15569 4797 15633
rect 4861 15569 4899 15633
rect 119 15552 4899 15569
rect 119 15488 157 15552
rect 221 15488 237 15552
rect 301 15488 317 15552
rect 381 15488 397 15552
rect 461 15488 477 15552
rect 541 15488 557 15552
rect 621 15488 637 15552
rect 701 15488 717 15552
rect 781 15488 797 15552
rect 861 15488 877 15552
rect 941 15488 957 15552
rect 1021 15488 1037 15552
rect 1101 15488 1117 15552
rect 1181 15488 1197 15552
rect 1261 15488 1277 15552
rect 1341 15488 1357 15552
rect 1421 15488 1437 15552
rect 1501 15488 1517 15552
rect 1581 15488 1597 15552
rect 1661 15488 1677 15552
rect 1741 15488 1757 15552
rect 1821 15488 1837 15552
rect 1901 15488 1917 15552
rect 1981 15488 1997 15552
rect 2061 15488 2077 15552
rect 2141 15488 2157 15552
rect 2221 15488 2237 15552
rect 2301 15488 2317 15552
rect 2381 15488 2397 15552
rect 2461 15488 2477 15552
rect 2541 15488 2557 15552
rect 2621 15488 2637 15552
rect 2701 15488 2717 15552
rect 2781 15488 2797 15552
rect 2861 15488 2877 15552
rect 2941 15488 2957 15552
rect 3021 15488 3037 15552
rect 3101 15488 3117 15552
rect 3181 15488 3197 15552
rect 3261 15488 3277 15552
rect 3341 15488 3357 15552
rect 3421 15488 3437 15552
rect 3501 15488 3517 15552
rect 3581 15488 3597 15552
rect 3661 15488 3677 15552
rect 3741 15488 3757 15552
rect 3821 15488 3837 15552
rect 3901 15488 3917 15552
rect 3981 15488 3997 15552
rect 4061 15488 4077 15552
rect 4141 15488 4157 15552
rect 4221 15488 4237 15552
rect 4301 15488 4317 15552
rect 4381 15488 4397 15552
rect 4461 15488 4477 15552
rect 4541 15488 4557 15552
rect 4621 15488 4637 15552
rect 4701 15488 4717 15552
rect 4781 15488 4797 15552
rect 4861 15488 4899 15552
rect 119 15471 4899 15488
rect 119 15407 157 15471
rect 221 15407 237 15471
rect 301 15407 317 15471
rect 381 15407 397 15471
rect 461 15407 477 15471
rect 541 15407 557 15471
rect 621 15407 637 15471
rect 701 15407 717 15471
rect 781 15407 797 15471
rect 861 15407 877 15471
rect 941 15407 957 15471
rect 1021 15407 1037 15471
rect 1101 15407 1117 15471
rect 1181 15407 1197 15471
rect 1261 15407 1277 15471
rect 1341 15407 1357 15471
rect 1421 15407 1437 15471
rect 1501 15407 1517 15471
rect 1581 15407 1597 15471
rect 1661 15407 1677 15471
rect 1741 15407 1757 15471
rect 1821 15407 1837 15471
rect 1901 15407 1917 15471
rect 1981 15407 1997 15471
rect 2061 15407 2077 15471
rect 2141 15407 2157 15471
rect 2221 15407 2237 15471
rect 2301 15407 2317 15471
rect 2381 15407 2397 15471
rect 2461 15407 2477 15471
rect 2541 15407 2557 15471
rect 2621 15407 2637 15471
rect 2701 15407 2717 15471
rect 2781 15407 2797 15471
rect 2861 15407 2877 15471
rect 2941 15407 2957 15471
rect 3021 15407 3037 15471
rect 3101 15407 3117 15471
rect 3181 15407 3197 15471
rect 3261 15407 3277 15471
rect 3341 15407 3357 15471
rect 3421 15407 3437 15471
rect 3501 15407 3517 15471
rect 3581 15407 3597 15471
rect 3661 15407 3677 15471
rect 3741 15407 3757 15471
rect 3821 15407 3837 15471
rect 3901 15407 3917 15471
rect 3981 15407 3997 15471
rect 4061 15407 4077 15471
rect 4141 15407 4157 15471
rect 4221 15407 4237 15471
rect 4301 15407 4317 15471
rect 4381 15407 4397 15471
rect 4461 15407 4477 15471
rect 4541 15407 4557 15471
rect 4621 15407 4637 15471
rect 4701 15407 4717 15471
rect 4781 15407 4797 15471
rect 4861 15407 4899 15471
rect 119 15390 4899 15407
rect 119 15326 157 15390
rect 221 15326 237 15390
rect 301 15326 317 15390
rect 381 15326 397 15390
rect 461 15326 477 15390
rect 541 15326 557 15390
rect 621 15326 637 15390
rect 701 15326 717 15390
rect 781 15326 797 15390
rect 861 15326 877 15390
rect 941 15326 957 15390
rect 1021 15326 1037 15390
rect 1101 15326 1117 15390
rect 1181 15326 1197 15390
rect 1261 15326 1277 15390
rect 1341 15326 1357 15390
rect 1421 15326 1437 15390
rect 1501 15326 1517 15390
rect 1581 15326 1597 15390
rect 1661 15326 1677 15390
rect 1741 15326 1757 15390
rect 1821 15326 1837 15390
rect 1901 15326 1917 15390
rect 1981 15326 1997 15390
rect 2061 15326 2077 15390
rect 2141 15326 2157 15390
rect 2221 15326 2237 15390
rect 2301 15326 2317 15390
rect 2381 15326 2397 15390
rect 2461 15326 2477 15390
rect 2541 15326 2557 15390
rect 2621 15326 2637 15390
rect 2701 15326 2717 15390
rect 2781 15326 2797 15390
rect 2861 15326 2877 15390
rect 2941 15326 2957 15390
rect 3021 15326 3037 15390
rect 3101 15326 3117 15390
rect 3181 15326 3197 15390
rect 3261 15326 3277 15390
rect 3341 15326 3357 15390
rect 3421 15326 3437 15390
rect 3501 15326 3517 15390
rect 3581 15326 3597 15390
rect 3661 15326 3677 15390
rect 3741 15326 3757 15390
rect 3821 15326 3837 15390
rect 3901 15326 3917 15390
rect 3981 15326 3997 15390
rect 4061 15326 4077 15390
rect 4141 15326 4157 15390
rect 4221 15326 4237 15390
rect 4301 15326 4317 15390
rect 4381 15326 4397 15390
rect 4461 15326 4477 15390
rect 4541 15326 4557 15390
rect 4621 15326 4637 15390
rect 4701 15326 4717 15390
rect 4781 15326 4797 15390
rect 4861 15326 4899 15390
rect 119 15309 4899 15326
rect 119 15245 157 15309
rect 221 15245 237 15309
rect 301 15245 317 15309
rect 381 15245 397 15309
rect 461 15245 477 15309
rect 541 15245 557 15309
rect 621 15245 637 15309
rect 701 15245 717 15309
rect 781 15245 797 15309
rect 861 15245 877 15309
rect 941 15245 957 15309
rect 1021 15245 1037 15309
rect 1101 15245 1117 15309
rect 1181 15245 1197 15309
rect 1261 15245 1277 15309
rect 1341 15245 1357 15309
rect 1421 15245 1437 15309
rect 1501 15245 1517 15309
rect 1581 15245 1597 15309
rect 1661 15245 1677 15309
rect 1741 15245 1757 15309
rect 1821 15245 1837 15309
rect 1901 15245 1917 15309
rect 1981 15245 1997 15309
rect 2061 15245 2077 15309
rect 2141 15245 2157 15309
rect 2221 15245 2237 15309
rect 2301 15245 2317 15309
rect 2381 15245 2397 15309
rect 2461 15245 2477 15309
rect 2541 15245 2557 15309
rect 2621 15245 2637 15309
rect 2701 15245 2717 15309
rect 2781 15245 2797 15309
rect 2861 15245 2877 15309
rect 2941 15245 2957 15309
rect 3021 15245 3037 15309
rect 3101 15245 3117 15309
rect 3181 15245 3197 15309
rect 3261 15245 3277 15309
rect 3341 15245 3357 15309
rect 3421 15245 3437 15309
rect 3501 15245 3517 15309
rect 3581 15245 3597 15309
rect 3661 15245 3677 15309
rect 3741 15245 3757 15309
rect 3821 15245 3837 15309
rect 3901 15245 3917 15309
rect 3981 15245 3997 15309
rect 4061 15245 4077 15309
rect 4141 15245 4157 15309
rect 4221 15245 4237 15309
rect 4301 15245 4317 15309
rect 4381 15245 4397 15309
rect 4461 15245 4477 15309
rect 4541 15245 4557 15309
rect 4621 15245 4637 15309
rect 4701 15245 4717 15309
rect 4781 15245 4797 15309
rect 4861 15245 4899 15309
rect 119 15228 4899 15245
rect 119 15164 157 15228
rect 221 15164 237 15228
rect 301 15164 317 15228
rect 381 15164 397 15228
rect 461 15164 477 15228
rect 541 15164 557 15228
rect 621 15164 637 15228
rect 701 15164 717 15228
rect 781 15164 797 15228
rect 861 15164 877 15228
rect 941 15164 957 15228
rect 1021 15164 1037 15228
rect 1101 15164 1117 15228
rect 1181 15164 1197 15228
rect 1261 15164 1277 15228
rect 1341 15164 1357 15228
rect 1421 15164 1437 15228
rect 1501 15164 1517 15228
rect 1581 15164 1597 15228
rect 1661 15164 1677 15228
rect 1741 15164 1757 15228
rect 1821 15164 1837 15228
rect 1901 15164 1917 15228
rect 1981 15164 1997 15228
rect 2061 15164 2077 15228
rect 2141 15164 2157 15228
rect 2221 15164 2237 15228
rect 2301 15164 2317 15228
rect 2381 15164 2397 15228
rect 2461 15164 2477 15228
rect 2541 15164 2557 15228
rect 2621 15164 2637 15228
rect 2701 15164 2717 15228
rect 2781 15164 2797 15228
rect 2861 15164 2877 15228
rect 2941 15164 2957 15228
rect 3021 15164 3037 15228
rect 3101 15164 3117 15228
rect 3181 15164 3197 15228
rect 3261 15164 3277 15228
rect 3341 15164 3357 15228
rect 3421 15164 3437 15228
rect 3501 15164 3517 15228
rect 3581 15164 3597 15228
rect 3661 15164 3677 15228
rect 3741 15164 3757 15228
rect 3821 15164 3837 15228
rect 3901 15164 3917 15228
rect 3981 15164 3997 15228
rect 4061 15164 4077 15228
rect 4141 15164 4157 15228
rect 4221 15164 4237 15228
rect 4301 15164 4317 15228
rect 4381 15164 4397 15228
rect 4461 15164 4477 15228
rect 4541 15164 4557 15228
rect 4621 15164 4637 15228
rect 4701 15164 4717 15228
rect 4781 15164 4797 15228
rect 4861 15164 4899 15228
rect 119 15147 4899 15164
rect 119 15083 157 15147
rect 221 15083 237 15147
rect 301 15083 317 15147
rect 381 15083 397 15147
rect 461 15083 477 15147
rect 541 15083 557 15147
rect 621 15083 637 15147
rect 701 15083 717 15147
rect 781 15083 797 15147
rect 861 15083 877 15147
rect 941 15083 957 15147
rect 1021 15083 1037 15147
rect 1101 15083 1117 15147
rect 1181 15083 1197 15147
rect 1261 15083 1277 15147
rect 1341 15083 1357 15147
rect 1421 15083 1437 15147
rect 1501 15083 1517 15147
rect 1581 15083 1597 15147
rect 1661 15083 1677 15147
rect 1741 15083 1757 15147
rect 1821 15083 1837 15147
rect 1901 15083 1917 15147
rect 1981 15083 1997 15147
rect 2061 15083 2077 15147
rect 2141 15083 2157 15147
rect 2221 15083 2237 15147
rect 2301 15083 2317 15147
rect 2381 15083 2397 15147
rect 2461 15083 2477 15147
rect 2541 15083 2557 15147
rect 2621 15083 2637 15147
rect 2701 15083 2717 15147
rect 2781 15083 2797 15147
rect 2861 15083 2877 15147
rect 2941 15083 2957 15147
rect 3021 15083 3037 15147
rect 3101 15083 3117 15147
rect 3181 15083 3197 15147
rect 3261 15083 3277 15147
rect 3341 15083 3357 15147
rect 3421 15083 3437 15147
rect 3501 15083 3517 15147
rect 3581 15083 3597 15147
rect 3661 15083 3677 15147
rect 3741 15083 3757 15147
rect 3821 15083 3837 15147
rect 3901 15083 3917 15147
rect 3981 15083 3997 15147
rect 4061 15083 4077 15147
rect 4141 15083 4157 15147
rect 4221 15083 4237 15147
rect 4301 15083 4317 15147
rect 4381 15083 4397 15147
rect 4461 15083 4477 15147
rect 4541 15083 4557 15147
rect 4621 15083 4637 15147
rect 4701 15083 4717 15147
rect 4781 15083 4797 15147
rect 4861 15083 4899 15147
rect 119 15066 4899 15083
rect 119 15002 157 15066
rect 221 15002 237 15066
rect 301 15002 317 15066
rect 381 15002 397 15066
rect 461 15002 477 15066
rect 541 15002 557 15066
rect 621 15002 637 15066
rect 701 15002 717 15066
rect 781 15002 797 15066
rect 861 15002 877 15066
rect 941 15002 957 15066
rect 1021 15002 1037 15066
rect 1101 15002 1117 15066
rect 1181 15002 1197 15066
rect 1261 15002 1277 15066
rect 1341 15002 1357 15066
rect 1421 15002 1437 15066
rect 1501 15002 1517 15066
rect 1581 15002 1597 15066
rect 1661 15002 1677 15066
rect 1741 15002 1757 15066
rect 1821 15002 1837 15066
rect 1901 15002 1917 15066
rect 1981 15002 1997 15066
rect 2061 15002 2077 15066
rect 2141 15002 2157 15066
rect 2221 15002 2237 15066
rect 2301 15002 2317 15066
rect 2381 15002 2397 15066
rect 2461 15002 2477 15066
rect 2541 15002 2557 15066
rect 2621 15002 2637 15066
rect 2701 15002 2717 15066
rect 2781 15002 2797 15066
rect 2861 15002 2877 15066
rect 2941 15002 2957 15066
rect 3021 15002 3037 15066
rect 3101 15002 3117 15066
rect 3181 15002 3197 15066
rect 3261 15002 3277 15066
rect 3341 15002 3357 15066
rect 3421 15002 3437 15066
rect 3501 15002 3517 15066
rect 3581 15002 3597 15066
rect 3661 15002 3677 15066
rect 3741 15002 3757 15066
rect 3821 15002 3837 15066
rect 3901 15002 3917 15066
rect 3981 15002 3997 15066
rect 4061 15002 4077 15066
rect 4141 15002 4157 15066
rect 4221 15002 4237 15066
rect 4301 15002 4317 15066
rect 4381 15002 4397 15066
rect 4461 15002 4477 15066
rect 4541 15002 4557 15066
rect 4621 15002 4637 15066
rect 4701 15002 4717 15066
rect 4781 15002 4797 15066
rect 4861 15002 4899 15066
rect 119 14985 4899 15002
rect 119 14921 157 14985
rect 221 14921 237 14985
rect 301 14921 317 14985
rect 381 14921 397 14985
rect 461 14921 477 14985
rect 541 14921 557 14985
rect 621 14921 637 14985
rect 701 14921 717 14985
rect 781 14921 797 14985
rect 861 14921 877 14985
rect 941 14921 957 14985
rect 1021 14921 1037 14985
rect 1101 14921 1117 14985
rect 1181 14921 1197 14985
rect 1261 14921 1277 14985
rect 1341 14921 1357 14985
rect 1421 14921 1437 14985
rect 1501 14921 1517 14985
rect 1581 14921 1597 14985
rect 1661 14921 1677 14985
rect 1741 14921 1757 14985
rect 1821 14921 1837 14985
rect 1901 14921 1917 14985
rect 1981 14921 1997 14985
rect 2061 14921 2077 14985
rect 2141 14921 2157 14985
rect 2221 14921 2237 14985
rect 2301 14921 2317 14985
rect 2381 14921 2397 14985
rect 2461 14921 2477 14985
rect 2541 14921 2557 14985
rect 2621 14921 2637 14985
rect 2701 14921 2717 14985
rect 2781 14921 2797 14985
rect 2861 14921 2877 14985
rect 2941 14921 2957 14985
rect 3021 14921 3037 14985
rect 3101 14921 3117 14985
rect 3181 14921 3197 14985
rect 3261 14921 3277 14985
rect 3341 14921 3357 14985
rect 3421 14921 3437 14985
rect 3501 14921 3517 14985
rect 3581 14921 3597 14985
rect 3661 14921 3677 14985
rect 3741 14921 3757 14985
rect 3821 14921 3837 14985
rect 3901 14921 3917 14985
rect 3981 14921 3997 14985
rect 4061 14921 4077 14985
rect 4141 14921 4157 14985
rect 4221 14921 4237 14985
rect 4301 14921 4317 14985
rect 4381 14921 4397 14985
rect 4461 14921 4477 14985
rect 4541 14921 4557 14985
rect 4621 14921 4637 14985
rect 4701 14921 4717 14985
rect 4781 14921 4797 14985
rect 4861 14921 4899 14985
rect 119 14904 4899 14921
rect 119 14840 157 14904
rect 221 14840 237 14904
rect 301 14840 317 14904
rect 381 14840 397 14904
rect 461 14840 477 14904
rect 541 14840 557 14904
rect 621 14840 637 14904
rect 701 14840 717 14904
rect 781 14840 797 14904
rect 861 14840 877 14904
rect 941 14840 957 14904
rect 1021 14840 1037 14904
rect 1101 14840 1117 14904
rect 1181 14840 1197 14904
rect 1261 14840 1277 14904
rect 1341 14840 1357 14904
rect 1421 14840 1437 14904
rect 1501 14840 1517 14904
rect 1581 14840 1597 14904
rect 1661 14840 1677 14904
rect 1741 14840 1757 14904
rect 1821 14840 1837 14904
rect 1901 14840 1917 14904
rect 1981 14840 1997 14904
rect 2061 14840 2077 14904
rect 2141 14840 2157 14904
rect 2221 14840 2237 14904
rect 2301 14840 2317 14904
rect 2381 14840 2397 14904
rect 2461 14840 2477 14904
rect 2541 14840 2557 14904
rect 2621 14840 2637 14904
rect 2701 14840 2717 14904
rect 2781 14840 2797 14904
rect 2861 14840 2877 14904
rect 2941 14840 2957 14904
rect 3021 14840 3037 14904
rect 3101 14840 3117 14904
rect 3181 14840 3197 14904
rect 3261 14840 3277 14904
rect 3341 14840 3357 14904
rect 3421 14840 3437 14904
rect 3501 14840 3517 14904
rect 3581 14840 3597 14904
rect 3661 14840 3677 14904
rect 3741 14840 3757 14904
rect 3821 14840 3837 14904
rect 3901 14840 3917 14904
rect 3981 14840 3997 14904
rect 4061 14840 4077 14904
rect 4141 14840 4157 14904
rect 4221 14840 4237 14904
rect 4301 14840 4317 14904
rect 4381 14840 4397 14904
rect 4461 14840 4477 14904
rect 4541 14840 4557 14904
rect 4621 14840 4637 14904
rect 4701 14840 4717 14904
rect 4781 14840 4797 14904
rect 4861 14840 4899 14904
rect 119 14823 4899 14840
rect 119 14759 157 14823
rect 221 14759 237 14823
rect 301 14759 317 14823
rect 381 14759 397 14823
rect 461 14759 477 14823
rect 541 14759 557 14823
rect 621 14759 637 14823
rect 701 14759 717 14823
rect 781 14759 797 14823
rect 861 14759 877 14823
rect 941 14759 957 14823
rect 1021 14759 1037 14823
rect 1101 14759 1117 14823
rect 1181 14759 1197 14823
rect 1261 14759 1277 14823
rect 1341 14759 1357 14823
rect 1421 14759 1437 14823
rect 1501 14759 1517 14823
rect 1581 14759 1597 14823
rect 1661 14759 1677 14823
rect 1741 14759 1757 14823
rect 1821 14759 1837 14823
rect 1901 14759 1917 14823
rect 1981 14759 1997 14823
rect 2061 14759 2077 14823
rect 2141 14759 2157 14823
rect 2221 14759 2237 14823
rect 2301 14759 2317 14823
rect 2381 14759 2397 14823
rect 2461 14759 2477 14823
rect 2541 14759 2557 14823
rect 2621 14759 2637 14823
rect 2701 14759 2717 14823
rect 2781 14759 2797 14823
rect 2861 14759 2877 14823
rect 2941 14759 2957 14823
rect 3021 14759 3037 14823
rect 3101 14759 3117 14823
rect 3181 14759 3197 14823
rect 3261 14759 3277 14823
rect 3341 14759 3357 14823
rect 3421 14759 3437 14823
rect 3501 14759 3517 14823
rect 3581 14759 3597 14823
rect 3661 14759 3677 14823
rect 3741 14759 3757 14823
rect 3821 14759 3837 14823
rect 3901 14759 3917 14823
rect 3981 14759 3997 14823
rect 4061 14759 4077 14823
rect 4141 14759 4157 14823
rect 4221 14759 4237 14823
rect 4301 14759 4317 14823
rect 4381 14759 4397 14823
rect 4461 14759 4477 14823
rect 4541 14759 4557 14823
rect 4621 14759 4637 14823
rect 4701 14759 4717 14823
rect 4781 14759 4797 14823
rect 4861 14759 4899 14823
rect 119 14742 4899 14759
rect 119 14678 157 14742
rect 221 14678 237 14742
rect 301 14678 317 14742
rect 381 14678 397 14742
rect 461 14678 477 14742
rect 541 14678 557 14742
rect 621 14678 637 14742
rect 701 14678 717 14742
rect 781 14678 797 14742
rect 861 14678 877 14742
rect 941 14678 957 14742
rect 1021 14678 1037 14742
rect 1101 14678 1117 14742
rect 1181 14678 1197 14742
rect 1261 14678 1277 14742
rect 1341 14678 1357 14742
rect 1421 14678 1437 14742
rect 1501 14678 1517 14742
rect 1581 14678 1597 14742
rect 1661 14678 1677 14742
rect 1741 14678 1757 14742
rect 1821 14678 1837 14742
rect 1901 14678 1917 14742
rect 1981 14678 1997 14742
rect 2061 14678 2077 14742
rect 2141 14678 2157 14742
rect 2221 14678 2237 14742
rect 2301 14678 2317 14742
rect 2381 14678 2397 14742
rect 2461 14678 2477 14742
rect 2541 14678 2557 14742
rect 2621 14678 2637 14742
rect 2701 14678 2717 14742
rect 2781 14678 2797 14742
rect 2861 14678 2877 14742
rect 2941 14678 2957 14742
rect 3021 14678 3037 14742
rect 3101 14678 3117 14742
rect 3181 14678 3197 14742
rect 3261 14678 3277 14742
rect 3341 14678 3357 14742
rect 3421 14678 3437 14742
rect 3501 14678 3517 14742
rect 3581 14678 3597 14742
rect 3661 14678 3677 14742
rect 3741 14678 3757 14742
rect 3821 14678 3837 14742
rect 3901 14678 3917 14742
rect 3981 14678 3997 14742
rect 4061 14678 4077 14742
rect 4141 14678 4157 14742
rect 4221 14678 4237 14742
rect 4301 14678 4317 14742
rect 4381 14678 4397 14742
rect 4461 14678 4477 14742
rect 4541 14678 4557 14742
rect 4621 14678 4637 14742
rect 4701 14678 4717 14742
rect 4781 14678 4797 14742
rect 4861 14678 4899 14742
rect 119 14661 4899 14678
rect 119 14597 157 14661
rect 221 14597 237 14661
rect 301 14597 317 14661
rect 381 14597 397 14661
rect 461 14597 477 14661
rect 541 14597 557 14661
rect 621 14597 637 14661
rect 701 14597 717 14661
rect 781 14597 797 14661
rect 861 14597 877 14661
rect 941 14597 957 14661
rect 1021 14597 1037 14661
rect 1101 14597 1117 14661
rect 1181 14597 1197 14661
rect 1261 14597 1277 14661
rect 1341 14597 1357 14661
rect 1421 14597 1437 14661
rect 1501 14597 1517 14661
rect 1581 14597 1597 14661
rect 1661 14597 1677 14661
rect 1741 14597 1757 14661
rect 1821 14597 1837 14661
rect 1901 14597 1917 14661
rect 1981 14597 1997 14661
rect 2061 14597 2077 14661
rect 2141 14597 2157 14661
rect 2221 14597 2237 14661
rect 2301 14597 2317 14661
rect 2381 14597 2397 14661
rect 2461 14597 2477 14661
rect 2541 14597 2557 14661
rect 2621 14597 2637 14661
rect 2701 14597 2717 14661
rect 2781 14597 2797 14661
rect 2861 14597 2877 14661
rect 2941 14597 2957 14661
rect 3021 14597 3037 14661
rect 3101 14597 3117 14661
rect 3181 14597 3197 14661
rect 3261 14597 3277 14661
rect 3341 14597 3357 14661
rect 3421 14597 3437 14661
rect 3501 14597 3517 14661
rect 3581 14597 3597 14661
rect 3661 14597 3677 14661
rect 3741 14597 3757 14661
rect 3821 14597 3837 14661
rect 3901 14597 3917 14661
rect 3981 14597 3997 14661
rect 4061 14597 4077 14661
rect 4141 14597 4157 14661
rect 4221 14597 4237 14661
rect 4301 14597 4317 14661
rect 4381 14597 4397 14661
rect 4461 14597 4477 14661
rect 4541 14597 4557 14661
rect 4621 14597 4637 14661
rect 4701 14597 4717 14661
rect 4781 14597 4797 14661
rect 4861 14597 4899 14661
rect 119 14579 4899 14597
rect 119 14515 157 14579
rect 221 14515 237 14579
rect 301 14515 317 14579
rect 381 14515 397 14579
rect 461 14515 477 14579
rect 541 14515 557 14579
rect 621 14515 637 14579
rect 701 14515 717 14579
rect 781 14515 797 14579
rect 861 14515 877 14579
rect 941 14515 957 14579
rect 1021 14515 1037 14579
rect 1101 14515 1117 14579
rect 1181 14515 1197 14579
rect 1261 14515 1277 14579
rect 1341 14515 1357 14579
rect 1421 14515 1437 14579
rect 1501 14515 1517 14579
rect 1581 14515 1597 14579
rect 1661 14515 1677 14579
rect 1741 14515 1757 14579
rect 1821 14515 1837 14579
rect 1901 14515 1917 14579
rect 1981 14515 1997 14579
rect 2061 14515 2077 14579
rect 2141 14515 2157 14579
rect 2221 14515 2237 14579
rect 2301 14515 2317 14579
rect 2381 14515 2397 14579
rect 2461 14515 2477 14579
rect 2541 14515 2557 14579
rect 2621 14515 2637 14579
rect 2701 14515 2717 14579
rect 2781 14515 2797 14579
rect 2861 14515 2877 14579
rect 2941 14515 2957 14579
rect 3021 14515 3037 14579
rect 3101 14515 3117 14579
rect 3181 14515 3197 14579
rect 3261 14515 3277 14579
rect 3341 14515 3357 14579
rect 3421 14515 3437 14579
rect 3501 14515 3517 14579
rect 3581 14515 3597 14579
rect 3661 14515 3677 14579
rect 3741 14515 3757 14579
rect 3821 14515 3837 14579
rect 3901 14515 3917 14579
rect 3981 14515 3997 14579
rect 4061 14515 4077 14579
rect 4141 14515 4157 14579
rect 4221 14515 4237 14579
rect 4301 14515 4317 14579
rect 4381 14515 4397 14579
rect 4461 14515 4477 14579
rect 4541 14515 4557 14579
rect 4621 14515 4637 14579
rect 4701 14515 4717 14579
rect 4781 14515 4797 14579
rect 4861 14515 4899 14579
rect 119 14497 4899 14515
rect 119 14433 157 14497
rect 221 14433 237 14497
rect 301 14433 317 14497
rect 381 14433 397 14497
rect 461 14433 477 14497
rect 541 14433 557 14497
rect 621 14433 637 14497
rect 701 14433 717 14497
rect 781 14433 797 14497
rect 861 14433 877 14497
rect 941 14433 957 14497
rect 1021 14433 1037 14497
rect 1101 14433 1117 14497
rect 1181 14433 1197 14497
rect 1261 14433 1277 14497
rect 1341 14433 1357 14497
rect 1421 14433 1437 14497
rect 1501 14433 1517 14497
rect 1581 14433 1597 14497
rect 1661 14433 1677 14497
rect 1741 14433 1757 14497
rect 1821 14433 1837 14497
rect 1901 14433 1917 14497
rect 1981 14433 1997 14497
rect 2061 14433 2077 14497
rect 2141 14433 2157 14497
rect 2221 14433 2237 14497
rect 2301 14433 2317 14497
rect 2381 14433 2397 14497
rect 2461 14433 2477 14497
rect 2541 14433 2557 14497
rect 2621 14433 2637 14497
rect 2701 14433 2717 14497
rect 2781 14433 2797 14497
rect 2861 14433 2877 14497
rect 2941 14433 2957 14497
rect 3021 14433 3037 14497
rect 3101 14433 3117 14497
rect 3181 14433 3197 14497
rect 3261 14433 3277 14497
rect 3341 14433 3357 14497
rect 3421 14433 3437 14497
rect 3501 14433 3517 14497
rect 3581 14433 3597 14497
rect 3661 14433 3677 14497
rect 3741 14433 3757 14497
rect 3821 14433 3837 14497
rect 3901 14433 3917 14497
rect 3981 14433 3997 14497
rect 4061 14433 4077 14497
rect 4141 14433 4157 14497
rect 4221 14433 4237 14497
rect 4301 14433 4317 14497
rect 4381 14433 4397 14497
rect 4461 14433 4477 14497
rect 4541 14433 4557 14497
rect 4621 14433 4637 14497
rect 4701 14433 4717 14497
rect 4781 14433 4797 14497
rect 4861 14433 4899 14497
rect 119 14415 4899 14433
rect 119 14351 157 14415
rect 221 14351 237 14415
rect 301 14351 317 14415
rect 381 14351 397 14415
rect 461 14351 477 14415
rect 541 14351 557 14415
rect 621 14351 637 14415
rect 701 14351 717 14415
rect 781 14351 797 14415
rect 861 14351 877 14415
rect 941 14351 957 14415
rect 1021 14351 1037 14415
rect 1101 14351 1117 14415
rect 1181 14351 1197 14415
rect 1261 14351 1277 14415
rect 1341 14351 1357 14415
rect 1421 14351 1437 14415
rect 1501 14351 1517 14415
rect 1581 14351 1597 14415
rect 1661 14351 1677 14415
rect 1741 14351 1757 14415
rect 1821 14351 1837 14415
rect 1901 14351 1917 14415
rect 1981 14351 1997 14415
rect 2061 14351 2077 14415
rect 2141 14351 2157 14415
rect 2221 14351 2237 14415
rect 2301 14351 2317 14415
rect 2381 14351 2397 14415
rect 2461 14351 2477 14415
rect 2541 14351 2557 14415
rect 2621 14351 2637 14415
rect 2701 14351 2717 14415
rect 2781 14351 2797 14415
rect 2861 14351 2877 14415
rect 2941 14351 2957 14415
rect 3021 14351 3037 14415
rect 3101 14351 3117 14415
rect 3181 14351 3197 14415
rect 3261 14351 3277 14415
rect 3341 14351 3357 14415
rect 3421 14351 3437 14415
rect 3501 14351 3517 14415
rect 3581 14351 3597 14415
rect 3661 14351 3677 14415
rect 3741 14351 3757 14415
rect 3821 14351 3837 14415
rect 3901 14351 3917 14415
rect 3981 14351 3997 14415
rect 4061 14351 4077 14415
rect 4141 14351 4157 14415
rect 4221 14351 4237 14415
rect 4301 14351 4317 14415
rect 4381 14351 4397 14415
rect 4461 14351 4477 14415
rect 4541 14351 4557 14415
rect 4621 14351 4637 14415
rect 4701 14351 4717 14415
rect 4781 14351 4797 14415
rect 4861 14351 4899 14415
rect 119 14333 4899 14351
rect 119 14269 157 14333
rect 221 14269 237 14333
rect 301 14269 317 14333
rect 381 14269 397 14333
rect 461 14269 477 14333
rect 541 14269 557 14333
rect 621 14269 637 14333
rect 701 14269 717 14333
rect 781 14269 797 14333
rect 861 14269 877 14333
rect 941 14269 957 14333
rect 1021 14269 1037 14333
rect 1101 14269 1117 14333
rect 1181 14269 1197 14333
rect 1261 14269 1277 14333
rect 1341 14269 1357 14333
rect 1421 14269 1437 14333
rect 1501 14269 1517 14333
rect 1581 14269 1597 14333
rect 1661 14269 1677 14333
rect 1741 14269 1757 14333
rect 1821 14269 1837 14333
rect 1901 14269 1917 14333
rect 1981 14269 1997 14333
rect 2061 14269 2077 14333
rect 2141 14269 2157 14333
rect 2221 14269 2237 14333
rect 2301 14269 2317 14333
rect 2381 14269 2397 14333
rect 2461 14269 2477 14333
rect 2541 14269 2557 14333
rect 2621 14269 2637 14333
rect 2701 14269 2717 14333
rect 2781 14269 2797 14333
rect 2861 14269 2877 14333
rect 2941 14269 2957 14333
rect 3021 14269 3037 14333
rect 3101 14269 3117 14333
rect 3181 14269 3197 14333
rect 3261 14269 3277 14333
rect 3341 14269 3357 14333
rect 3421 14269 3437 14333
rect 3501 14269 3517 14333
rect 3581 14269 3597 14333
rect 3661 14269 3677 14333
rect 3741 14269 3757 14333
rect 3821 14269 3837 14333
rect 3901 14269 3917 14333
rect 3981 14269 3997 14333
rect 4061 14269 4077 14333
rect 4141 14269 4157 14333
rect 4221 14269 4237 14333
rect 4301 14269 4317 14333
rect 4381 14269 4397 14333
rect 4461 14269 4477 14333
rect 4541 14269 4557 14333
rect 4621 14269 4637 14333
rect 4701 14269 4717 14333
rect 4781 14269 4797 14333
rect 4861 14269 4899 14333
rect 119 14251 4899 14269
rect 119 14187 157 14251
rect 221 14187 237 14251
rect 301 14187 317 14251
rect 381 14187 397 14251
rect 461 14187 477 14251
rect 541 14187 557 14251
rect 621 14187 637 14251
rect 701 14187 717 14251
rect 781 14187 797 14251
rect 861 14187 877 14251
rect 941 14187 957 14251
rect 1021 14187 1037 14251
rect 1101 14187 1117 14251
rect 1181 14187 1197 14251
rect 1261 14187 1277 14251
rect 1341 14187 1357 14251
rect 1421 14187 1437 14251
rect 1501 14187 1517 14251
rect 1581 14187 1597 14251
rect 1661 14187 1677 14251
rect 1741 14187 1757 14251
rect 1821 14187 1837 14251
rect 1901 14187 1917 14251
rect 1981 14187 1997 14251
rect 2061 14187 2077 14251
rect 2141 14187 2157 14251
rect 2221 14187 2237 14251
rect 2301 14187 2317 14251
rect 2381 14187 2397 14251
rect 2461 14187 2477 14251
rect 2541 14187 2557 14251
rect 2621 14187 2637 14251
rect 2701 14187 2717 14251
rect 2781 14187 2797 14251
rect 2861 14187 2877 14251
rect 2941 14187 2957 14251
rect 3021 14187 3037 14251
rect 3101 14187 3117 14251
rect 3181 14187 3197 14251
rect 3261 14187 3277 14251
rect 3341 14187 3357 14251
rect 3421 14187 3437 14251
rect 3501 14187 3517 14251
rect 3581 14187 3597 14251
rect 3661 14187 3677 14251
rect 3741 14187 3757 14251
rect 3821 14187 3837 14251
rect 3901 14187 3917 14251
rect 3981 14187 3997 14251
rect 4061 14187 4077 14251
rect 4141 14187 4157 14251
rect 4221 14187 4237 14251
rect 4301 14187 4317 14251
rect 4381 14187 4397 14251
rect 4461 14187 4477 14251
rect 4541 14187 4557 14251
rect 4621 14187 4637 14251
rect 4701 14187 4717 14251
rect 4781 14187 4797 14251
rect 4861 14187 4899 14251
rect 119 14169 4899 14187
rect 119 14105 157 14169
rect 221 14105 237 14169
rect 301 14105 317 14169
rect 381 14105 397 14169
rect 461 14105 477 14169
rect 541 14105 557 14169
rect 621 14105 637 14169
rect 701 14105 717 14169
rect 781 14105 797 14169
rect 861 14105 877 14169
rect 941 14105 957 14169
rect 1021 14105 1037 14169
rect 1101 14105 1117 14169
rect 1181 14105 1197 14169
rect 1261 14105 1277 14169
rect 1341 14105 1357 14169
rect 1421 14105 1437 14169
rect 1501 14105 1517 14169
rect 1581 14105 1597 14169
rect 1661 14105 1677 14169
rect 1741 14105 1757 14169
rect 1821 14105 1837 14169
rect 1901 14105 1917 14169
rect 1981 14105 1997 14169
rect 2061 14105 2077 14169
rect 2141 14105 2157 14169
rect 2221 14105 2237 14169
rect 2301 14105 2317 14169
rect 2381 14105 2397 14169
rect 2461 14105 2477 14169
rect 2541 14105 2557 14169
rect 2621 14105 2637 14169
rect 2701 14105 2717 14169
rect 2781 14105 2797 14169
rect 2861 14105 2877 14169
rect 2941 14105 2957 14169
rect 3021 14105 3037 14169
rect 3101 14105 3117 14169
rect 3181 14105 3197 14169
rect 3261 14105 3277 14169
rect 3341 14105 3357 14169
rect 3421 14105 3437 14169
rect 3501 14105 3517 14169
rect 3581 14105 3597 14169
rect 3661 14105 3677 14169
rect 3741 14105 3757 14169
rect 3821 14105 3837 14169
rect 3901 14105 3917 14169
rect 3981 14105 3997 14169
rect 4061 14105 4077 14169
rect 4141 14105 4157 14169
rect 4221 14105 4237 14169
rect 4301 14105 4317 14169
rect 4381 14105 4397 14169
rect 4461 14105 4477 14169
rect 4541 14105 4557 14169
rect 4621 14105 4637 14169
rect 4701 14105 4717 14169
rect 4781 14105 4797 14169
rect 4861 14105 4899 14169
rect 119 14087 4899 14105
rect 119 14023 157 14087
rect 221 14023 237 14087
rect 301 14023 317 14087
rect 381 14023 397 14087
rect 461 14023 477 14087
rect 541 14023 557 14087
rect 621 14023 637 14087
rect 701 14023 717 14087
rect 781 14023 797 14087
rect 861 14023 877 14087
rect 941 14023 957 14087
rect 1021 14023 1037 14087
rect 1101 14023 1117 14087
rect 1181 14023 1197 14087
rect 1261 14023 1277 14087
rect 1341 14023 1357 14087
rect 1421 14023 1437 14087
rect 1501 14023 1517 14087
rect 1581 14023 1597 14087
rect 1661 14023 1677 14087
rect 1741 14023 1757 14087
rect 1821 14023 1837 14087
rect 1901 14023 1917 14087
rect 1981 14023 1997 14087
rect 2061 14023 2077 14087
rect 2141 14023 2157 14087
rect 2221 14023 2237 14087
rect 2301 14023 2317 14087
rect 2381 14023 2397 14087
rect 2461 14023 2477 14087
rect 2541 14023 2557 14087
rect 2621 14023 2637 14087
rect 2701 14023 2717 14087
rect 2781 14023 2797 14087
rect 2861 14023 2877 14087
rect 2941 14023 2957 14087
rect 3021 14023 3037 14087
rect 3101 14023 3117 14087
rect 3181 14023 3197 14087
rect 3261 14023 3277 14087
rect 3341 14023 3357 14087
rect 3421 14023 3437 14087
rect 3501 14023 3517 14087
rect 3581 14023 3597 14087
rect 3661 14023 3677 14087
rect 3741 14023 3757 14087
rect 3821 14023 3837 14087
rect 3901 14023 3917 14087
rect 3981 14023 3997 14087
rect 4061 14023 4077 14087
rect 4141 14023 4157 14087
rect 4221 14023 4237 14087
rect 4301 14023 4317 14087
rect 4381 14023 4397 14087
rect 4461 14023 4477 14087
rect 4541 14023 4557 14087
rect 4621 14023 4637 14087
rect 4701 14023 4717 14087
rect 4781 14023 4797 14087
rect 4861 14023 4899 14087
rect 119 14005 4899 14023
rect 119 13941 157 14005
rect 221 13941 237 14005
rect 301 13941 317 14005
rect 381 13941 397 14005
rect 461 13941 477 14005
rect 541 13941 557 14005
rect 621 13941 637 14005
rect 701 13941 717 14005
rect 781 13941 797 14005
rect 861 13941 877 14005
rect 941 13941 957 14005
rect 1021 13941 1037 14005
rect 1101 13941 1117 14005
rect 1181 13941 1197 14005
rect 1261 13941 1277 14005
rect 1341 13941 1357 14005
rect 1421 13941 1437 14005
rect 1501 13941 1517 14005
rect 1581 13941 1597 14005
rect 1661 13941 1677 14005
rect 1741 13941 1757 14005
rect 1821 13941 1837 14005
rect 1901 13941 1917 14005
rect 1981 13941 1997 14005
rect 2061 13941 2077 14005
rect 2141 13941 2157 14005
rect 2221 13941 2237 14005
rect 2301 13941 2317 14005
rect 2381 13941 2397 14005
rect 2461 13941 2477 14005
rect 2541 13941 2557 14005
rect 2621 13941 2637 14005
rect 2701 13941 2717 14005
rect 2781 13941 2797 14005
rect 2861 13941 2877 14005
rect 2941 13941 2957 14005
rect 3021 13941 3037 14005
rect 3101 13941 3117 14005
rect 3181 13941 3197 14005
rect 3261 13941 3277 14005
rect 3341 13941 3357 14005
rect 3421 13941 3437 14005
rect 3501 13941 3517 14005
rect 3581 13941 3597 14005
rect 3661 13941 3677 14005
rect 3741 13941 3757 14005
rect 3821 13941 3837 14005
rect 3901 13941 3917 14005
rect 3981 13941 3997 14005
rect 4061 13941 4077 14005
rect 4141 13941 4157 14005
rect 4221 13941 4237 14005
rect 4301 13941 4317 14005
rect 4381 13941 4397 14005
rect 4461 13941 4477 14005
rect 4541 13941 4557 14005
rect 4621 13941 4637 14005
rect 4701 13941 4717 14005
rect 4781 13941 4797 14005
rect 4861 13941 4899 14005
rect 119 13923 4899 13941
rect 119 13859 157 13923
rect 221 13859 237 13923
rect 301 13859 317 13923
rect 381 13859 397 13923
rect 461 13859 477 13923
rect 541 13859 557 13923
rect 621 13859 637 13923
rect 701 13859 717 13923
rect 781 13859 797 13923
rect 861 13859 877 13923
rect 941 13859 957 13923
rect 1021 13859 1037 13923
rect 1101 13859 1117 13923
rect 1181 13859 1197 13923
rect 1261 13859 1277 13923
rect 1341 13859 1357 13923
rect 1421 13859 1437 13923
rect 1501 13859 1517 13923
rect 1581 13859 1597 13923
rect 1661 13859 1677 13923
rect 1741 13859 1757 13923
rect 1821 13859 1837 13923
rect 1901 13859 1917 13923
rect 1981 13859 1997 13923
rect 2061 13859 2077 13923
rect 2141 13859 2157 13923
rect 2221 13859 2237 13923
rect 2301 13859 2317 13923
rect 2381 13859 2397 13923
rect 2461 13859 2477 13923
rect 2541 13859 2557 13923
rect 2621 13859 2637 13923
rect 2701 13859 2717 13923
rect 2781 13859 2797 13923
rect 2861 13859 2877 13923
rect 2941 13859 2957 13923
rect 3021 13859 3037 13923
rect 3101 13859 3117 13923
rect 3181 13859 3197 13923
rect 3261 13859 3277 13923
rect 3341 13859 3357 13923
rect 3421 13859 3437 13923
rect 3501 13859 3517 13923
rect 3581 13859 3597 13923
rect 3661 13859 3677 13923
rect 3741 13859 3757 13923
rect 3821 13859 3837 13923
rect 3901 13859 3917 13923
rect 3981 13859 3997 13923
rect 4061 13859 4077 13923
rect 4141 13859 4157 13923
rect 4221 13859 4237 13923
rect 4301 13859 4317 13923
rect 4381 13859 4397 13923
rect 4461 13859 4477 13923
rect 4541 13859 4557 13923
rect 4621 13859 4637 13923
rect 4701 13859 4717 13923
rect 4781 13859 4797 13923
rect 4861 13859 4899 13923
rect 119 13841 4899 13859
rect 119 13777 157 13841
rect 221 13777 237 13841
rect 301 13777 317 13841
rect 381 13777 397 13841
rect 461 13777 477 13841
rect 541 13777 557 13841
rect 621 13777 637 13841
rect 701 13777 717 13841
rect 781 13777 797 13841
rect 861 13777 877 13841
rect 941 13777 957 13841
rect 1021 13777 1037 13841
rect 1101 13777 1117 13841
rect 1181 13777 1197 13841
rect 1261 13777 1277 13841
rect 1341 13777 1357 13841
rect 1421 13777 1437 13841
rect 1501 13777 1517 13841
rect 1581 13777 1597 13841
rect 1661 13777 1677 13841
rect 1741 13777 1757 13841
rect 1821 13777 1837 13841
rect 1901 13777 1917 13841
rect 1981 13777 1997 13841
rect 2061 13777 2077 13841
rect 2141 13777 2157 13841
rect 2221 13777 2237 13841
rect 2301 13777 2317 13841
rect 2381 13777 2397 13841
rect 2461 13777 2477 13841
rect 2541 13777 2557 13841
rect 2621 13777 2637 13841
rect 2701 13777 2717 13841
rect 2781 13777 2797 13841
rect 2861 13777 2877 13841
rect 2941 13777 2957 13841
rect 3021 13777 3037 13841
rect 3101 13777 3117 13841
rect 3181 13777 3197 13841
rect 3261 13777 3277 13841
rect 3341 13777 3357 13841
rect 3421 13777 3437 13841
rect 3501 13777 3517 13841
rect 3581 13777 3597 13841
rect 3661 13777 3677 13841
rect 3741 13777 3757 13841
rect 3821 13777 3837 13841
rect 3901 13777 3917 13841
rect 3981 13777 3997 13841
rect 4061 13777 4077 13841
rect 4141 13777 4157 13841
rect 4221 13777 4237 13841
rect 4301 13777 4317 13841
rect 4381 13777 4397 13841
rect 4461 13777 4477 13841
rect 4541 13777 4557 13841
rect 4621 13777 4637 13841
rect 4701 13777 4717 13841
rect 4781 13777 4797 13841
rect 4861 13777 4899 13841
rect 119 13759 4899 13777
rect 119 13695 157 13759
rect 221 13695 237 13759
rect 301 13695 317 13759
rect 381 13695 397 13759
rect 461 13695 477 13759
rect 541 13695 557 13759
rect 621 13695 637 13759
rect 701 13695 717 13759
rect 781 13695 797 13759
rect 861 13695 877 13759
rect 941 13695 957 13759
rect 1021 13695 1037 13759
rect 1101 13695 1117 13759
rect 1181 13695 1197 13759
rect 1261 13695 1277 13759
rect 1341 13695 1357 13759
rect 1421 13695 1437 13759
rect 1501 13695 1517 13759
rect 1581 13695 1597 13759
rect 1661 13695 1677 13759
rect 1741 13695 1757 13759
rect 1821 13695 1837 13759
rect 1901 13695 1917 13759
rect 1981 13695 1997 13759
rect 2061 13695 2077 13759
rect 2141 13695 2157 13759
rect 2221 13695 2237 13759
rect 2301 13695 2317 13759
rect 2381 13695 2397 13759
rect 2461 13695 2477 13759
rect 2541 13695 2557 13759
rect 2621 13695 2637 13759
rect 2701 13695 2717 13759
rect 2781 13695 2797 13759
rect 2861 13695 2877 13759
rect 2941 13695 2957 13759
rect 3021 13695 3037 13759
rect 3101 13695 3117 13759
rect 3181 13695 3197 13759
rect 3261 13695 3277 13759
rect 3341 13695 3357 13759
rect 3421 13695 3437 13759
rect 3501 13695 3517 13759
rect 3581 13695 3597 13759
rect 3661 13695 3677 13759
rect 3741 13695 3757 13759
rect 3821 13695 3837 13759
rect 3901 13695 3917 13759
rect 3981 13695 3997 13759
rect 4061 13695 4077 13759
rect 4141 13695 4157 13759
rect 4221 13695 4237 13759
rect 4301 13695 4317 13759
rect 4381 13695 4397 13759
rect 4461 13695 4477 13759
rect 4541 13695 4557 13759
rect 4621 13695 4637 13759
rect 4701 13695 4717 13759
rect 4781 13695 4797 13759
rect 4861 13695 4899 13759
rect 119 13677 4899 13695
rect 119 13613 157 13677
rect 221 13613 237 13677
rect 301 13613 317 13677
rect 381 13613 397 13677
rect 461 13613 477 13677
rect 541 13613 557 13677
rect 621 13613 637 13677
rect 701 13613 717 13677
rect 781 13613 797 13677
rect 861 13613 877 13677
rect 941 13613 957 13677
rect 1021 13613 1037 13677
rect 1101 13613 1117 13677
rect 1181 13613 1197 13677
rect 1261 13613 1277 13677
rect 1341 13613 1357 13677
rect 1421 13613 1437 13677
rect 1501 13613 1517 13677
rect 1581 13613 1597 13677
rect 1661 13613 1677 13677
rect 1741 13613 1757 13677
rect 1821 13613 1837 13677
rect 1901 13613 1917 13677
rect 1981 13613 1997 13677
rect 2061 13613 2077 13677
rect 2141 13613 2157 13677
rect 2221 13613 2237 13677
rect 2301 13613 2317 13677
rect 2381 13613 2397 13677
rect 2461 13613 2477 13677
rect 2541 13613 2557 13677
rect 2621 13613 2637 13677
rect 2701 13613 2717 13677
rect 2781 13613 2797 13677
rect 2861 13613 2877 13677
rect 2941 13613 2957 13677
rect 3021 13613 3037 13677
rect 3101 13613 3117 13677
rect 3181 13613 3197 13677
rect 3261 13613 3277 13677
rect 3341 13613 3357 13677
rect 3421 13613 3437 13677
rect 3501 13613 3517 13677
rect 3581 13613 3597 13677
rect 3661 13613 3677 13677
rect 3741 13613 3757 13677
rect 3821 13613 3837 13677
rect 3901 13613 3917 13677
rect 3981 13613 3997 13677
rect 4061 13613 4077 13677
rect 4141 13613 4157 13677
rect 4221 13613 4237 13677
rect 4301 13613 4317 13677
rect 4381 13613 4397 13677
rect 4461 13613 4477 13677
rect 4541 13613 4557 13677
rect 4621 13613 4637 13677
rect 4701 13613 4717 13677
rect 4781 13613 4797 13677
rect 4861 13613 4899 13677
rect 119 13607 4899 13613
tri 10152 16533 10177 16558 se
rect 10177 16533 14932 16558
rect 10152 16524 14932 16533
rect 10152 16460 10190 16524
rect 10254 16460 10270 16524
rect 10334 16460 10350 16524
rect 10414 16460 10430 16524
rect 10494 16460 10510 16524
rect 10574 16460 10590 16524
rect 10654 16460 10670 16524
rect 10734 16460 10750 16524
rect 10814 16460 10830 16524
rect 10894 16460 10910 16524
rect 10974 16460 10990 16524
rect 11054 16460 11070 16524
rect 11134 16460 11150 16524
rect 11214 16460 11230 16524
rect 11294 16460 11310 16524
rect 11374 16460 11390 16524
rect 11454 16460 11470 16524
rect 11534 16460 11550 16524
rect 11614 16460 11630 16524
rect 11694 16460 11710 16524
rect 11774 16460 11790 16524
rect 11854 16460 11870 16524
rect 11934 16460 11950 16524
rect 12014 16460 12030 16524
rect 12094 16460 12110 16524
rect 12174 16460 12190 16524
rect 12254 16460 12270 16524
rect 12334 16460 12350 16524
rect 12414 16460 12430 16524
rect 12494 16460 12510 16524
rect 12574 16460 12590 16524
rect 12654 16460 12670 16524
rect 12734 16460 12750 16524
rect 12814 16460 12830 16524
rect 12894 16460 12910 16524
rect 12974 16460 12990 16524
rect 13054 16460 13070 16524
rect 13134 16460 13150 16524
rect 13214 16460 13230 16524
rect 13294 16460 13310 16524
rect 13374 16460 13390 16524
rect 13454 16460 13470 16524
rect 13534 16460 13550 16524
rect 13614 16460 13630 16524
rect 13694 16460 13710 16524
rect 13774 16460 13790 16524
rect 13854 16460 13870 16524
rect 13934 16460 13950 16524
rect 14014 16460 14030 16524
rect 14094 16460 14110 16524
rect 14174 16460 14190 16524
rect 14254 16460 14270 16524
rect 14334 16460 14350 16524
rect 14414 16460 14430 16524
rect 14494 16460 14510 16524
rect 14574 16460 14590 16524
rect 14654 16460 14670 16524
rect 14734 16460 14750 16524
rect 14814 16460 14830 16524
rect 14894 16460 14932 16524
rect 10152 16443 14932 16460
rect 10152 16379 10190 16443
rect 10254 16379 10270 16443
rect 10334 16379 10350 16443
rect 10414 16379 10430 16443
rect 10494 16379 10510 16443
rect 10574 16379 10590 16443
rect 10654 16379 10670 16443
rect 10734 16379 10750 16443
rect 10814 16379 10830 16443
rect 10894 16379 10910 16443
rect 10974 16379 10990 16443
rect 11054 16379 11070 16443
rect 11134 16379 11150 16443
rect 11214 16379 11230 16443
rect 11294 16379 11310 16443
rect 11374 16379 11390 16443
rect 11454 16379 11470 16443
rect 11534 16379 11550 16443
rect 11614 16379 11630 16443
rect 11694 16379 11710 16443
rect 11774 16379 11790 16443
rect 11854 16379 11870 16443
rect 11934 16379 11950 16443
rect 12014 16379 12030 16443
rect 12094 16379 12110 16443
rect 12174 16379 12190 16443
rect 12254 16379 12270 16443
rect 12334 16379 12350 16443
rect 12414 16379 12430 16443
rect 12494 16379 12510 16443
rect 12574 16379 12590 16443
rect 12654 16379 12670 16443
rect 12734 16379 12750 16443
rect 12814 16379 12830 16443
rect 12894 16379 12910 16443
rect 12974 16379 12990 16443
rect 13054 16379 13070 16443
rect 13134 16379 13150 16443
rect 13214 16379 13230 16443
rect 13294 16379 13310 16443
rect 13374 16379 13390 16443
rect 13454 16379 13470 16443
rect 13534 16379 13550 16443
rect 13614 16379 13630 16443
rect 13694 16379 13710 16443
rect 13774 16379 13790 16443
rect 13854 16379 13870 16443
rect 13934 16379 13950 16443
rect 14014 16379 14030 16443
rect 14094 16379 14110 16443
rect 14174 16379 14190 16443
rect 14254 16379 14270 16443
rect 14334 16379 14350 16443
rect 14414 16379 14430 16443
rect 14494 16379 14510 16443
rect 14574 16379 14590 16443
rect 14654 16379 14670 16443
rect 14734 16379 14750 16443
rect 14814 16379 14830 16443
rect 14894 16379 14932 16443
rect 10152 16362 14932 16379
rect 10152 16298 10190 16362
rect 10254 16298 10270 16362
rect 10334 16298 10350 16362
rect 10414 16298 10430 16362
rect 10494 16298 10510 16362
rect 10574 16298 10590 16362
rect 10654 16298 10670 16362
rect 10734 16298 10750 16362
rect 10814 16298 10830 16362
rect 10894 16298 10910 16362
rect 10974 16298 10990 16362
rect 11054 16298 11070 16362
rect 11134 16298 11150 16362
rect 11214 16298 11230 16362
rect 11294 16298 11310 16362
rect 11374 16298 11390 16362
rect 11454 16298 11470 16362
rect 11534 16298 11550 16362
rect 11614 16298 11630 16362
rect 11694 16298 11710 16362
rect 11774 16298 11790 16362
rect 11854 16298 11870 16362
rect 11934 16298 11950 16362
rect 12014 16298 12030 16362
rect 12094 16298 12110 16362
rect 12174 16298 12190 16362
rect 12254 16298 12270 16362
rect 12334 16298 12350 16362
rect 12414 16298 12430 16362
rect 12494 16298 12510 16362
rect 12574 16298 12590 16362
rect 12654 16298 12670 16362
rect 12734 16298 12750 16362
rect 12814 16298 12830 16362
rect 12894 16298 12910 16362
rect 12974 16298 12990 16362
rect 13054 16298 13070 16362
rect 13134 16298 13150 16362
rect 13214 16298 13230 16362
rect 13294 16298 13310 16362
rect 13374 16298 13390 16362
rect 13454 16298 13470 16362
rect 13534 16298 13550 16362
rect 13614 16298 13630 16362
rect 13694 16298 13710 16362
rect 13774 16298 13790 16362
rect 13854 16298 13870 16362
rect 13934 16298 13950 16362
rect 14014 16298 14030 16362
rect 14094 16298 14110 16362
rect 14174 16298 14190 16362
rect 14254 16298 14270 16362
rect 14334 16298 14350 16362
rect 14414 16298 14430 16362
rect 14494 16298 14510 16362
rect 14574 16298 14590 16362
rect 14654 16298 14670 16362
rect 14734 16298 14750 16362
rect 14814 16298 14830 16362
rect 14894 16298 14932 16362
rect 10152 16281 14932 16298
rect 10152 16217 10190 16281
rect 10254 16217 10270 16281
rect 10334 16217 10350 16281
rect 10414 16217 10430 16281
rect 10494 16217 10510 16281
rect 10574 16217 10590 16281
rect 10654 16217 10670 16281
rect 10734 16217 10750 16281
rect 10814 16217 10830 16281
rect 10894 16217 10910 16281
rect 10974 16217 10990 16281
rect 11054 16217 11070 16281
rect 11134 16217 11150 16281
rect 11214 16217 11230 16281
rect 11294 16217 11310 16281
rect 11374 16217 11390 16281
rect 11454 16217 11470 16281
rect 11534 16217 11550 16281
rect 11614 16217 11630 16281
rect 11694 16217 11710 16281
rect 11774 16217 11790 16281
rect 11854 16217 11870 16281
rect 11934 16217 11950 16281
rect 12014 16217 12030 16281
rect 12094 16217 12110 16281
rect 12174 16217 12190 16281
rect 12254 16217 12270 16281
rect 12334 16217 12350 16281
rect 12414 16217 12430 16281
rect 12494 16217 12510 16281
rect 12574 16217 12590 16281
rect 12654 16217 12670 16281
rect 12734 16217 12750 16281
rect 12814 16217 12830 16281
rect 12894 16217 12910 16281
rect 12974 16217 12990 16281
rect 13054 16217 13070 16281
rect 13134 16217 13150 16281
rect 13214 16217 13230 16281
rect 13294 16217 13310 16281
rect 13374 16217 13390 16281
rect 13454 16217 13470 16281
rect 13534 16217 13550 16281
rect 13614 16217 13630 16281
rect 13694 16217 13710 16281
rect 13774 16217 13790 16281
rect 13854 16217 13870 16281
rect 13934 16217 13950 16281
rect 14014 16217 14030 16281
rect 14094 16217 14110 16281
rect 14174 16217 14190 16281
rect 14254 16217 14270 16281
rect 14334 16217 14350 16281
rect 14414 16217 14430 16281
rect 14494 16217 14510 16281
rect 14574 16217 14590 16281
rect 14654 16217 14670 16281
rect 14734 16217 14750 16281
rect 14814 16217 14830 16281
rect 14894 16217 14932 16281
rect 10152 16200 14932 16217
rect 10152 16136 10190 16200
rect 10254 16136 10270 16200
rect 10334 16136 10350 16200
rect 10414 16136 10430 16200
rect 10494 16136 10510 16200
rect 10574 16136 10590 16200
rect 10654 16136 10670 16200
rect 10734 16136 10750 16200
rect 10814 16136 10830 16200
rect 10894 16136 10910 16200
rect 10974 16136 10990 16200
rect 11054 16136 11070 16200
rect 11134 16136 11150 16200
rect 11214 16136 11230 16200
rect 11294 16136 11310 16200
rect 11374 16136 11390 16200
rect 11454 16136 11470 16200
rect 11534 16136 11550 16200
rect 11614 16136 11630 16200
rect 11694 16136 11710 16200
rect 11774 16136 11790 16200
rect 11854 16136 11870 16200
rect 11934 16136 11950 16200
rect 12014 16136 12030 16200
rect 12094 16136 12110 16200
rect 12174 16136 12190 16200
rect 12254 16136 12270 16200
rect 12334 16136 12350 16200
rect 12414 16136 12430 16200
rect 12494 16136 12510 16200
rect 12574 16136 12590 16200
rect 12654 16136 12670 16200
rect 12734 16136 12750 16200
rect 12814 16136 12830 16200
rect 12894 16136 12910 16200
rect 12974 16136 12990 16200
rect 13054 16136 13070 16200
rect 13134 16136 13150 16200
rect 13214 16136 13230 16200
rect 13294 16136 13310 16200
rect 13374 16136 13390 16200
rect 13454 16136 13470 16200
rect 13534 16136 13550 16200
rect 13614 16136 13630 16200
rect 13694 16136 13710 16200
rect 13774 16136 13790 16200
rect 13854 16136 13870 16200
rect 13934 16136 13950 16200
rect 14014 16136 14030 16200
rect 14094 16136 14110 16200
rect 14174 16136 14190 16200
rect 14254 16136 14270 16200
rect 14334 16136 14350 16200
rect 14414 16136 14430 16200
rect 14494 16136 14510 16200
rect 14574 16136 14590 16200
rect 14654 16136 14670 16200
rect 14734 16136 14750 16200
rect 14814 16136 14830 16200
rect 14894 16136 14932 16200
rect 10152 16119 14932 16136
rect 10152 16055 10190 16119
rect 10254 16055 10270 16119
rect 10334 16055 10350 16119
rect 10414 16055 10430 16119
rect 10494 16055 10510 16119
rect 10574 16055 10590 16119
rect 10654 16055 10670 16119
rect 10734 16055 10750 16119
rect 10814 16055 10830 16119
rect 10894 16055 10910 16119
rect 10974 16055 10990 16119
rect 11054 16055 11070 16119
rect 11134 16055 11150 16119
rect 11214 16055 11230 16119
rect 11294 16055 11310 16119
rect 11374 16055 11390 16119
rect 11454 16055 11470 16119
rect 11534 16055 11550 16119
rect 11614 16055 11630 16119
rect 11694 16055 11710 16119
rect 11774 16055 11790 16119
rect 11854 16055 11870 16119
rect 11934 16055 11950 16119
rect 12014 16055 12030 16119
rect 12094 16055 12110 16119
rect 12174 16055 12190 16119
rect 12254 16055 12270 16119
rect 12334 16055 12350 16119
rect 12414 16055 12430 16119
rect 12494 16055 12510 16119
rect 12574 16055 12590 16119
rect 12654 16055 12670 16119
rect 12734 16055 12750 16119
rect 12814 16055 12830 16119
rect 12894 16055 12910 16119
rect 12974 16055 12990 16119
rect 13054 16055 13070 16119
rect 13134 16055 13150 16119
rect 13214 16055 13230 16119
rect 13294 16055 13310 16119
rect 13374 16055 13390 16119
rect 13454 16055 13470 16119
rect 13534 16055 13550 16119
rect 13614 16055 13630 16119
rect 13694 16055 13710 16119
rect 13774 16055 13790 16119
rect 13854 16055 13870 16119
rect 13934 16055 13950 16119
rect 14014 16055 14030 16119
rect 14094 16055 14110 16119
rect 14174 16055 14190 16119
rect 14254 16055 14270 16119
rect 14334 16055 14350 16119
rect 14414 16055 14430 16119
rect 14494 16055 14510 16119
rect 14574 16055 14590 16119
rect 14654 16055 14670 16119
rect 14734 16055 14750 16119
rect 14814 16055 14830 16119
rect 14894 16055 14932 16119
rect 10152 16038 14932 16055
rect 10152 15974 10190 16038
rect 10254 15974 10270 16038
rect 10334 15974 10350 16038
rect 10414 15974 10430 16038
rect 10494 15974 10510 16038
rect 10574 15974 10590 16038
rect 10654 15974 10670 16038
rect 10734 15974 10750 16038
rect 10814 15974 10830 16038
rect 10894 15974 10910 16038
rect 10974 15974 10990 16038
rect 11054 15974 11070 16038
rect 11134 15974 11150 16038
rect 11214 15974 11230 16038
rect 11294 15974 11310 16038
rect 11374 15974 11390 16038
rect 11454 15974 11470 16038
rect 11534 15974 11550 16038
rect 11614 15974 11630 16038
rect 11694 15974 11710 16038
rect 11774 15974 11790 16038
rect 11854 15974 11870 16038
rect 11934 15974 11950 16038
rect 12014 15974 12030 16038
rect 12094 15974 12110 16038
rect 12174 15974 12190 16038
rect 12254 15974 12270 16038
rect 12334 15974 12350 16038
rect 12414 15974 12430 16038
rect 12494 15974 12510 16038
rect 12574 15974 12590 16038
rect 12654 15974 12670 16038
rect 12734 15974 12750 16038
rect 12814 15974 12830 16038
rect 12894 15974 12910 16038
rect 12974 15974 12990 16038
rect 13054 15974 13070 16038
rect 13134 15974 13150 16038
rect 13214 15974 13230 16038
rect 13294 15974 13310 16038
rect 13374 15974 13390 16038
rect 13454 15974 13470 16038
rect 13534 15974 13550 16038
rect 13614 15974 13630 16038
rect 13694 15974 13710 16038
rect 13774 15974 13790 16038
rect 13854 15974 13870 16038
rect 13934 15974 13950 16038
rect 14014 15974 14030 16038
rect 14094 15974 14110 16038
rect 14174 15974 14190 16038
rect 14254 15974 14270 16038
rect 14334 15974 14350 16038
rect 14414 15974 14430 16038
rect 14494 15974 14510 16038
rect 14574 15974 14590 16038
rect 14654 15974 14670 16038
rect 14734 15974 14750 16038
rect 14814 15974 14830 16038
rect 14894 15974 14932 16038
rect 10152 15957 14932 15974
rect 10152 15893 10190 15957
rect 10254 15893 10270 15957
rect 10334 15893 10350 15957
rect 10414 15893 10430 15957
rect 10494 15893 10510 15957
rect 10574 15893 10590 15957
rect 10654 15893 10670 15957
rect 10734 15893 10750 15957
rect 10814 15893 10830 15957
rect 10894 15893 10910 15957
rect 10974 15893 10990 15957
rect 11054 15893 11070 15957
rect 11134 15893 11150 15957
rect 11214 15893 11230 15957
rect 11294 15893 11310 15957
rect 11374 15893 11390 15957
rect 11454 15893 11470 15957
rect 11534 15893 11550 15957
rect 11614 15893 11630 15957
rect 11694 15893 11710 15957
rect 11774 15893 11790 15957
rect 11854 15893 11870 15957
rect 11934 15893 11950 15957
rect 12014 15893 12030 15957
rect 12094 15893 12110 15957
rect 12174 15893 12190 15957
rect 12254 15893 12270 15957
rect 12334 15893 12350 15957
rect 12414 15893 12430 15957
rect 12494 15893 12510 15957
rect 12574 15893 12590 15957
rect 12654 15893 12670 15957
rect 12734 15893 12750 15957
rect 12814 15893 12830 15957
rect 12894 15893 12910 15957
rect 12974 15893 12990 15957
rect 13054 15893 13070 15957
rect 13134 15893 13150 15957
rect 13214 15893 13230 15957
rect 13294 15893 13310 15957
rect 13374 15893 13390 15957
rect 13454 15893 13470 15957
rect 13534 15893 13550 15957
rect 13614 15893 13630 15957
rect 13694 15893 13710 15957
rect 13774 15893 13790 15957
rect 13854 15893 13870 15957
rect 13934 15893 13950 15957
rect 14014 15893 14030 15957
rect 14094 15893 14110 15957
rect 14174 15893 14190 15957
rect 14254 15893 14270 15957
rect 14334 15893 14350 15957
rect 14414 15893 14430 15957
rect 14494 15893 14510 15957
rect 14574 15893 14590 15957
rect 14654 15893 14670 15957
rect 14734 15893 14750 15957
rect 14814 15893 14830 15957
rect 14894 15893 14932 15957
rect 10152 15876 14932 15893
rect 10152 15812 10190 15876
rect 10254 15812 10270 15876
rect 10334 15812 10350 15876
rect 10414 15812 10430 15876
rect 10494 15812 10510 15876
rect 10574 15812 10590 15876
rect 10654 15812 10670 15876
rect 10734 15812 10750 15876
rect 10814 15812 10830 15876
rect 10894 15812 10910 15876
rect 10974 15812 10990 15876
rect 11054 15812 11070 15876
rect 11134 15812 11150 15876
rect 11214 15812 11230 15876
rect 11294 15812 11310 15876
rect 11374 15812 11390 15876
rect 11454 15812 11470 15876
rect 11534 15812 11550 15876
rect 11614 15812 11630 15876
rect 11694 15812 11710 15876
rect 11774 15812 11790 15876
rect 11854 15812 11870 15876
rect 11934 15812 11950 15876
rect 12014 15812 12030 15876
rect 12094 15812 12110 15876
rect 12174 15812 12190 15876
rect 12254 15812 12270 15876
rect 12334 15812 12350 15876
rect 12414 15812 12430 15876
rect 12494 15812 12510 15876
rect 12574 15812 12590 15876
rect 12654 15812 12670 15876
rect 12734 15812 12750 15876
rect 12814 15812 12830 15876
rect 12894 15812 12910 15876
rect 12974 15812 12990 15876
rect 13054 15812 13070 15876
rect 13134 15812 13150 15876
rect 13214 15812 13230 15876
rect 13294 15812 13310 15876
rect 13374 15812 13390 15876
rect 13454 15812 13470 15876
rect 13534 15812 13550 15876
rect 13614 15812 13630 15876
rect 13694 15812 13710 15876
rect 13774 15812 13790 15876
rect 13854 15812 13870 15876
rect 13934 15812 13950 15876
rect 14014 15812 14030 15876
rect 14094 15812 14110 15876
rect 14174 15812 14190 15876
rect 14254 15812 14270 15876
rect 14334 15812 14350 15876
rect 14414 15812 14430 15876
rect 14494 15812 14510 15876
rect 14574 15812 14590 15876
rect 14654 15812 14670 15876
rect 14734 15812 14750 15876
rect 14814 15812 14830 15876
rect 14894 15812 14932 15876
rect 10152 15795 14932 15812
rect 10152 15731 10190 15795
rect 10254 15731 10270 15795
rect 10334 15731 10350 15795
rect 10414 15731 10430 15795
rect 10494 15731 10510 15795
rect 10574 15731 10590 15795
rect 10654 15731 10670 15795
rect 10734 15731 10750 15795
rect 10814 15731 10830 15795
rect 10894 15731 10910 15795
rect 10974 15731 10990 15795
rect 11054 15731 11070 15795
rect 11134 15731 11150 15795
rect 11214 15731 11230 15795
rect 11294 15731 11310 15795
rect 11374 15731 11390 15795
rect 11454 15731 11470 15795
rect 11534 15731 11550 15795
rect 11614 15731 11630 15795
rect 11694 15731 11710 15795
rect 11774 15731 11790 15795
rect 11854 15731 11870 15795
rect 11934 15731 11950 15795
rect 12014 15731 12030 15795
rect 12094 15731 12110 15795
rect 12174 15731 12190 15795
rect 12254 15731 12270 15795
rect 12334 15731 12350 15795
rect 12414 15731 12430 15795
rect 12494 15731 12510 15795
rect 12574 15731 12590 15795
rect 12654 15731 12670 15795
rect 12734 15731 12750 15795
rect 12814 15731 12830 15795
rect 12894 15731 12910 15795
rect 12974 15731 12990 15795
rect 13054 15731 13070 15795
rect 13134 15731 13150 15795
rect 13214 15731 13230 15795
rect 13294 15731 13310 15795
rect 13374 15731 13390 15795
rect 13454 15731 13470 15795
rect 13534 15731 13550 15795
rect 13614 15731 13630 15795
rect 13694 15731 13710 15795
rect 13774 15731 13790 15795
rect 13854 15731 13870 15795
rect 13934 15731 13950 15795
rect 14014 15731 14030 15795
rect 14094 15731 14110 15795
rect 14174 15731 14190 15795
rect 14254 15731 14270 15795
rect 14334 15731 14350 15795
rect 14414 15731 14430 15795
rect 14494 15731 14510 15795
rect 14574 15731 14590 15795
rect 14654 15731 14670 15795
rect 14734 15731 14750 15795
rect 14814 15731 14830 15795
rect 14894 15731 14932 15795
rect 10152 15714 14932 15731
rect 10152 15650 10190 15714
rect 10254 15650 10270 15714
rect 10334 15650 10350 15714
rect 10414 15650 10430 15714
rect 10494 15650 10510 15714
rect 10574 15650 10590 15714
rect 10654 15650 10670 15714
rect 10734 15650 10750 15714
rect 10814 15650 10830 15714
rect 10894 15650 10910 15714
rect 10974 15650 10990 15714
rect 11054 15650 11070 15714
rect 11134 15650 11150 15714
rect 11214 15650 11230 15714
rect 11294 15650 11310 15714
rect 11374 15650 11390 15714
rect 11454 15650 11470 15714
rect 11534 15650 11550 15714
rect 11614 15650 11630 15714
rect 11694 15650 11710 15714
rect 11774 15650 11790 15714
rect 11854 15650 11870 15714
rect 11934 15650 11950 15714
rect 12014 15650 12030 15714
rect 12094 15650 12110 15714
rect 12174 15650 12190 15714
rect 12254 15650 12270 15714
rect 12334 15650 12350 15714
rect 12414 15650 12430 15714
rect 12494 15650 12510 15714
rect 12574 15650 12590 15714
rect 12654 15650 12670 15714
rect 12734 15650 12750 15714
rect 12814 15650 12830 15714
rect 12894 15650 12910 15714
rect 12974 15650 12990 15714
rect 13054 15650 13070 15714
rect 13134 15650 13150 15714
rect 13214 15650 13230 15714
rect 13294 15650 13310 15714
rect 13374 15650 13390 15714
rect 13454 15650 13470 15714
rect 13534 15650 13550 15714
rect 13614 15650 13630 15714
rect 13694 15650 13710 15714
rect 13774 15650 13790 15714
rect 13854 15650 13870 15714
rect 13934 15650 13950 15714
rect 14014 15650 14030 15714
rect 14094 15650 14110 15714
rect 14174 15650 14190 15714
rect 14254 15650 14270 15714
rect 14334 15650 14350 15714
rect 14414 15650 14430 15714
rect 14494 15650 14510 15714
rect 14574 15650 14590 15714
rect 14654 15650 14670 15714
rect 14734 15650 14750 15714
rect 14814 15650 14830 15714
rect 14894 15650 14932 15714
rect 10152 15633 14932 15650
rect 10152 15569 10190 15633
rect 10254 15569 10270 15633
rect 10334 15569 10350 15633
rect 10414 15569 10430 15633
rect 10494 15569 10510 15633
rect 10574 15569 10590 15633
rect 10654 15569 10670 15633
rect 10734 15569 10750 15633
rect 10814 15569 10830 15633
rect 10894 15569 10910 15633
rect 10974 15569 10990 15633
rect 11054 15569 11070 15633
rect 11134 15569 11150 15633
rect 11214 15569 11230 15633
rect 11294 15569 11310 15633
rect 11374 15569 11390 15633
rect 11454 15569 11470 15633
rect 11534 15569 11550 15633
rect 11614 15569 11630 15633
rect 11694 15569 11710 15633
rect 11774 15569 11790 15633
rect 11854 15569 11870 15633
rect 11934 15569 11950 15633
rect 12014 15569 12030 15633
rect 12094 15569 12110 15633
rect 12174 15569 12190 15633
rect 12254 15569 12270 15633
rect 12334 15569 12350 15633
rect 12414 15569 12430 15633
rect 12494 15569 12510 15633
rect 12574 15569 12590 15633
rect 12654 15569 12670 15633
rect 12734 15569 12750 15633
rect 12814 15569 12830 15633
rect 12894 15569 12910 15633
rect 12974 15569 12990 15633
rect 13054 15569 13070 15633
rect 13134 15569 13150 15633
rect 13214 15569 13230 15633
rect 13294 15569 13310 15633
rect 13374 15569 13390 15633
rect 13454 15569 13470 15633
rect 13534 15569 13550 15633
rect 13614 15569 13630 15633
rect 13694 15569 13710 15633
rect 13774 15569 13790 15633
rect 13854 15569 13870 15633
rect 13934 15569 13950 15633
rect 14014 15569 14030 15633
rect 14094 15569 14110 15633
rect 14174 15569 14190 15633
rect 14254 15569 14270 15633
rect 14334 15569 14350 15633
rect 14414 15569 14430 15633
rect 14494 15569 14510 15633
rect 14574 15569 14590 15633
rect 14654 15569 14670 15633
rect 14734 15569 14750 15633
rect 14814 15569 14830 15633
rect 14894 15569 14932 15633
rect 10152 15552 14932 15569
rect 10152 15488 10190 15552
rect 10254 15488 10270 15552
rect 10334 15488 10350 15552
rect 10414 15488 10430 15552
rect 10494 15488 10510 15552
rect 10574 15488 10590 15552
rect 10654 15488 10670 15552
rect 10734 15488 10750 15552
rect 10814 15488 10830 15552
rect 10894 15488 10910 15552
rect 10974 15488 10990 15552
rect 11054 15488 11070 15552
rect 11134 15488 11150 15552
rect 11214 15488 11230 15552
rect 11294 15488 11310 15552
rect 11374 15488 11390 15552
rect 11454 15488 11470 15552
rect 11534 15488 11550 15552
rect 11614 15488 11630 15552
rect 11694 15488 11710 15552
rect 11774 15488 11790 15552
rect 11854 15488 11870 15552
rect 11934 15488 11950 15552
rect 12014 15488 12030 15552
rect 12094 15488 12110 15552
rect 12174 15488 12190 15552
rect 12254 15488 12270 15552
rect 12334 15488 12350 15552
rect 12414 15488 12430 15552
rect 12494 15488 12510 15552
rect 12574 15488 12590 15552
rect 12654 15488 12670 15552
rect 12734 15488 12750 15552
rect 12814 15488 12830 15552
rect 12894 15488 12910 15552
rect 12974 15488 12990 15552
rect 13054 15488 13070 15552
rect 13134 15488 13150 15552
rect 13214 15488 13230 15552
rect 13294 15488 13310 15552
rect 13374 15488 13390 15552
rect 13454 15488 13470 15552
rect 13534 15488 13550 15552
rect 13614 15488 13630 15552
rect 13694 15488 13710 15552
rect 13774 15488 13790 15552
rect 13854 15488 13870 15552
rect 13934 15488 13950 15552
rect 14014 15488 14030 15552
rect 14094 15488 14110 15552
rect 14174 15488 14190 15552
rect 14254 15488 14270 15552
rect 14334 15488 14350 15552
rect 14414 15488 14430 15552
rect 14494 15488 14510 15552
rect 14574 15488 14590 15552
rect 14654 15488 14670 15552
rect 14734 15488 14750 15552
rect 14814 15488 14830 15552
rect 14894 15488 14932 15552
rect 10152 15471 14932 15488
rect 10152 15407 10190 15471
rect 10254 15407 10270 15471
rect 10334 15407 10350 15471
rect 10414 15407 10430 15471
rect 10494 15407 10510 15471
rect 10574 15407 10590 15471
rect 10654 15407 10670 15471
rect 10734 15407 10750 15471
rect 10814 15407 10830 15471
rect 10894 15407 10910 15471
rect 10974 15407 10990 15471
rect 11054 15407 11070 15471
rect 11134 15407 11150 15471
rect 11214 15407 11230 15471
rect 11294 15407 11310 15471
rect 11374 15407 11390 15471
rect 11454 15407 11470 15471
rect 11534 15407 11550 15471
rect 11614 15407 11630 15471
rect 11694 15407 11710 15471
rect 11774 15407 11790 15471
rect 11854 15407 11870 15471
rect 11934 15407 11950 15471
rect 12014 15407 12030 15471
rect 12094 15407 12110 15471
rect 12174 15407 12190 15471
rect 12254 15407 12270 15471
rect 12334 15407 12350 15471
rect 12414 15407 12430 15471
rect 12494 15407 12510 15471
rect 12574 15407 12590 15471
rect 12654 15407 12670 15471
rect 12734 15407 12750 15471
rect 12814 15407 12830 15471
rect 12894 15407 12910 15471
rect 12974 15407 12990 15471
rect 13054 15407 13070 15471
rect 13134 15407 13150 15471
rect 13214 15407 13230 15471
rect 13294 15407 13310 15471
rect 13374 15407 13390 15471
rect 13454 15407 13470 15471
rect 13534 15407 13550 15471
rect 13614 15407 13630 15471
rect 13694 15407 13710 15471
rect 13774 15407 13790 15471
rect 13854 15407 13870 15471
rect 13934 15407 13950 15471
rect 14014 15407 14030 15471
rect 14094 15407 14110 15471
rect 14174 15407 14190 15471
rect 14254 15407 14270 15471
rect 14334 15407 14350 15471
rect 14414 15407 14430 15471
rect 14494 15407 14510 15471
rect 14574 15407 14590 15471
rect 14654 15407 14670 15471
rect 14734 15407 14750 15471
rect 14814 15407 14830 15471
rect 14894 15407 14932 15471
rect 10152 15390 14932 15407
rect 10152 15326 10190 15390
rect 10254 15326 10270 15390
rect 10334 15326 10350 15390
rect 10414 15326 10430 15390
rect 10494 15326 10510 15390
rect 10574 15326 10590 15390
rect 10654 15326 10670 15390
rect 10734 15326 10750 15390
rect 10814 15326 10830 15390
rect 10894 15326 10910 15390
rect 10974 15326 10990 15390
rect 11054 15326 11070 15390
rect 11134 15326 11150 15390
rect 11214 15326 11230 15390
rect 11294 15326 11310 15390
rect 11374 15326 11390 15390
rect 11454 15326 11470 15390
rect 11534 15326 11550 15390
rect 11614 15326 11630 15390
rect 11694 15326 11710 15390
rect 11774 15326 11790 15390
rect 11854 15326 11870 15390
rect 11934 15326 11950 15390
rect 12014 15326 12030 15390
rect 12094 15326 12110 15390
rect 12174 15326 12190 15390
rect 12254 15326 12270 15390
rect 12334 15326 12350 15390
rect 12414 15326 12430 15390
rect 12494 15326 12510 15390
rect 12574 15326 12590 15390
rect 12654 15326 12670 15390
rect 12734 15326 12750 15390
rect 12814 15326 12830 15390
rect 12894 15326 12910 15390
rect 12974 15326 12990 15390
rect 13054 15326 13070 15390
rect 13134 15326 13150 15390
rect 13214 15326 13230 15390
rect 13294 15326 13310 15390
rect 13374 15326 13390 15390
rect 13454 15326 13470 15390
rect 13534 15326 13550 15390
rect 13614 15326 13630 15390
rect 13694 15326 13710 15390
rect 13774 15326 13790 15390
rect 13854 15326 13870 15390
rect 13934 15326 13950 15390
rect 14014 15326 14030 15390
rect 14094 15326 14110 15390
rect 14174 15326 14190 15390
rect 14254 15326 14270 15390
rect 14334 15326 14350 15390
rect 14414 15326 14430 15390
rect 14494 15326 14510 15390
rect 14574 15326 14590 15390
rect 14654 15326 14670 15390
rect 14734 15326 14750 15390
rect 14814 15326 14830 15390
rect 14894 15326 14932 15390
rect 10152 15309 14932 15326
rect 10152 15245 10190 15309
rect 10254 15245 10270 15309
rect 10334 15245 10350 15309
rect 10414 15245 10430 15309
rect 10494 15245 10510 15309
rect 10574 15245 10590 15309
rect 10654 15245 10670 15309
rect 10734 15245 10750 15309
rect 10814 15245 10830 15309
rect 10894 15245 10910 15309
rect 10974 15245 10990 15309
rect 11054 15245 11070 15309
rect 11134 15245 11150 15309
rect 11214 15245 11230 15309
rect 11294 15245 11310 15309
rect 11374 15245 11390 15309
rect 11454 15245 11470 15309
rect 11534 15245 11550 15309
rect 11614 15245 11630 15309
rect 11694 15245 11710 15309
rect 11774 15245 11790 15309
rect 11854 15245 11870 15309
rect 11934 15245 11950 15309
rect 12014 15245 12030 15309
rect 12094 15245 12110 15309
rect 12174 15245 12190 15309
rect 12254 15245 12270 15309
rect 12334 15245 12350 15309
rect 12414 15245 12430 15309
rect 12494 15245 12510 15309
rect 12574 15245 12590 15309
rect 12654 15245 12670 15309
rect 12734 15245 12750 15309
rect 12814 15245 12830 15309
rect 12894 15245 12910 15309
rect 12974 15245 12990 15309
rect 13054 15245 13070 15309
rect 13134 15245 13150 15309
rect 13214 15245 13230 15309
rect 13294 15245 13310 15309
rect 13374 15245 13390 15309
rect 13454 15245 13470 15309
rect 13534 15245 13550 15309
rect 13614 15245 13630 15309
rect 13694 15245 13710 15309
rect 13774 15245 13790 15309
rect 13854 15245 13870 15309
rect 13934 15245 13950 15309
rect 14014 15245 14030 15309
rect 14094 15245 14110 15309
rect 14174 15245 14190 15309
rect 14254 15245 14270 15309
rect 14334 15245 14350 15309
rect 14414 15245 14430 15309
rect 14494 15245 14510 15309
rect 14574 15245 14590 15309
rect 14654 15245 14670 15309
rect 14734 15245 14750 15309
rect 14814 15245 14830 15309
rect 14894 15245 14932 15309
rect 10152 15228 14932 15245
rect 10152 15164 10190 15228
rect 10254 15164 10270 15228
rect 10334 15164 10350 15228
rect 10414 15164 10430 15228
rect 10494 15164 10510 15228
rect 10574 15164 10590 15228
rect 10654 15164 10670 15228
rect 10734 15164 10750 15228
rect 10814 15164 10830 15228
rect 10894 15164 10910 15228
rect 10974 15164 10990 15228
rect 11054 15164 11070 15228
rect 11134 15164 11150 15228
rect 11214 15164 11230 15228
rect 11294 15164 11310 15228
rect 11374 15164 11390 15228
rect 11454 15164 11470 15228
rect 11534 15164 11550 15228
rect 11614 15164 11630 15228
rect 11694 15164 11710 15228
rect 11774 15164 11790 15228
rect 11854 15164 11870 15228
rect 11934 15164 11950 15228
rect 12014 15164 12030 15228
rect 12094 15164 12110 15228
rect 12174 15164 12190 15228
rect 12254 15164 12270 15228
rect 12334 15164 12350 15228
rect 12414 15164 12430 15228
rect 12494 15164 12510 15228
rect 12574 15164 12590 15228
rect 12654 15164 12670 15228
rect 12734 15164 12750 15228
rect 12814 15164 12830 15228
rect 12894 15164 12910 15228
rect 12974 15164 12990 15228
rect 13054 15164 13070 15228
rect 13134 15164 13150 15228
rect 13214 15164 13230 15228
rect 13294 15164 13310 15228
rect 13374 15164 13390 15228
rect 13454 15164 13470 15228
rect 13534 15164 13550 15228
rect 13614 15164 13630 15228
rect 13694 15164 13710 15228
rect 13774 15164 13790 15228
rect 13854 15164 13870 15228
rect 13934 15164 13950 15228
rect 14014 15164 14030 15228
rect 14094 15164 14110 15228
rect 14174 15164 14190 15228
rect 14254 15164 14270 15228
rect 14334 15164 14350 15228
rect 14414 15164 14430 15228
rect 14494 15164 14510 15228
rect 14574 15164 14590 15228
rect 14654 15164 14670 15228
rect 14734 15164 14750 15228
rect 14814 15164 14830 15228
rect 14894 15164 14932 15228
rect 10152 15147 14932 15164
rect 10152 15083 10190 15147
rect 10254 15083 10270 15147
rect 10334 15083 10350 15147
rect 10414 15083 10430 15147
rect 10494 15083 10510 15147
rect 10574 15083 10590 15147
rect 10654 15083 10670 15147
rect 10734 15083 10750 15147
rect 10814 15083 10830 15147
rect 10894 15083 10910 15147
rect 10974 15083 10990 15147
rect 11054 15083 11070 15147
rect 11134 15083 11150 15147
rect 11214 15083 11230 15147
rect 11294 15083 11310 15147
rect 11374 15083 11390 15147
rect 11454 15083 11470 15147
rect 11534 15083 11550 15147
rect 11614 15083 11630 15147
rect 11694 15083 11710 15147
rect 11774 15083 11790 15147
rect 11854 15083 11870 15147
rect 11934 15083 11950 15147
rect 12014 15083 12030 15147
rect 12094 15083 12110 15147
rect 12174 15083 12190 15147
rect 12254 15083 12270 15147
rect 12334 15083 12350 15147
rect 12414 15083 12430 15147
rect 12494 15083 12510 15147
rect 12574 15083 12590 15147
rect 12654 15083 12670 15147
rect 12734 15083 12750 15147
rect 12814 15083 12830 15147
rect 12894 15083 12910 15147
rect 12974 15083 12990 15147
rect 13054 15083 13070 15147
rect 13134 15083 13150 15147
rect 13214 15083 13230 15147
rect 13294 15083 13310 15147
rect 13374 15083 13390 15147
rect 13454 15083 13470 15147
rect 13534 15083 13550 15147
rect 13614 15083 13630 15147
rect 13694 15083 13710 15147
rect 13774 15083 13790 15147
rect 13854 15083 13870 15147
rect 13934 15083 13950 15147
rect 14014 15083 14030 15147
rect 14094 15083 14110 15147
rect 14174 15083 14190 15147
rect 14254 15083 14270 15147
rect 14334 15083 14350 15147
rect 14414 15083 14430 15147
rect 14494 15083 14510 15147
rect 14574 15083 14590 15147
rect 14654 15083 14670 15147
rect 14734 15083 14750 15147
rect 14814 15083 14830 15147
rect 14894 15083 14932 15147
rect 10152 15066 14932 15083
rect 10152 15002 10190 15066
rect 10254 15002 10270 15066
rect 10334 15002 10350 15066
rect 10414 15002 10430 15066
rect 10494 15002 10510 15066
rect 10574 15002 10590 15066
rect 10654 15002 10670 15066
rect 10734 15002 10750 15066
rect 10814 15002 10830 15066
rect 10894 15002 10910 15066
rect 10974 15002 10990 15066
rect 11054 15002 11070 15066
rect 11134 15002 11150 15066
rect 11214 15002 11230 15066
rect 11294 15002 11310 15066
rect 11374 15002 11390 15066
rect 11454 15002 11470 15066
rect 11534 15002 11550 15066
rect 11614 15002 11630 15066
rect 11694 15002 11710 15066
rect 11774 15002 11790 15066
rect 11854 15002 11870 15066
rect 11934 15002 11950 15066
rect 12014 15002 12030 15066
rect 12094 15002 12110 15066
rect 12174 15002 12190 15066
rect 12254 15002 12270 15066
rect 12334 15002 12350 15066
rect 12414 15002 12430 15066
rect 12494 15002 12510 15066
rect 12574 15002 12590 15066
rect 12654 15002 12670 15066
rect 12734 15002 12750 15066
rect 12814 15002 12830 15066
rect 12894 15002 12910 15066
rect 12974 15002 12990 15066
rect 13054 15002 13070 15066
rect 13134 15002 13150 15066
rect 13214 15002 13230 15066
rect 13294 15002 13310 15066
rect 13374 15002 13390 15066
rect 13454 15002 13470 15066
rect 13534 15002 13550 15066
rect 13614 15002 13630 15066
rect 13694 15002 13710 15066
rect 13774 15002 13790 15066
rect 13854 15002 13870 15066
rect 13934 15002 13950 15066
rect 14014 15002 14030 15066
rect 14094 15002 14110 15066
rect 14174 15002 14190 15066
rect 14254 15002 14270 15066
rect 14334 15002 14350 15066
rect 14414 15002 14430 15066
rect 14494 15002 14510 15066
rect 14574 15002 14590 15066
rect 14654 15002 14670 15066
rect 14734 15002 14750 15066
rect 14814 15002 14830 15066
rect 14894 15002 14932 15066
rect 10152 14985 14932 15002
rect 10152 14921 10190 14985
rect 10254 14921 10270 14985
rect 10334 14921 10350 14985
rect 10414 14921 10430 14985
rect 10494 14921 10510 14985
rect 10574 14921 10590 14985
rect 10654 14921 10670 14985
rect 10734 14921 10750 14985
rect 10814 14921 10830 14985
rect 10894 14921 10910 14985
rect 10974 14921 10990 14985
rect 11054 14921 11070 14985
rect 11134 14921 11150 14985
rect 11214 14921 11230 14985
rect 11294 14921 11310 14985
rect 11374 14921 11390 14985
rect 11454 14921 11470 14985
rect 11534 14921 11550 14985
rect 11614 14921 11630 14985
rect 11694 14921 11710 14985
rect 11774 14921 11790 14985
rect 11854 14921 11870 14985
rect 11934 14921 11950 14985
rect 12014 14921 12030 14985
rect 12094 14921 12110 14985
rect 12174 14921 12190 14985
rect 12254 14921 12270 14985
rect 12334 14921 12350 14985
rect 12414 14921 12430 14985
rect 12494 14921 12510 14985
rect 12574 14921 12590 14985
rect 12654 14921 12670 14985
rect 12734 14921 12750 14985
rect 12814 14921 12830 14985
rect 12894 14921 12910 14985
rect 12974 14921 12990 14985
rect 13054 14921 13070 14985
rect 13134 14921 13150 14985
rect 13214 14921 13230 14985
rect 13294 14921 13310 14985
rect 13374 14921 13390 14985
rect 13454 14921 13470 14985
rect 13534 14921 13550 14985
rect 13614 14921 13630 14985
rect 13694 14921 13710 14985
rect 13774 14921 13790 14985
rect 13854 14921 13870 14985
rect 13934 14921 13950 14985
rect 14014 14921 14030 14985
rect 14094 14921 14110 14985
rect 14174 14921 14190 14985
rect 14254 14921 14270 14985
rect 14334 14921 14350 14985
rect 14414 14921 14430 14985
rect 14494 14921 14510 14985
rect 14574 14921 14590 14985
rect 14654 14921 14670 14985
rect 14734 14921 14750 14985
rect 14814 14921 14830 14985
rect 14894 14921 14932 14985
rect 10152 14904 14932 14921
rect 10152 14840 10190 14904
rect 10254 14840 10270 14904
rect 10334 14840 10350 14904
rect 10414 14840 10430 14904
rect 10494 14840 10510 14904
rect 10574 14840 10590 14904
rect 10654 14840 10670 14904
rect 10734 14840 10750 14904
rect 10814 14840 10830 14904
rect 10894 14840 10910 14904
rect 10974 14840 10990 14904
rect 11054 14840 11070 14904
rect 11134 14840 11150 14904
rect 11214 14840 11230 14904
rect 11294 14840 11310 14904
rect 11374 14840 11390 14904
rect 11454 14840 11470 14904
rect 11534 14840 11550 14904
rect 11614 14840 11630 14904
rect 11694 14840 11710 14904
rect 11774 14840 11790 14904
rect 11854 14840 11870 14904
rect 11934 14840 11950 14904
rect 12014 14840 12030 14904
rect 12094 14840 12110 14904
rect 12174 14840 12190 14904
rect 12254 14840 12270 14904
rect 12334 14840 12350 14904
rect 12414 14840 12430 14904
rect 12494 14840 12510 14904
rect 12574 14840 12590 14904
rect 12654 14840 12670 14904
rect 12734 14840 12750 14904
rect 12814 14840 12830 14904
rect 12894 14840 12910 14904
rect 12974 14840 12990 14904
rect 13054 14840 13070 14904
rect 13134 14840 13150 14904
rect 13214 14840 13230 14904
rect 13294 14840 13310 14904
rect 13374 14840 13390 14904
rect 13454 14840 13470 14904
rect 13534 14840 13550 14904
rect 13614 14840 13630 14904
rect 13694 14840 13710 14904
rect 13774 14840 13790 14904
rect 13854 14840 13870 14904
rect 13934 14840 13950 14904
rect 14014 14840 14030 14904
rect 14094 14840 14110 14904
rect 14174 14840 14190 14904
rect 14254 14840 14270 14904
rect 14334 14840 14350 14904
rect 14414 14840 14430 14904
rect 14494 14840 14510 14904
rect 14574 14840 14590 14904
rect 14654 14840 14670 14904
rect 14734 14840 14750 14904
rect 14814 14840 14830 14904
rect 14894 14840 14932 14904
rect 10152 14823 14932 14840
rect 10152 14759 10190 14823
rect 10254 14759 10270 14823
rect 10334 14759 10350 14823
rect 10414 14759 10430 14823
rect 10494 14759 10510 14823
rect 10574 14759 10590 14823
rect 10654 14759 10670 14823
rect 10734 14759 10750 14823
rect 10814 14759 10830 14823
rect 10894 14759 10910 14823
rect 10974 14759 10990 14823
rect 11054 14759 11070 14823
rect 11134 14759 11150 14823
rect 11214 14759 11230 14823
rect 11294 14759 11310 14823
rect 11374 14759 11390 14823
rect 11454 14759 11470 14823
rect 11534 14759 11550 14823
rect 11614 14759 11630 14823
rect 11694 14759 11710 14823
rect 11774 14759 11790 14823
rect 11854 14759 11870 14823
rect 11934 14759 11950 14823
rect 12014 14759 12030 14823
rect 12094 14759 12110 14823
rect 12174 14759 12190 14823
rect 12254 14759 12270 14823
rect 12334 14759 12350 14823
rect 12414 14759 12430 14823
rect 12494 14759 12510 14823
rect 12574 14759 12590 14823
rect 12654 14759 12670 14823
rect 12734 14759 12750 14823
rect 12814 14759 12830 14823
rect 12894 14759 12910 14823
rect 12974 14759 12990 14823
rect 13054 14759 13070 14823
rect 13134 14759 13150 14823
rect 13214 14759 13230 14823
rect 13294 14759 13310 14823
rect 13374 14759 13390 14823
rect 13454 14759 13470 14823
rect 13534 14759 13550 14823
rect 13614 14759 13630 14823
rect 13694 14759 13710 14823
rect 13774 14759 13790 14823
rect 13854 14759 13870 14823
rect 13934 14759 13950 14823
rect 14014 14759 14030 14823
rect 14094 14759 14110 14823
rect 14174 14759 14190 14823
rect 14254 14759 14270 14823
rect 14334 14759 14350 14823
rect 14414 14759 14430 14823
rect 14494 14759 14510 14823
rect 14574 14759 14590 14823
rect 14654 14759 14670 14823
rect 14734 14759 14750 14823
rect 14814 14759 14830 14823
rect 14894 14759 14932 14823
rect 10152 14742 14932 14759
rect 10152 14678 10190 14742
rect 10254 14678 10270 14742
rect 10334 14678 10350 14742
rect 10414 14678 10430 14742
rect 10494 14678 10510 14742
rect 10574 14678 10590 14742
rect 10654 14678 10670 14742
rect 10734 14678 10750 14742
rect 10814 14678 10830 14742
rect 10894 14678 10910 14742
rect 10974 14678 10990 14742
rect 11054 14678 11070 14742
rect 11134 14678 11150 14742
rect 11214 14678 11230 14742
rect 11294 14678 11310 14742
rect 11374 14678 11390 14742
rect 11454 14678 11470 14742
rect 11534 14678 11550 14742
rect 11614 14678 11630 14742
rect 11694 14678 11710 14742
rect 11774 14678 11790 14742
rect 11854 14678 11870 14742
rect 11934 14678 11950 14742
rect 12014 14678 12030 14742
rect 12094 14678 12110 14742
rect 12174 14678 12190 14742
rect 12254 14678 12270 14742
rect 12334 14678 12350 14742
rect 12414 14678 12430 14742
rect 12494 14678 12510 14742
rect 12574 14678 12590 14742
rect 12654 14678 12670 14742
rect 12734 14678 12750 14742
rect 12814 14678 12830 14742
rect 12894 14678 12910 14742
rect 12974 14678 12990 14742
rect 13054 14678 13070 14742
rect 13134 14678 13150 14742
rect 13214 14678 13230 14742
rect 13294 14678 13310 14742
rect 13374 14678 13390 14742
rect 13454 14678 13470 14742
rect 13534 14678 13550 14742
rect 13614 14678 13630 14742
rect 13694 14678 13710 14742
rect 13774 14678 13790 14742
rect 13854 14678 13870 14742
rect 13934 14678 13950 14742
rect 14014 14678 14030 14742
rect 14094 14678 14110 14742
rect 14174 14678 14190 14742
rect 14254 14678 14270 14742
rect 14334 14678 14350 14742
rect 14414 14678 14430 14742
rect 14494 14678 14510 14742
rect 14574 14678 14590 14742
rect 14654 14678 14670 14742
rect 14734 14678 14750 14742
rect 14814 14678 14830 14742
rect 14894 14678 14932 14742
rect 10152 14661 14932 14678
rect 10152 14597 10190 14661
rect 10254 14597 10270 14661
rect 10334 14597 10350 14661
rect 10414 14597 10430 14661
rect 10494 14597 10510 14661
rect 10574 14597 10590 14661
rect 10654 14597 10670 14661
rect 10734 14597 10750 14661
rect 10814 14597 10830 14661
rect 10894 14597 10910 14661
rect 10974 14597 10990 14661
rect 11054 14597 11070 14661
rect 11134 14597 11150 14661
rect 11214 14597 11230 14661
rect 11294 14597 11310 14661
rect 11374 14597 11390 14661
rect 11454 14597 11470 14661
rect 11534 14597 11550 14661
rect 11614 14597 11630 14661
rect 11694 14597 11710 14661
rect 11774 14597 11790 14661
rect 11854 14597 11870 14661
rect 11934 14597 11950 14661
rect 12014 14597 12030 14661
rect 12094 14597 12110 14661
rect 12174 14597 12190 14661
rect 12254 14597 12270 14661
rect 12334 14597 12350 14661
rect 12414 14597 12430 14661
rect 12494 14597 12510 14661
rect 12574 14597 12590 14661
rect 12654 14597 12670 14661
rect 12734 14597 12750 14661
rect 12814 14597 12830 14661
rect 12894 14597 12910 14661
rect 12974 14597 12990 14661
rect 13054 14597 13070 14661
rect 13134 14597 13150 14661
rect 13214 14597 13230 14661
rect 13294 14597 13310 14661
rect 13374 14597 13390 14661
rect 13454 14597 13470 14661
rect 13534 14597 13550 14661
rect 13614 14597 13630 14661
rect 13694 14597 13710 14661
rect 13774 14597 13790 14661
rect 13854 14597 13870 14661
rect 13934 14597 13950 14661
rect 14014 14597 14030 14661
rect 14094 14597 14110 14661
rect 14174 14597 14190 14661
rect 14254 14597 14270 14661
rect 14334 14597 14350 14661
rect 14414 14597 14430 14661
rect 14494 14597 14510 14661
rect 14574 14597 14590 14661
rect 14654 14597 14670 14661
rect 14734 14597 14750 14661
rect 14814 14597 14830 14661
rect 14894 14597 14932 14661
rect 10152 14579 14932 14597
rect 10152 14515 10190 14579
rect 10254 14515 10270 14579
rect 10334 14515 10350 14579
rect 10414 14515 10430 14579
rect 10494 14515 10510 14579
rect 10574 14515 10590 14579
rect 10654 14515 10670 14579
rect 10734 14515 10750 14579
rect 10814 14515 10830 14579
rect 10894 14515 10910 14579
rect 10974 14515 10990 14579
rect 11054 14515 11070 14579
rect 11134 14515 11150 14579
rect 11214 14515 11230 14579
rect 11294 14515 11310 14579
rect 11374 14515 11390 14579
rect 11454 14515 11470 14579
rect 11534 14515 11550 14579
rect 11614 14515 11630 14579
rect 11694 14515 11710 14579
rect 11774 14515 11790 14579
rect 11854 14515 11870 14579
rect 11934 14515 11950 14579
rect 12014 14515 12030 14579
rect 12094 14515 12110 14579
rect 12174 14515 12190 14579
rect 12254 14515 12270 14579
rect 12334 14515 12350 14579
rect 12414 14515 12430 14579
rect 12494 14515 12510 14579
rect 12574 14515 12590 14579
rect 12654 14515 12670 14579
rect 12734 14515 12750 14579
rect 12814 14515 12830 14579
rect 12894 14515 12910 14579
rect 12974 14515 12990 14579
rect 13054 14515 13070 14579
rect 13134 14515 13150 14579
rect 13214 14515 13230 14579
rect 13294 14515 13310 14579
rect 13374 14515 13390 14579
rect 13454 14515 13470 14579
rect 13534 14515 13550 14579
rect 13614 14515 13630 14579
rect 13694 14515 13710 14579
rect 13774 14515 13790 14579
rect 13854 14515 13870 14579
rect 13934 14515 13950 14579
rect 14014 14515 14030 14579
rect 14094 14515 14110 14579
rect 14174 14515 14190 14579
rect 14254 14515 14270 14579
rect 14334 14515 14350 14579
rect 14414 14515 14430 14579
rect 14494 14515 14510 14579
rect 14574 14515 14590 14579
rect 14654 14515 14670 14579
rect 14734 14515 14750 14579
rect 14814 14515 14830 14579
rect 14894 14515 14932 14579
rect 10152 14497 14932 14515
rect 10152 14433 10190 14497
rect 10254 14433 10270 14497
rect 10334 14433 10350 14497
rect 10414 14433 10430 14497
rect 10494 14433 10510 14497
rect 10574 14433 10590 14497
rect 10654 14433 10670 14497
rect 10734 14433 10750 14497
rect 10814 14433 10830 14497
rect 10894 14433 10910 14497
rect 10974 14433 10990 14497
rect 11054 14433 11070 14497
rect 11134 14433 11150 14497
rect 11214 14433 11230 14497
rect 11294 14433 11310 14497
rect 11374 14433 11390 14497
rect 11454 14433 11470 14497
rect 11534 14433 11550 14497
rect 11614 14433 11630 14497
rect 11694 14433 11710 14497
rect 11774 14433 11790 14497
rect 11854 14433 11870 14497
rect 11934 14433 11950 14497
rect 12014 14433 12030 14497
rect 12094 14433 12110 14497
rect 12174 14433 12190 14497
rect 12254 14433 12270 14497
rect 12334 14433 12350 14497
rect 12414 14433 12430 14497
rect 12494 14433 12510 14497
rect 12574 14433 12590 14497
rect 12654 14433 12670 14497
rect 12734 14433 12750 14497
rect 12814 14433 12830 14497
rect 12894 14433 12910 14497
rect 12974 14433 12990 14497
rect 13054 14433 13070 14497
rect 13134 14433 13150 14497
rect 13214 14433 13230 14497
rect 13294 14433 13310 14497
rect 13374 14433 13390 14497
rect 13454 14433 13470 14497
rect 13534 14433 13550 14497
rect 13614 14433 13630 14497
rect 13694 14433 13710 14497
rect 13774 14433 13790 14497
rect 13854 14433 13870 14497
rect 13934 14433 13950 14497
rect 14014 14433 14030 14497
rect 14094 14433 14110 14497
rect 14174 14433 14190 14497
rect 14254 14433 14270 14497
rect 14334 14433 14350 14497
rect 14414 14433 14430 14497
rect 14494 14433 14510 14497
rect 14574 14433 14590 14497
rect 14654 14433 14670 14497
rect 14734 14433 14750 14497
rect 14814 14433 14830 14497
rect 14894 14433 14932 14497
rect 10152 14415 14932 14433
rect 10152 14351 10190 14415
rect 10254 14351 10270 14415
rect 10334 14351 10350 14415
rect 10414 14351 10430 14415
rect 10494 14351 10510 14415
rect 10574 14351 10590 14415
rect 10654 14351 10670 14415
rect 10734 14351 10750 14415
rect 10814 14351 10830 14415
rect 10894 14351 10910 14415
rect 10974 14351 10990 14415
rect 11054 14351 11070 14415
rect 11134 14351 11150 14415
rect 11214 14351 11230 14415
rect 11294 14351 11310 14415
rect 11374 14351 11390 14415
rect 11454 14351 11470 14415
rect 11534 14351 11550 14415
rect 11614 14351 11630 14415
rect 11694 14351 11710 14415
rect 11774 14351 11790 14415
rect 11854 14351 11870 14415
rect 11934 14351 11950 14415
rect 12014 14351 12030 14415
rect 12094 14351 12110 14415
rect 12174 14351 12190 14415
rect 12254 14351 12270 14415
rect 12334 14351 12350 14415
rect 12414 14351 12430 14415
rect 12494 14351 12510 14415
rect 12574 14351 12590 14415
rect 12654 14351 12670 14415
rect 12734 14351 12750 14415
rect 12814 14351 12830 14415
rect 12894 14351 12910 14415
rect 12974 14351 12990 14415
rect 13054 14351 13070 14415
rect 13134 14351 13150 14415
rect 13214 14351 13230 14415
rect 13294 14351 13310 14415
rect 13374 14351 13390 14415
rect 13454 14351 13470 14415
rect 13534 14351 13550 14415
rect 13614 14351 13630 14415
rect 13694 14351 13710 14415
rect 13774 14351 13790 14415
rect 13854 14351 13870 14415
rect 13934 14351 13950 14415
rect 14014 14351 14030 14415
rect 14094 14351 14110 14415
rect 14174 14351 14190 14415
rect 14254 14351 14270 14415
rect 14334 14351 14350 14415
rect 14414 14351 14430 14415
rect 14494 14351 14510 14415
rect 14574 14351 14590 14415
rect 14654 14351 14670 14415
rect 14734 14351 14750 14415
rect 14814 14351 14830 14415
rect 14894 14351 14932 14415
rect 10152 14333 14932 14351
rect 10152 14269 10190 14333
rect 10254 14269 10270 14333
rect 10334 14269 10350 14333
rect 10414 14269 10430 14333
rect 10494 14269 10510 14333
rect 10574 14269 10590 14333
rect 10654 14269 10670 14333
rect 10734 14269 10750 14333
rect 10814 14269 10830 14333
rect 10894 14269 10910 14333
rect 10974 14269 10990 14333
rect 11054 14269 11070 14333
rect 11134 14269 11150 14333
rect 11214 14269 11230 14333
rect 11294 14269 11310 14333
rect 11374 14269 11390 14333
rect 11454 14269 11470 14333
rect 11534 14269 11550 14333
rect 11614 14269 11630 14333
rect 11694 14269 11710 14333
rect 11774 14269 11790 14333
rect 11854 14269 11870 14333
rect 11934 14269 11950 14333
rect 12014 14269 12030 14333
rect 12094 14269 12110 14333
rect 12174 14269 12190 14333
rect 12254 14269 12270 14333
rect 12334 14269 12350 14333
rect 12414 14269 12430 14333
rect 12494 14269 12510 14333
rect 12574 14269 12590 14333
rect 12654 14269 12670 14333
rect 12734 14269 12750 14333
rect 12814 14269 12830 14333
rect 12894 14269 12910 14333
rect 12974 14269 12990 14333
rect 13054 14269 13070 14333
rect 13134 14269 13150 14333
rect 13214 14269 13230 14333
rect 13294 14269 13310 14333
rect 13374 14269 13390 14333
rect 13454 14269 13470 14333
rect 13534 14269 13550 14333
rect 13614 14269 13630 14333
rect 13694 14269 13710 14333
rect 13774 14269 13790 14333
rect 13854 14269 13870 14333
rect 13934 14269 13950 14333
rect 14014 14269 14030 14333
rect 14094 14269 14110 14333
rect 14174 14269 14190 14333
rect 14254 14269 14270 14333
rect 14334 14269 14350 14333
rect 14414 14269 14430 14333
rect 14494 14269 14510 14333
rect 14574 14269 14590 14333
rect 14654 14269 14670 14333
rect 14734 14269 14750 14333
rect 14814 14269 14830 14333
rect 14894 14269 14932 14333
rect 10152 14251 14932 14269
rect 10152 14187 10190 14251
rect 10254 14187 10270 14251
rect 10334 14187 10350 14251
rect 10414 14187 10430 14251
rect 10494 14187 10510 14251
rect 10574 14187 10590 14251
rect 10654 14187 10670 14251
rect 10734 14187 10750 14251
rect 10814 14187 10830 14251
rect 10894 14187 10910 14251
rect 10974 14187 10990 14251
rect 11054 14187 11070 14251
rect 11134 14187 11150 14251
rect 11214 14187 11230 14251
rect 11294 14187 11310 14251
rect 11374 14187 11390 14251
rect 11454 14187 11470 14251
rect 11534 14187 11550 14251
rect 11614 14187 11630 14251
rect 11694 14187 11710 14251
rect 11774 14187 11790 14251
rect 11854 14187 11870 14251
rect 11934 14187 11950 14251
rect 12014 14187 12030 14251
rect 12094 14187 12110 14251
rect 12174 14187 12190 14251
rect 12254 14187 12270 14251
rect 12334 14187 12350 14251
rect 12414 14187 12430 14251
rect 12494 14187 12510 14251
rect 12574 14187 12590 14251
rect 12654 14187 12670 14251
rect 12734 14187 12750 14251
rect 12814 14187 12830 14251
rect 12894 14187 12910 14251
rect 12974 14187 12990 14251
rect 13054 14187 13070 14251
rect 13134 14187 13150 14251
rect 13214 14187 13230 14251
rect 13294 14187 13310 14251
rect 13374 14187 13390 14251
rect 13454 14187 13470 14251
rect 13534 14187 13550 14251
rect 13614 14187 13630 14251
rect 13694 14187 13710 14251
rect 13774 14187 13790 14251
rect 13854 14187 13870 14251
rect 13934 14187 13950 14251
rect 14014 14187 14030 14251
rect 14094 14187 14110 14251
rect 14174 14187 14190 14251
rect 14254 14187 14270 14251
rect 14334 14187 14350 14251
rect 14414 14187 14430 14251
rect 14494 14187 14510 14251
rect 14574 14187 14590 14251
rect 14654 14187 14670 14251
rect 14734 14187 14750 14251
rect 14814 14187 14830 14251
rect 14894 14187 14932 14251
rect 10152 14169 14932 14187
rect 10152 14105 10190 14169
rect 10254 14105 10270 14169
rect 10334 14105 10350 14169
rect 10414 14105 10430 14169
rect 10494 14105 10510 14169
rect 10574 14105 10590 14169
rect 10654 14105 10670 14169
rect 10734 14105 10750 14169
rect 10814 14105 10830 14169
rect 10894 14105 10910 14169
rect 10974 14105 10990 14169
rect 11054 14105 11070 14169
rect 11134 14105 11150 14169
rect 11214 14105 11230 14169
rect 11294 14105 11310 14169
rect 11374 14105 11390 14169
rect 11454 14105 11470 14169
rect 11534 14105 11550 14169
rect 11614 14105 11630 14169
rect 11694 14105 11710 14169
rect 11774 14105 11790 14169
rect 11854 14105 11870 14169
rect 11934 14105 11950 14169
rect 12014 14105 12030 14169
rect 12094 14105 12110 14169
rect 12174 14105 12190 14169
rect 12254 14105 12270 14169
rect 12334 14105 12350 14169
rect 12414 14105 12430 14169
rect 12494 14105 12510 14169
rect 12574 14105 12590 14169
rect 12654 14105 12670 14169
rect 12734 14105 12750 14169
rect 12814 14105 12830 14169
rect 12894 14105 12910 14169
rect 12974 14105 12990 14169
rect 13054 14105 13070 14169
rect 13134 14105 13150 14169
rect 13214 14105 13230 14169
rect 13294 14105 13310 14169
rect 13374 14105 13390 14169
rect 13454 14105 13470 14169
rect 13534 14105 13550 14169
rect 13614 14105 13630 14169
rect 13694 14105 13710 14169
rect 13774 14105 13790 14169
rect 13854 14105 13870 14169
rect 13934 14105 13950 14169
rect 14014 14105 14030 14169
rect 14094 14105 14110 14169
rect 14174 14105 14190 14169
rect 14254 14105 14270 14169
rect 14334 14105 14350 14169
rect 14414 14105 14430 14169
rect 14494 14105 14510 14169
rect 14574 14105 14590 14169
rect 14654 14105 14670 14169
rect 14734 14105 14750 14169
rect 14814 14105 14830 14169
rect 14894 14105 14932 14169
rect 10152 14087 14932 14105
rect 10152 14023 10190 14087
rect 10254 14023 10270 14087
rect 10334 14023 10350 14087
rect 10414 14023 10430 14087
rect 10494 14023 10510 14087
rect 10574 14023 10590 14087
rect 10654 14023 10670 14087
rect 10734 14023 10750 14087
rect 10814 14023 10830 14087
rect 10894 14023 10910 14087
rect 10974 14023 10990 14087
rect 11054 14023 11070 14087
rect 11134 14023 11150 14087
rect 11214 14023 11230 14087
rect 11294 14023 11310 14087
rect 11374 14023 11390 14087
rect 11454 14023 11470 14087
rect 11534 14023 11550 14087
rect 11614 14023 11630 14087
rect 11694 14023 11710 14087
rect 11774 14023 11790 14087
rect 11854 14023 11870 14087
rect 11934 14023 11950 14087
rect 12014 14023 12030 14087
rect 12094 14023 12110 14087
rect 12174 14023 12190 14087
rect 12254 14023 12270 14087
rect 12334 14023 12350 14087
rect 12414 14023 12430 14087
rect 12494 14023 12510 14087
rect 12574 14023 12590 14087
rect 12654 14023 12670 14087
rect 12734 14023 12750 14087
rect 12814 14023 12830 14087
rect 12894 14023 12910 14087
rect 12974 14023 12990 14087
rect 13054 14023 13070 14087
rect 13134 14023 13150 14087
rect 13214 14023 13230 14087
rect 13294 14023 13310 14087
rect 13374 14023 13390 14087
rect 13454 14023 13470 14087
rect 13534 14023 13550 14087
rect 13614 14023 13630 14087
rect 13694 14023 13710 14087
rect 13774 14023 13790 14087
rect 13854 14023 13870 14087
rect 13934 14023 13950 14087
rect 14014 14023 14030 14087
rect 14094 14023 14110 14087
rect 14174 14023 14190 14087
rect 14254 14023 14270 14087
rect 14334 14023 14350 14087
rect 14414 14023 14430 14087
rect 14494 14023 14510 14087
rect 14574 14023 14590 14087
rect 14654 14023 14670 14087
rect 14734 14023 14750 14087
rect 14814 14023 14830 14087
rect 14894 14023 14932 14087
rect 10152 14005 14932 14023
rect 10152 13941 10190 14005
rect 10254 13941 10270 14005
rect 10334 13941 10350 14005
rect 10414 13941 10430 14005
rect 10494 13941 10510 14005
rect 10574 13941 10590 14005
rect 10654 13941 10670 14005
rect 10734 13941 10750 14005
rect 10814 13941 10830 14005
rect 10894 13941 10910 14005
rect 10974 13941 10990 14005
rect 11054 13941 11070 14005
rect 11134 13941 11150 14005
rect 11214 13941 11230 14005
rect 11294 13941 11310 14005
rect 11374 13941 11390 14005
rect 11454 13941 11470 14005
rect 11534 13941 11550 14005
rect 11614 13941 11630 14005
rect 11694 13941 11710 14005
rect 11774 13941 11790 14005
rect 11854 13941 11870 14005
rect 11934 13941 11950 14005
rect 12014 13941 12030 14005
rect 12094 13941 12110 14005
rect 12174 13941 12190 14005
rect 12254 13941 12270 14005
rect 12334 13941 12350 14005
rect 12414 13941 12430 14005
rect 12494 13941 12510 14005
rect 12574 13941 12590 14005
rect 12654 13941 12670 14005
rect 12734 13941 12750 14005
rect 12814 13941 12830 14005
rect 12894 13941 12910 14005
rect 12974 13941 12990 14005
rect 13054 13941 13070 14005
rect 13134 13941 13150 14005
rect 13214 13941 13230 14005
rect 13294 13941 13310 14005
rect 13374 13941 13390 14005
rect 13454 13941 13470 14005
rect 13534 13941 13550 14005
rect 13614 13941 13630 14005
rect 13694 13941 13710 14005
rect 13774 13941 13790 14005
rect 13854 13941 13870 14005
rect 13934 13941 13950 14005
rect 14014 13941 14030 14005
rect 14094 13941 14110 14005
rect 14174 13941 14190 14005
rect 14254 13941 14270 14005
rect 14334 13941 14350 14005
rect 14414 13941 14430 14005
rect 14494 13941 14510 14005
rect 14574 13941 14590 14005
rect 14654 13941 14670 14005
rect 14734 13941 14750 14005
rect 14814 13941 14830 14005
rect 14894 13941 14932 14005
rect 10152 13923 14932 13941
rect 10152 13859 10190 13923
rect 10254 13859 10270 13923
rect 10334 13859 10350 13923
rect 10414 13859 10430 13923
rect 10494 13859 10510 13923
rect 10574 13859 10590 13923
rect 10654 13859 10670 13923
rect 10734 13859 10750 13923
rect 10814 13859 10830 13923
rect 10894 13859 10910 13923
rect 10974 13859 10990 13923
rect 11054 13859 11070 13923
rect 11134 13859 11150 13923
rect 11214 13859 11230 13923
rect 11294 13859 11310 13923
rect 11374 13859 11390 13923
rect 11454 13859 11470 13923
rect 11534 13859 11550 13923
rect 11614 13859 11630 13923
rect 11694 13859 11710 13923
rect 11774 13859 11790 13923
rect 11854 13859 11870 13923
rect 11934 13859 11950 13923
rect 12014 13859 12030 13923
rect 12094 13859 12110 13923
rect 12174 13859 12190 13923
rect 12254 13859 12270 13923
rect 12334 13859 12350 13923
rect 12414 13859 12430 13923
rect 12494 13859 12510 13923
rect 12574 13859 12590 13923
rect 12654 13859 12670 13923
rect 12734 13859 12750 13923
rect 12814 13859 12830 13923
rect 12894 13859 12910 13923
rect 12974 13859 12990 13923
rect 13054 13859 13070 13923
rect 13134 13859 13150 13923
rect 13214 13859 13230 13923
rect 13294 13859 13310 13923
rect 13374 13859 13390 13923
rect 13454 13859 13470 13923
rect 13534 13859 13550 13923
rect 13614 13859 13630 13923
rect 13694 13859 13710 13923
rect 13774 13859 13790 13923
rect 13854 13859 13870 13923
rect 13934 13859 13950 13923
rect 14014 13859 14030 13923
rect 14094 13859 14110 13923
rect 14174 13859 14190 13923
rect 14254 13859 14270 13923
rect 14334 13859 14350 13923
rect 14414 13859 14430 13923
rect 14494 13859 14510 13923
rect 14574 13859 14590 13923
rect 14654 13859 14670 13923
rect 14734 13859 14750 13923
rect 14814 13859 14830 13923
rect 14894 13859 14932 13923
rect 10152 13841 14932 13859
rect 10152 13777 10190 13841
rect 10254 13777 10270 13841
rect 10334 13777 10350 13841
rect 10414 13777 10430 13841
rect 10494 13777 10510 13841
rect 10574 13777 10590 13841
rect 10654 13777 10670 13841
rect 10734 13777 10750 13841
rect 10814 13777 10830 13841
rect 10894 13777 10910 13841
rect 10974 13777 10990 13841
rect 11054 13777 11070 13841
rect 11134 13777 11150 13841
rect 11214 13777 11230 13841
rect 11294 13777 11310 13841
rect 11374 13777 11390 13841
rect 11454 13777 11470 13841
rect 11534 13777 11550 13841
rect 11614 13777 11630 13841
rect 11694 13777 11710 13841
rect 11774 13777 11790 13841
rect 11854 13777 11870 13841
rect 11934 13777 11950 13841
rect 12014 13777 12030 13841
rect 12094 13777 12110 13841
rect 12174 13777 12190 13841
rect 12254 13777 12270 13841
rect 12334 13777 12350 13841
rect 12414 13777 12430 13841
rect 12494 13777 12510 13841
rect 12574 13777 12590 13841
rect 12654 13777 12670 13841
rect 12734 13777 12750 13841
rect 12814 13777 12830 13841
rect 12894 13777 12910 13841
rect 12974 13777 12990 13841
rect 13054 13777 13070 13841
rect 13134 13777 13150 13841
rect 13214 13777 13230 13841
rect 13294 13777 13310 13841
rect 13374 13777 13390 13841
rect 13454 13777 13470 13841
rect 13534 13777 13550 13841
rect 13614 13777 13630 13841
rect 13694 13777 13710 13841
rect 13774 13777 13790 13841
rect 13854 13777 13870 13841
rect 13934 13777 13950 13841
rect 14014 13777 14030 13841
rect 14094 13777 14110 13841
rect 14174 13777 14190 13841
rect 14254 13777 14270 13841
rect 14334 13777 14350 13841
rect 14414 13777 14430 13841
rect 14494 13777 14510 13841
rect 14574 13777 14590 13841
rect 14654 13777 14670 13841
rect 14734 13777 14750 13841
rect 14814 13777 14830 13841
rect 14894 13777 14932 13841
rect 10152 13759 14932 13777
rect 10152 13695 10190 13759
rect 10254 13695 10270 13759
rect 10334 13695 10350 13759
rect 10414 13695 10430 13759
rect 10494 13695 10510 13759
rect 10574 13695 10590 13759
rect 10654 13695 10670 13759
rect 10734 13695 10750 13759
rect 10814 13695 10830 13759
rect 10894 13695 10910 13759
rect 10974 13695 10990 13759
rect 11054 13695 11070 13759
rect 11134 13695 11150 13759
rect 11214 13695 11230 13759
rect 11294 13695 11310 13759
rect 11374 13695 11390 13759
rect 11454 13695 11470 13759
rect 11534 13695 11550 13759
rect 11614 13695 11630 13759
rect 11694 13695 11710 13759
rect 11774 13695 11790 13759
rect 11854 13695 11870 13759
rect 11934 13695 11950 13759
rect 12014 13695 12030 13759
rect 12094 13695 12110 13759
rect 12174 13695 12190 13759
rect 12254 13695 12270 13759
rect 12334 13695 12350 13759
rect 12414 13695 12430 13759
rect 12494 13695 12510 13759
rect 12574 13695 12590 13759
rect 12654 13695 12670 13759
rect 12734 13695 12750 13759
rect 12814 13695 12830 13759
rect 12894 13695 12910 13759
rect 12974 13695 12990 13759
rect 13054 13695 13070 13759
rect 13134 13695 13150 13759
rect 13214 13695 13230 13759
rect 13294 13695 13310 13759
rect 13374 13695 13390 13759
rect 13454 13695 13470 13759
rect 13534 13695 13550 13759
rect 13614 13695 13630 13759
rect 13694 13695 13710 13759
rect 13774 13695 13790 13759
rect 13854 13695 13870 13759
rect 13934 13695 13950 13759
rect 14014 13695 14030 13759
rect 14094 13695 14110 13759
rect 14174 13695 14190 13759
rect 14254 13695 14270 13759
rect 14334 13695 14350 13759
rect 14414 13695 14430 13759
rect 14494 13695 14510 13759
rect 14574 13695 14590 13759
rect 14654 13695 14670 13759
rect 14734 13695 14750 13759
rect 14814 13695 14830 13759
rect 14894 13695 14932 13759
rect 10152 13677 14932 13695
rect 10152 13613 10190 13677
rect 10254 13613 10270 13677
rect 10334 13613 10350 13677
rect 10414 13613 10430 13677
rect 10494 13613 10510 13677
rect 10574 13613 10590 13677
rect 10654 13613 10670 13677
rect 10734 13613 10750 13677
rect 10814 13613 10830 13677
rect 10894 13613 10910 13677
rect 10974 13613 10990 13677
rect 11054 13613 11070 13677
rect 11134 13613 11150 13677
rect 11214 13613 11230 13677
rect 11294 13613 11310 13677
rect 11374 13613 11390 13677
rect 11454 13613 11470 13677
rect 11534 13613 11550 13677
rect 11614 13613 11630 13677
rect 11694 13613 11710 13677
rect 11774 13613 11790 13677
rect 11854 13613 11870 13677
rect 11934 13613 11950 13677
rect 12014 13613 12030 13677
rect 12094 13613 12110 13677
rect 12174 13613 12190 13677
rect 12254 13613 12270 13677
rect 12334 13613 12350 13677
rect 12414 13613 12430 13677
rect 12494 13613 12510 13677
rect 12574 13613 12590 13677
rect 12654 13613 12670 13677
rect 12734 13613 12750 13677
rect 12814 13613 12830 13677
rect 12894 13613 12910 13677
rect 12974 13613 12990 13677
rect 13054 13613 13070 13677
rect 13134 13613 13150 13677
rect 13214 13613 13230 13677
rect 13294 13613 13310 13677
rect 13374 13613 13390 13677
rect 13454 13613 13470 13677
rect 13534 13613 13550 13677
rect 13614 13613 13630 13677
rect 13694 13613 13710 13677
rect 13774 13613 13790 13677
rect 13854 13613 13870 13677
rect 13934 13613 13950 13677
rect 14014 13613 14030 13677
rect 14094 13613 14110 13677
rect 14174 13613 14190 13677
rect 14254 13613 14270 13677
rect 14334 13613 14350 13677
rect 14414 13613 14430 13677
rect 14494 13613 14510 13677
rect 14574 13613 14590 13677
rect 14654 13613 14670 13677
rect 14734 13613 14750 13677
rect 14814 13613 14830 13677
rect 14894 13613 14932 13677
rect 10152 13607 14932 13613
rect 120 13304 4900 13306
rect 120 13240 126 13304
rect 190 13240 207 13304
rect 271 13240 288 13304
rect 352 13240 369 13304
rect 433 13240 450 13304
rect 514 13240 531 13304
rect 595 13240 612 13304
rect 676 13240 693 13304
rect 757 13240 774 13304
rect 838 13240 855 13304
rect 919 13240 936 13304
rect 1000 13240 1017 13304
rect 1081 13240 1098 13304
rect 1162 13240 1179 13304
rect 1243 13240 1260 13304
rect 1324 13240 1341 13304
rect 1405 13240 1422 13304
rect 1486 13240 1503 13304
rect 1567 13240 1584 13304
rect 1648 13240 1665 13304
rect 1729 13240 1746 13304
rect 1810 13240 1827 13304
rect 1891 13240 1908 13304
rect 1972 13240 1989 13304
rect 2053 13240 2070 13304
rect 2134 13240 2151 13304
rect 2215 13240 2232 13304
rect 2296 13240 2313 13304
rect 2377 13240 2394 13304
rect 2458 13240 2475 13304
rect 2539 13240 2556 13304
rect 2620 13240 2637 13304
rect 2701 13240 2718 13304
rect 2782 13240 2799 13304
rect 2863 13240 2880 13304
rect 2944 13240 2961 13304
rect 3025 13240 3042 13304
rect 3106 13240 3123 13304
rect 3187 13240 3204 13304
rect 3268 13240 3285 13304
rect 3349 13240 3366 13304
rect 3430 13240 3447 13304
rect 3511 13240 3528 13304
rect 3592 13240 3609 13304
rect 3673 13240 3690 13304
rect 3754 13240 3771 13304
rect 3835 13240 3852 13304
rect 3916 13240 3933 13304
rect 3997 13240 4014 13304
rect 4078 13240 4095 13304
rect 4159 13240 4176 13304
rect 4240 13240 4257 13304
rect 4321 13240 4338 13304
rect 4402 13240 4420 13304
rect 4484 13240 4502 13304
rect 4566 13240 4584 13304
rect 4648 13240 4666 13304
rect 4730 13240 4748 13304
rect 4812 13240 4830 13304
rect 4894 13240 4900 13304
rect 120 13222 4900 13240
rect 120 13158 126 13222
rect 190 13158 207 13222
rect 271 13158 288 13222
rect 352 13158 369 13222
rect 433 13158 450 13222
rect 514 13158 531 13222
rect 595 13158 612 13222
rect 676 13158 693 13222
rect 757 13158 774 13222
rect 838 13158 855 13222
rect 919 13158 936 13222
rect 1000 13158 1017 13222
rect 1081 13158 1098 13222
rect 1162 13158 1179 13222
rect 1243 13158 1260 13222
rect 1324 13158 1341 13222
rect 1405 13158 1422 13222
rect 1486 13158 1503 13222
rect 1567 13158 1584 13222
rect 1648 13158 1665 13222
rect 1729 13158 1746 13222
rect 1810 13158 1827 13222
rect 1891 13158 1908 13222
rect 1972 13158 1989 13222
rect 2053 13158 2070 13222
rect 2134 13158 2151 13222
rect 2215 13158 2232 13222
rect 2296 13158 2313 13222
rect 2377 13158 2394 13222
rect 2458 13158 2475 13222
rect 2539 13158 2556 13222
rect 2620 13158 2637 13222
rect 2701 13158 2718 13222
rect 2782 13158 2799 13222
rect 2863 13158 2880 13222
rect 2944 13158 2961 13222
rect 3025 13158 3042 13222
rect 3106 13158 3123 13222
rect 3187 13158 3204 13222
rect 3268 13158 3285 13222
rect 3349 13158 3366 13222
rect 3430 13158 3447 13222
rect 3511 13158 3528 13222
rect 3592 13158 3609 13222
rect 3673 13158 3690 13222
rect 3754 13158 3771 13222
rect 3835 13158 3852 13222
rect 3916 13158 3933 13222
rect 3997 13158 4014 13222
rect 4078 13158 4095 13222
rect 4159 13158 4176 13222
rect 4240 13158 4257 13222
rect 4321 13158 4338 13222
rect 4402 13158 4420 13222
rect 4484 13158 4502 13222
rect 4566 13158 4584 13222
rect 4648 13158 4666 13222
rect 4730 13158 4748 13222
rect 4812 13158 4830 13222
rect 4894 13158 4900 13222
rect 120 13140 4900 13158
rect 120 13076 126 13140
rect 190 13076 207 13140
rect 271 13076 288 13140
rect 352 13076 369 13140
rect 433 13076 450 13140
rect 514 13076 531 13140
rect 595 13076 612 13140
rect 676 13076 693 13140
rect 757 13076 774 13140
rect 838 13076 855 13140
rect 919 13076 936 13140
rect 1000 13076 1017 13140
rect 1081 13076 1098 13140
rect 1162 13076 1179 13140
rect 1243 13076 1260 13140
rect 1324 13076 1341 13140
rect 1405 13076 1422 13140
rect 1486 13076 1503 13140
rect 1567 13076 1584 13140
rect 1648 13076 1665 13140
rect 1729 13076 1746 13140
rect 1810 13076 1827 13140
rect 1891 13076 1908 13140
rect 1972 13076 1989 13140
rect 2053 13076 2070 13140
rect 2134 13076 2151 13140
rect 2215 13076 2232 13140
rect 2296 13076 2313 13140
rect 2377 13076 2394 13140
rect 2458 13076 2475 13140
rect 2539 13076 2556 13140
rect 2620 13076 2637 13140
rect 2701 13076 2718 13140
rect 2782 13076 2799 13140
rect 2863 13076 2880 13140
rect 2944 13076 2961 13140
rect 3025 13076 3042 13140
rect 3106 13076 3123 13140
rect 3187 13076 3204 13140
rect 3268 13076 3285 13140
rect 3349 13076 3366 13140
rect 3430 13076 3447 13140
rect 3511 13076 3528 13140
rect 3592 13076 3609 13140
rect 3673 13076 3690 13140
rect 3754 13076 3771 13140
rect 3835 13076 3852 13140
rect 3916 13076 3933 13140
rect 3997 13076 4014 13140
rect 4078 13076 4095 13140
rect 4159 13076 4176 13140
rect 4240 13076 4257 13140
rect 4321 13076 4338 13140
rect 4402 13076 4420 13140
rect 4484 13076 4502 13140
rect 4566 13076 4584 13140
rect 4648 13076 4666 13140
rect 4730 13076 4748 13140
rect 4812 13076 4830 13140
rect 4894 13076 4900 13140
rect 120 13058 4900 13076
rect 120 12994 126 13058
rect 190 12994 207 13058
rect 271 12994 288 13058
rect 352 12994 369 13058
rect 433 12994 450 13058
rect 514 12994 531 13058
rect 595 12994 612 13058
rect 676 12994 693 13058
rect 757 12994 774 13058
rect 838 12994 855 13058
rect 919 12994 936 13058
rect 1000 12994 1017 13058
rect 1081 12994 1098 13058
rect 1162 12994 1179 13058
rect 1243 12994 1260 13058
rect 1324 12994 1341 13058
rect 1405 12994 1422 13058
rect 1486 12994 1503 13058
rect 1567 12994 1584 13058
rect 1648 12994 1665 13058
rect 1729 12994 1746 13058
rect 1810 12994 1827 13058
rect 1891 12994 1908 13058
rect 1972 12994 1989 13058
rect 2053 12994 2070 13058
rect 2134 12994 2151 13058
rect 2215 12994 2232 13058
rect 2296 12994 2313 13058
rect 2377 12994 2394 13058
rect 2458 12994 2475 13058
rect 2539 12994 2556 13058
rect 2620 12994 2637 13058
rect 2701 12994 2718 13058
rect 2782 12994 2799 13058
rect 2863 12994 2880 13058
rect 2944 12994 2961 13058
rect 3025 12994 3042 13058
rect 3106 12994 3123 13058
rect 3187 12994 3204 13058
rect 3268 12994 3285 13058
rect 3349 12994 3366 13058
rect 3430 12994 3447 13058
rect 3511 12994 3528 13058
rect 3592 12994 3609 13058
rect 3673 12994 3690 13058
rect 3754 12994 3771 13058
rect 3835 12994 3852 13058
rect 3916 12994 3933 13058
rect 3997 12994 4014 13058
rect 4078 12994 4095 13058
rect 4159 12994 4176 13058
rect 4240 12994 4257 13058
rect 4321 12994 4338 13058
rect 4402 12994 4420 13058
rect 4484 12994 4502 13058
rect 4566 12994 4584 13058
rect 4648 12994 4666 13058
rect 4730 12994 4748 13058
rect 4812 12994 4830 13058
rect 4894 12994 4900 13058
rect 120 12976 4900 12994
rect 120 12912 126 12976
rect 190 12912 207 12976
rect 271 12912 288 12976
rect 352 12912 369 12976
rect 433 12912 450 12976
rect 514 12912 531 12976
rect 595 12912 612 12976
rect 676 12912 693 12976
rect 757 12912 774 12976
rect 838 12912 855 12976
rect 919 12912 936 12976
rect 1000 12912 1017 12976
rect 1081 12912 1098 12976
rect 1162 12912 1179 12976
rect 1243 12912 1260 12976
rect 1324 12912 1341 12976
rect 1405 12912 1422 12976
rect 1486 12912 1503 12976
rect 1567 12912 1584 12976
rect 1648 12912 1665 12976
rect 1729 12912 1746 12976
rect 1810 12912 1827 12976
rect 1891 12912 1908 12976
rect 1972 12912 1989 12976
rect 2053 12912 2070 12976
rect 2134 12912 2151 12976
rect 2215 12912 2232 12976
rect 2296 12912 2313 12976
rect 2377 12912 2394 12976
rect 2458 12912 2475 12976
rect 2539 12912 2556 12976
rect 2620 12912 2637 12976
rect 2701 12912 2718 12976
rect 2782 12912 2799 12976
rect 2863 12912 2880 12976
rect 2944 12912 2961 12976
rect 3025 12912 3042 12976
rect 3106 12912 3123 12976
rect 3187 12912 3204 12976
rect 3268 12912 3285 12976
rect 3349 12912 3366 12976
rect 3430 12912 3447 12976
rect 3511 12912 3528 12976
rect 3592 12912 3609 12976
rect 3673 12912 3690 12976
rect 3754 12912 3771 12976
rect 3835 12912 3852 12976
rect 3916 12912 3933 12976
rect 3997 12912 4014 12976
rect 4078 12912 4095 12976
rect 4159 12912 4176 12976
rect 4240 12912 4257 12976
rect 4321 12912 4338 12976
rect 4402 12912 4420 12976
rect 4484 12912 4502 12976
rect 4566 12912 4584 12976
rect 4648 12912 4666 12976
rect 4730 12912 4748 12976
rect 4812 12912 4830 12976
rect 4894 12912 4900 12976
rect 120 12894 4900 12912
rect 120 12830 126 12894
rect 190 12830 207 12894
rect 271 12830 288 12894
rect 352 12830 369 12894
rect 433 12830 450 12894
rect 514 12830 531 12894
rect 595 12830 612 12894
rect 676 12830 693 12894
rect 757 12830 774 12894
rect 838 12830 855 12894
rect 919 12830 936 12894
rect 1000 12830 1017 12894
rect 1081 12830 1098 12894
rect 1162 12830 1179 12894
rect 1243 12830 1260 12894
rect 1324 12830 1341 12894
rect 1405 12830 1422 12894
rect 1486 12830 1503 12894
rect 1567 12830 1584 12894
rect 1648 12830 1665 12894
rect 1729 12830 1746 12894
rect 1810 12830 1827 12894
rect 1891 12830 1908 12894
rect 1972 12830 1989 12894
rect 2053 12830 2070 12894
rect 2134 12830 2151 12894
rect 2215 12830 2232 12894
rect 2296 12830 2313 12894
rect 2377 12830 2394 12894
rect 2458 12830 2475 12894
rect 2539 12830 2556 12894
rect 2620 12830 2637 12894
rect 2701 12830 2718 12894
rect 2782 12830 2799 12894
rect 2863 12830 2880 12894
rect 2944 12830 2961 12894
rect 3025 12830 3042 12894
rect 3106 12830 3123 12894
rect 3187 12830 3204 12894
rect 3268 12830 3285 12894
rect 3349 12830 3366 12894
rect 3430 12830 3447 12894
rect 3511 12830 3528 12894
rect 3592 12830 3609 12894
rect 3673 12830 3690 12894
rect 3754 12830 3771 12894
rect 3835 12830 3852 12894
rect 3916 12830 3933 12894
rect 3997 12830 4014 12894
rect 4078 12830 4095 12894
rect 4159 12830 4176 12894
rect 4240 12830 4257 12894
rect 4321 12830 4338 12894
rect 4402 12830 4420 12894
rect 4484 12830 4502 12894
rect 4566 12830 4584 12894
rect 4648 12830 4666 12894
rect 4730 12830 4748 12894
rect 4812 12830 4830 12894
rect 4894 12830 4900 12894
rect 120 12812 4900 12830
rect 120 12748 126 12812
rect 190 12748 207 12812
rect 271 12748 288 12812
rect 352 12748 369 12812
rect 433 12748 450 12812
rect 514 12748 531 12812
rect 595 12748 612 12812
rect 676 12748 693 12812
rect 757 12748 774 12812
rect 838 12748 855 12812
rect 919 12748 936 12812
rect 1000 12748 1017 12812
rect 1081 12748 1098 12812
rect 1162 12748 1179 12812
rect 1243 12748 1260 12812
rect 1324 12748 1341 12812
rect 1405 12748 1422 12812
rect 1486 12748 1503 12812
rect 1567 12748 1584 12812
rect 1648 12748 1665 12812
rect 1729 12748 1746 12812
rect 1810 12748 1827 12812
rect 1891 12748 1908 12812
rect 1972 12748 1989 12812
rect 2053 12748 2070 12812
rect 2134 12748 2151 12812
rect 2215 12748 2232 12812
rect 2296 12748 2313 12812
rect 2377 12748 2394 12812
rect 2458 12748 2475 12812
rect 2539 12748 2556 12812
rect 2620 12748 2637 12812
rect 2701 12748 2718 12812
rect 2782 12748 2799 12812
rect 2863 12748 2880 12812
rect 2944 12748 2961 12812
rect 3025 12748 3042 12812
rect 3106 12748 3123 12812
rect 3187 12748 3204 12812
rect 3268 12748 3285 12812
rect 3349 12748 3366 12812
rect 3430 12748 3447 12812
rect 3511 12748 3528 12812
rect 3592 12748 3609 12812
rect 3673 12748 3690 12812
rect 3754 12748 3771 12812
rect 3835 12748 3852 12812
rect 3916 12748 3933 12812
rect 3997 12748 4014 12812
rect 4078 12748 4095 12812
rect 4159 12748 4176 12812
rect 4240 12748 4257 12812
rect 4321 12748 4338 12812
rect 4402 12748 4420 12812
rect 4484 12748 4502 12812
rect 4566 12748 4584 12812
rect 4648 12748 4666 12812
rect 4730 12748 4748 12812
rect 4812 12748 4830 12812
rect 4894 12748 4900 12812
rect 120 12730 4900 12748
rect 120 12666 126 12730
rect 190 12666 207 12730
rect 271 12666 288 12730
rect 352 12666 369 12730
rect 433 12666 450 12730
rect 514 12666 531 12730
rect 595 12666 612 12730
rect 676 12666 693 12730
rect 757 12666 774 12730
rect 838 12666 855 12730
rect 919 12666 936 12730
rect 1000 12666 1017 12730
rect 1081 12666 1098 12730
rect 1162 12666 1179 12730
rect 1243 12666 1260 12730
rect 1324 12666 1341 12730
rect 1405 12666 1422 12730
rect 1486 12666 1503 12730
rect 1567 12666 1584 12730
rect 1648 12666 1665 12730
rect 1729 12666 1746 12730
rect 1810 12666 1827 12730
rect 1891 12666 1908 12730
rect 1972 12666 1989 12730
rect 2053 12666 2070 12730
rect 2134 12666 2151 12730
rect 2215 12666 2232 12730
rect 2296 12666 2313 12730
rect 2377 12666 2394 12730
rect 2458 12666 2475 12730
rect 2539 12666 2556 12730
rect 2620 12666 2637 12730
rect 2701 12666 2718 12730
rect 2782 12666 2799 12730
rect 2863 12666 2880 12730
rect 2944 12666 2961 12730
rect 3025 12666 3042 12730
rect 3106 12666 3123 12730
rect 3187 12666 3204 12730
rect 3268 12666 3285 12730
rect 3349 12666 3366 12730
rect 3430 12666 3447 12730
rect 3511 12666 3528 12730
rect 3592 12666 3609 12730
rect 3673 12666 3690 12730
rect 3754 12666 3771 12730
rect 3835 12666 3852 12730
rect 3916 12666 3933 12730
rect 3997 12666 4014 12730
rect 4078 12666 4095 12730
rect 4159 12666 4176 12730
rect 4240 12666 4257 12730
rect 4321 12666 4338 12730
rect 4402 12666 4420 12730
rect 4484 12666 4502 12730
rect 4566 12666 4584 12730
rect 4648 12666 4666 12730
rect 4730 12666 4748 12730
rect 4812 12666 4830 12730
rect 4894 12666 4900 12730
rect 120 12648 4900 12666
rect 120 12584 126 12648
rect 190 12584 207 12648
rect 271 12584 288 12648
rect 352 12584 369 12648
rect 433 12584 450 12648
rect 514 12584 531 12648
rect 595 12584 612 12648
rect 676 12584 693 12648
rect 757 12584 774 12648
rect 838 12584 855 12648
rect 919 12584 936 12648
rect 1000 12584 1017 12648
rect 1081 12584 1098 12648
rect 1162 12584 1179 12648
rect 1243 12584 1260 12648
rect 1324 12584 1341 12648
rect 1405 12584 1422 12648
rect 1486 12584 1503 12648
rect 1567 12584 1584 12648
rect 1648 12584 1665 12648
rect 1729 12584 1746 12648
rect 1810 12584 1827 12648
rect 1891 12584 1908 12648
rect 1972 12584 1989 12648
rect 2053 12584 2070 12648
rect 2134 12584 2151 12648
rect 2215 12584 2232 12648
rect 2296 12584 2313 12648
rect 2377 12584 2394 12648
rect 2458 12584 2475 12648
rect 2539 12584 2556 12648
rect 2620 12584 2637 12648
rect 2701 12584 2718 12648
rect 2782 12584 2799 12648
rect 2863 12584 2880 12648
rect 2944 12584 2961 12648
rect 3025 12584 3042 12648
rect 3106 12584 3123 12648
rect 3187 12584 3204 12648
rect 3268 12584 3285 12648
rect 3349 12584 3366 12648
rect 3430 12584 3447 12648
rect 3511 12584 3528 12648
rect 3592 12584 3609 12648
rect 3673 12584 3690 12648
rect 3754 12584 3771 12648
rect 3835 12584 3852 12648
rect 3916 12584 3933 12648
rect 3997 12584 4014 12648
rect 4078 12584 4095 12648
rect 4159 12584 4176 12648
rect 4240 12584 4257 12648
rect 4321 12584 4338 12648
rect 4402 12584 4420 12648
rect 4484 12584 4502 12648
rect 4566 12584 4584 12648
rect 4648 12584 4666 12648
rect 4730 12584 4748 12648
rect 4812 12584 4830 12648
rect 4894 12584 4900 12648
rect 120 12566 4900 12584
rect 120 12502 126 12566
rect 190 12502 207 12566
rect 271 12502 288 12566
rect 352 12502 369 12566
rect 433 12502 450 12566
rect 514 12502 531 12566
rect 595 12502 612 12566
rect 676 12502 693 12566
rect 757 12502 774 12566
rect 838 12502 855 12566
rect 919 12502 936 12566
rect 1000 12502 1017 12566
rect 1081 12502 1098 12566
rect 1162 12502 1179 12566
rect 1243 12502 1260 12566
rect 1324 12502 1341 12566
rect 1405 12502 1422 12566
rect 1486 12502 1503 12566
rect 1567 12502 1584 12566
rect 1648 12502 1665 12566
rect 1729 12502 1746 12566
rect 1810 12502 1827 12566
rect 1891 12502 1908 12566
rect 1972 12502 1989 12566
rect 2053 12502 2070 12566
rect 2134 12502 2151 12566
rect 2215 12502 2232 12566
rect 2296 12502 2313 12566
rect 2377 12502 2394 12566
rect 2458 12502 2475 12566
rect 2539 12502 2556 12566
rect 2620 12502 2637 12566
rect 2701 12502 2718 12566
rect 2782 12502 2799 12566
rect 2863 12502 2880 12566
rect 2944 12502 2961 12566
rect 3025 12502 3042 12566
rect 3106 12502 3123 12566
rect 3187 12502 3204 12566
rect 3268 12502 3285 12566
rect 3349 12502 3366 12566
rect 3430 12502 3447 12566
rect 3511 12502 3528 12566
rect 3592 12502 3609 12566
rect 3673 12502 3690 12566
rect 3754 12502 3771 12566
rect 3835 12502 3852 12566
rect 3916 12502 3933 12566
rect 3997 12502 4014 12566
rect 4078 12502 4095 12566
rect 4159 12502 4176 12566
rect 4240 12502 4257 12566
rect 4321 12502 4338 12566
rect 4402 12502 4420 12566
rect 4484 12502 4502 12566
rect 4566 12502 4584 12566
rect 4648 12502 4666 12566
rect 4730 12502 4748 12566
rect 4812 12502 4830 12566
rect 4894 12502 4900 12566
rect 120 12484 4900 12502
rect 120 12420 126 12484
rect 190 12420 207 12484
rect 271 12420 288 12484
rect 352 12420 369 12484
rect 433 12420 450 12484
rect 514 12420 531 12484
rect 595 12420 612 12484
rect 676 12420 693 12484
rect 757 12420 774 12484
rect 838 12420 855 12484
rect 919 12420 936 12484
rect 1000 12420 1017 12484
rect 1081 12420 1098 12484
rect 1162 12420 1179 12484
rect 1243 12420 1260 12484
rect 1324 12420 1341 12484
rect 1405 12420 1422 12484
rect 1486 12420 1503 12484
rect 1567 12420 1584 12484
rect 1648 12420 1665 12484
rect 1729 12420 1746 12484
rect 1810 12420 1827 12484
rect 1891 12420 1908 12484
rect 1972 12420 1989 12484
rect 2053 12420 2070 12484
rect 2134 12420 2151 12484
rect 2215 12420 2232 12484
rect 2296 12420 2313 12484
rect 2377 12420 2394 12484
rect 2458 12420 2475 12484
rect 2539 12420 2556 12484
rect 2620 12420 2637 12484
rect 2701 12420 2718 12484
rect 2782 12420 2799 12484
rect 2863 12420 2880 12484
rect 2944 12420 2961 12484
rect 3025 12420 3042 12484
rect 3106 12420 3123 12484
rect 3187 12420 3204 12484
rect 3268 12420 3285 12484
rect 3349 12420 3366 12484
rect 3430 12420 3447 12484
rect 3511 12420 3528 12484
rect 3592 12420 3609 12484
rect 3673 12420 3690 12484
rect 3754 12420 3771 12484
rect 3835 12420 3852 12484
rect 3916 12420 3933 12484
rect 3997 12420 4014 12484
rect 4078 12420 4095 12484
rect 4159 12420 4176 12484
rect 4240 12420 4257 12484
rect 4321 12420 4338 12484
rect 4402 12420 4420 12484
rect 4484 12420 4502 12484
rect 4566 12420 4584 12484
rect 4648 12420 4666 12484
rect 4730 12420 4748 12484
rect 4812 12420 4830 12484
rect 4894 12420 4900 12484
rect 120 12418 4900 12420
rect 10151 13304 14931 13306
rect 10151 13240 10157 13304
rect 10221 13240 10238 13304
rect 10302 13240 10319 13304
rect 10383 13240 10400 13304
rect 10464 13240 10481 13304
rect 10545 13240 10562 13304
rect 10626 13240 10643 13304
rect 10707 13240 10724 13304
rect 10788 13240 10805 13304
rect 10869 13240 10886 13304
rect 10950 13240 10967 13304
rect 11031 13240 11048 13304
rect 11112 13240 11129 13304
rect 11193 13240 11210 13304
rect 11274 13240 11291 13304
rect 11355 13240 11372 13304
rect 11436 13240 11453 13304
rect 11517 13240 11534 13304
rect 11598 13240 11615 13304
rect 11679 13240 11696 13304
rect 11760 13240 11777 13304
rect 11841 13240 11858 13304
rect 11922 13240 11939 13304
rect 12003 13240 12020 13304
rect 12084 13240 12101 13304
rect 12165 13240 12182 13304
rect 12246 13240 12263 13304
rect 12327 13240 12344 13304
rect 12408 13240 12425 13304
rect 12489 13240 12506 13304
rect 12570 13240 12587 13304
rect 12651 13240 12668 13304
rect 12732 13240 12749 13304
rect 12813 13240 12830 13304
rect 12894 13240 12911 13304
rect 12975 13240 12992 13304
rect 13056 13240 13073 13304
rect 13137 13240 13154 13304
rect 13218 13240 13235 13304
rect 13299 13240 13316 13304
rect 13380 13240 13397 13304
rect 13461 13240 13478 13304
rect 13542 13240 13559 13304
rect 13623 13240 13640 13304
rect 13704 13240 13721 13304
rect 13785 13240 13802 13304
rect 13866 13240 13883 13304
rect 13947 13240 13964 13304
rect 14028 13240 14045 13304
rect 14109 13240 14126 13304
rect 14190 13240 14207 13304
rect 14271 13240 14288 13304
rect 14352 13240 14369 13304
rect 14433 13240 14451 13304
rect 14515 13240 14533 13304
rect 14597 13240 14615 13304
rect 14679 13240 14697 13304
rect 14761 13240 14779 13304
rect 14843 13240 14861 13304
rect 14925 13240 14931 13304
rect 10151 13222 14931 13240
rect 10151 13158 10157 13222
rect 10221 13158 10238 13222
rect 10302 13158 10319 13222
rect 10383 13158 10400 13222
rect 10464 13158 10481 13222
rect 10545 13158 10562 13222
rect 10626 13158 10643 13222
rect 10707 13158 10724 13222
rect 10788 13158 10805 13222
rect 10869 13158 10886 13222
rect 10950 13158 10967 13222
rect 11031 13158 11048 13222
rect 11112 13158 11129 13222
rect 11193 13158 11210 13222
rect 11274 13158 11291 13222
rect 11355 13158 11372 13222
rect 11436 13158 11453 13222
rect 11517 13158 11534 13222
rect 11598 13158 11615 13222
rect 11679 13158 11696 13222
rect 11760 13158 11777 13222
rect 11841 13158 11858 13222
rect 11922 13158 11939 13222
rect 12003 13158 12020 13222
rect 12084 13158 12101 13222
rect 12165 13158 12182 13222
rect 12246 13158 12263 13222
rect 12327 13158 12344 13222
rect 12408 13158 12425 13222
rect 12489 13158 12506 13222
rect 12570 13158 12587 13222
rect 12651 13158 12668 13222
rect 12732 13158 12749 13222
rect 12813 13158 12830 13222
rect 12894 13158 12911 13222
rect 12975 13158 12992 13222
rect 13056 13158 13073 13222
rect 13137 13158 13154 13222
rect 13218 13158 13235 13222
rect 13299 13158 13316 13222
rect 13380 13158 13397 13222
rect 13461 13158 13478 13222
rect 13542 13158 13559 13222
rect 13623 13158 13640 13222
rect 13704 13158 13721 13222
rect 13785 13158 13802 13222
rect 13866 13158 13883 13222
rect 13947 13158 13964 13222
rect 14028 13158 14045 13222
rect 14109 13158 14126 13222
rect 14190 13158 14207 13222
rect 14271 13158 14288 13222
rect 14352 13158 14369 13222
rect 14433 13158 14451 13222
rect 14515 13158 14533 13222
rect 14597 13158 14615 13222
rect 14679 13158 14697 13222
rect 14761 13158 14779 13222
rect 14843 13158 14861 13222
rect 14925 13158 14931 13222
rect 10151 13140 14931 13158
rect 10151 13076 10157 13140
rect 10221 13076 10238 13140
rect 10302 13076 10319 13140
rect 10383 13076 10400 13140
rect 10464 13076 10481 13140
rect 10545 13076 10562 13140
rect 10626 13076 10643 13140
rect 10707 13076 10724 13140
rect 10788 13076 10805 13140
rect 10869 13076 10886 13140
rect 10950 13076 10967 13140
rect 11031 13076 11048 13140
rect 11112 13076 11129 13140
rect 11193 13076 11210 13140
rect 11274 13076 11291 13140
rect 11355 13076 11372 13140
rect 11436 13076 11453 13140
rect 11517 13076 11534 13140
rect 11598 13076 11615 13140
rect 11679 13076 11696 13140
rect 11760 13076 11777 13140
rect 11841 13076 11858 13140
rect 11922 13076 11939 13140
rect 12003 13076 12020 13140
rect 12084 13076 12101 13140
rect 12165 13076 12182 13140
rect 12246 13076 12263 13140
rect 12327 13076 12344 13140
rect 12408 13076 12425 13140
rect 12489 13076 12506 13140
rect 12570 13076 12587 13140
rect 12651 13076 12668 13140
rect 12732 13076 12749 13140
rect 12813 13076 12830 13140
rect 12894 13076 12911 13140
rect 12975 13076 12992 13140
rect 13056 13076 13073 13140
rect 13137 13076 13154 13140
rect 13218 13076 13235 13140
rect 13299 13076 13316 13140
rect 13380 13076 13397 13140
rect 13461 13076 13478 13140
rect 13542 13076 13559 13140
rect 13623 13076 13640 13140
rect 13704 13076 13721 13140
rect 13785 13076 13802 13140
rect 13866 13076 13883 13140
rect 13947 13076 13964 13140
rect 14028 13076 14045 13140
rect 14109 13076 14126 13140
rect 14190 13076 14207 13140
rect 14271 13076 14288 13140
rect 14352 13076 14369 13140
rect 14433 13076 14451 13140
rect 14515 13076 14533 13140
rect 14597 13076 14615 13140
rect 14679 13076 14697 13140
rect 14761 13076 14779 13140
rect 14843 13076 14861 13140
rect 14925 13076 14931 13140
rect 10151 13058 14931 13076
rect 10151 12994 10157 13058
rect 10221 12994 10238 13058
rect 10302 12994 10319 13058
rect 10383 12994 10400 13058
rect 10464 12994 10481 13058
rect 10545 12994 10562 13058
rect 10626 12994 10643 13058
rect 10707 12994 10724 13058
rect 10788 12994 10805 13058
rect 10869 12994 10886 13058
rect 10950 12994 10967 13058
rect 11031 12994 11048 13058
rect 11112 12994 11129 13058
rect 11193 12994 11210 13058
rect 11274 12994 11291 13058
rect 11355 12994 11372 13058
rect 11436 12994 11453 13058
rect 11517 12994 11534 13058
rect 11598 12994 11615 13058
rect 11679 12994 11696 13058
rect 11760 12994 11777 13058
rect 11841 12994 11858 13058
rect 11922 12994 11939 13058
rect 12003 12994 12020 13058
rect 12084 12994 12101 13058
rect 12165 12994 12182 13058
rect 12246 12994 12263 13058
rect 12327 12994 12344 13058
rect 12408 12994 12425 13058
rect 12489 12994 12506 13058
rect 12570 12994 12587 13058
rect 12651 12994 12668 13058
rect 12732 12994 12749 13058
rect 12813 12994 12830 13058
rect 12894 12994 12911 13058
rect 12975 12994 12992 13058
rect 13056 12994 13073 13058
rect 13137 12994 13154 13058
rect 13218 12994 13235 13058
rect 13299 12994 13316 13058
rect 13380 12994 13397 13058
rect 13461 12994 13478 13058
rect 13542 12994 13559 13058
rect 13623 12994 13640 13058
rect 13704 12994 13721 13058
rect 13785 12994 13802 13058
rect 13866 12994 13883 13058
rect 13947 12994 13964 13058
rect 14028 12994 14045 13058
rect 14109 12994 14126 13058
rect 14190 12994 14207 13058
rect 14271 12994 14288 13058
rect 14352 12994 14369 13058
rect 14433 12994 14451 13058
rect 14515 12994 14533 13058
rect 14597 12994 14615 13058
rect 14679 12994 14697 13058
rect 14761 12994 14779 13058
rect 14843 12994 14861 13058
rect 14925 12994 14931 13058
rect 10151 12976 14931 12994
rect 10151 12912 10157 12976
rect 10221 12912 10238 12976
rect 10302 12912 10319 12976
rect 10383 12912 10400 12976
rect 10464 12912 10481 12976
rect 10545 12912 10562 12976
rect 10626 12912 10643 12976
rect 10707 12912 10724 12976
rect 10788 12912 10805 12976
rect 10869 12912 10886 12976
rect 10950 12912 10967 12976
rect 11031 12912 11048 12976
rect 11112 12912 11129 12976
rect 11193 12912 11210 12976
rect 11274 12912 11291 12976
rect 11355 12912 11372 12976
rect 11436 12912 11453 12976
rect 11517 12912 11534 12976
rect 11598 12912 11615 12976
rect 11679 12912 11696 12976
rect 11760 12912 11777 12976
rect 11841 12912 11858 12976
rect 11922 12912 11939 12976
rect 12003 12912 12020 12976
rect 12084 12912 12101 12976
rect 12165 12912 12182 12976
rect 12246 12912 12263 12976
rect 12327 12912 12344 12976
rect 12408 12912 12425 12976
rect 12489 12912 12506 12976
rect 12570 12912 12587 12976
rect 12651 12912 12668 12976
rect 12732 12912 12749 12976
rect 12813 12912 12830 12976
rect 12894 12912 12911 12976
rect 12975 12912 12992 12976
rect 13056 12912 13073 12976
rect 13137 12912 13154 12976
rect 13218 12912 13235 12976
rect 13299 12912 13316 12976
rect 13380 12912 13397 12976
rect 13461 12912 13478 12976
rect 13542 12912 13559 12976
rect 13623 12912 13640 12976
rect 13704 12912 13721 12976
rect 13785 12912 13802 12976
rect 13866 12912 13883 12976
rect 13947 12912 13964 12976
rect 14028 12912 14045 12976
rect 14109 12912 14126 12976
rect 14190 12912 14207 12976
rect 14271 12912 14288 12976
rect 14352 12912 14369 12976
rect 14433 12912 14451 12976
rect 14515 12912 14533 12976
rect 14597 12912 14615 12976
rect 14679 12912 14697 12976
rect 14761 12912 14779 12976
rect 14843 12912 14861 12976
rect 14925 12912 14931 12976
rect 10151 12894 14931 12912
rect 10151 12830 10157 12894
rect 10221 12830 10238 12894
rect 10302 12830 10319 12894
rect 10383 12830 10400 12894
rect 10464 12830 10481 12894
rect 10545 12830 10562 12894
rect 10626 12830 10643 12894
rect 10707 12830 10724 12894
rect 10788 12830 10805 12894
rect 10869 12830 10886 12894
rect 10950 12830 10967 12894
rect 11031 12830 11048 12894
rect 11112 12830 11129 12894
rect 11193 12830 11210 12894
rect 11274 12830 11291 12894
rect 11355 12830 11372 12894
rect 11436 12830 11453 12894
rect 11517 12830 11534 12894
rect 11598 12830 11615 12894
rect 11679 12830 11696 12894
rect 11760 12830 11777 12894
rect 11841 12830 11858 12894
rect 11922 12830 11939 12894
rect 12003 12830 12020 12894
rect 12084 12830 12101 12894
rect 12165 12830 12182 12894
rect 12246 12830 12263 12894
rect 12327 12830 12344 12894
rect 12408 12830 12425 12894
rect 12489 12830 12506 12894
rect 12570 12830 12587 12894
rect 12651 12830 12668 12894
rect 12732 12830 12749 12894
rect 12813 12830 12830 12894
rect 12894 12830 12911 12894
rect 12975 12830 12992 12894
rect 13056 12830 13073 12894
rect 13137 12830 13154 12894
rect 13218 12830 13235 12894
rect 13299 12830 13316 12894
rect 13380 12830 13397 12894
rect 13461 12830 13478 12894
rect 13542 12830 13559 12894
rect 13623 12830 13640 12894
rect 13704 12830 13721 12894
rect 13785 12830 13802 12894
rect 13866 12830 13883 12894
rect 13947 12830 13964 12894
rect 14028 12830 14045 12894
rect 14109 12830 14126 12894
rect 14190 12830 14207 12894
rect 14271 12830 14288 12894
rect 14352 12830 14369 12894
rect 14433 12830 14451 12894
rect 14515 12830 14533 12894
rect 14597 12830 14615 12894
rect 14679 12830 14697 12894
rect 14761 12830 14779 12894
rect 14843 12830 14861 12894
rect 14925 12830 14931 12894
rect 10151 12812 14931 12830
rect 10151 12748 10157 12812
rect 10221 12748 10238 12812
rect 10302 12748 10319 12812
rect 10383 12748 10400 12812
rect 10464 12748 10481 12812
rect 10545 12748 10562 12812
rect 10626 12748 10643 12812
rect 10707 12748 10724 12812
rect 10788 12748 10805 12812
rect 10869 12748 10886 12812
rect 10950 12748 10967 12812
rect 11031 12748 11048 12812
rect 11112 12748 11129 12812
rect 11193 12748 11210 12812
rect 11274 12748 11291 12812
rect 11355 12748 11372 12812
rect 11436 12748 11453 12812
rect 11517 12748 11534 12812
rect 11598 12748 11615 12812
rect 11679 12748 11696 12812
rect 11760 12748 11777 12812
rect 11841 12748 11858 12812
rect 11922 12748 11939 12812
rect 12003 12748 12020 12812
rect 12084 12748 12101 12812
rect 12165 12748 12182 12812
rect 12246 12748 12263 12812
rect 12327 12748 12344 12812
rect 12408 12748 12425 12812
rect 12489 12748 12506 12812
rect 12570 12748 12587 12812
rect 12651 12748 12668 12812
rect 12732 12748 12749 12812
rect 12813 12748 12830 12812
rect 12894 12748 12911 12812
rect 12975 12748 12992 12812
rect 13056 12748 13073 12812
rect 13137 12748 13154 12812
rect 13218 12748 13235 12812
rect 13299 12748 13316 12812
rect 13380 12748 13397 12812
rect 13461 12748 13478 12812
rect 13542 12748 13559 12812
rect 13623 12748 13640 12812
rect 13704 12748 13721 12812
rect 13785 12748 13802 12812
rect 13866 12748 13883 12812
rect 13947 12748 13964 12812
rect 14028 12748 14045 12812
rect 14109 12748 14126 12812
rect 14190 12748 14207 12812
rect 14271 12748 14288 12812
rect 14352 12748 14369 12812
rect 14433 12748 14451 12812
rect 14515 12748 14533 12812
rect 14597 12748 14615 12812
rect 14679 12748 14697 12812
rect 14761 12748 14779 12812
rect 14843 12748 14861 12812
rect 14925 12748 14931 12812
rect 10151 12730 14931 12748
rect 10151 12666 10157 12730
rect 10221 12666 10238 12730
rect 10302 12666 10319 12730
rect 10383 12666 10400 12730
rect 10464 12666 10481 12730
rect 10545 12666 10562 12730
rect 10626 12666 10643 12730
rect 10707 12666 10724 12730
rect 10788 12666 10805 12730
rect 10869 12666 10886 12730
rect 10950 12666 10967 12730
rect 11031 12666 11048 12730
rect 11112 12666 11129 12730
rect 11193 12666 11210 12730
rect 11274 12666 11291 12730
rect 11355 12666 11372 12730
rect 11436 12666 11453 12730
rect 11517 12666 11534 12730
rect 11598 12666 11615 12730
rect 11679 12666 11696 12730
rect 11760 12666 11777 12730
rect 11841 12666 11858 12730
rect 11922 12666 11939 12730
rect 12003 12666 12020 12730
rect 12084 12666 12101 12730
rect 12165 12666 12182 12730
rect 12246 12666 12263 12730
rect 12327 12666 12344 12730
rect 12408 12666 12425 12730
rect 12489 12666 12506 12730
rect 12570 12666 12587 12730
rect 12651 12666 12668 12730
rect 12732 12666 12749 12730
rect 12813 12666 12830 12730
rect 12894 12666 12911 12730
rect 12975 12666 12992 12730
rect 13056 12666 13073 12730
rect 13137 12666 13154 12730
rect 13218 12666 13235 12730
rect 13299 12666 13316 12730
rect 13380 12666 13397 12730
rect 13461 12666 13478 12730
rect 13542 12666 13559 12730
rect 13623 12666 13640 12730
rect 13704 12666 13721 12730
rect 13785 12666 13802 12730
rect 13866 12666 13883 12730
rect 13947 12666 13964 12730
rect 14028 12666 14045 12730
rect 14109 12666 14126 12730
rect 14190 12666 14207 12730
rect 14271 12666 14288 12730
rect 14352 12666 14369 12730
rect 14433 12666 14451 12730
rect 14515 12666 14533 12730
rect 14597 12666 14615 12730
rect 14679 12666 14697 12730
rect 14761 12666 14779 12730
rect 14843 12666 14861 12730
rect 14925 12666 14931 12730
rect 10151 12648 14931 12666
rect 10151 12584 10157 12648
rect 10221 12584 10238 12648
rect 10302 12584 10319 12648
rect 10383 12584 10400 12648
rect 10464 12584 10481 12648
rect 10545 12584 10562 12648
rect 10626 12584 10643 12648
rect 10707 12584 10724 12648
rect 10788 12584 10805 12648
rect 10869 12584 10886 12648
rect 10950 12584 10967 12648
rect 11031 12584 11048 12648
rect 11112 12584 11129 12648
rect 11193 12584 11210 12648
rect 11274 12584 11291 12648
rect 11355 12584 11372 12648
rect 11436 12584 11453 12648
rect 11517 12584 11534 12648
rect 11598 12584 11615 12648
rect 11679 12584 11696 12648
rect 11760 12584 11777 12648
rect 11841 12584 11858 12648
rect 11922 12584 11939 12648
rect 12003 12584 12020 12648
rect 12084 12584 12101 12648
rect 12165 12584 12182 12648
rect 12246 12584 12263 12648
rect 12327 12584 12344 12648
rect 12408 12584 12425 12648
rect 12489 12584 12506 12648
rect 12570 12584 12587 12648
rect 12651 12584 12668 12648
rect 12732 12584 12749 12648
rect 12813 12584 12830 12648
rect 12894 12584 12911 12648
rect 12975 12584 12992 12648
rect 13056 12584 13073 12648
rect 13137 12584 13154 12648
rect 13218 12584 13235 12648
rect 13299 12584 13316 12648
rect 13380 12584 13397 12648
rect 13461 12584 13478 12648
rect 13542 12584 13559 12648
rect 13623 12584 13640 12648
rect 13704 12584 13721 12648
rect 13785 12584 13802 12648
rect 13866 12584 13883 12648
rect 13947 12584 13964 12648
rect 14028 12584 14045 12648
rect 14109 12584 14126 12648
rect 14190 12584 14207 12648
rect 14271 12584 14288 12648
rect 14352 12584 14369 12648
rect 14433 12584 14451 12648
rect 14515 12584 14533 12648
rect 14597 12584 14615 12648
rect 14679 12584 14697 12648
rect 14761 12584 14779 12648
rect 14843 12584 14861 12648
rect 14925 12584 14931 12648
rect 10151 12566 14931 12584
rect 10151 12502 10157 12566
rect 10221 12502 10238 12566
rect 10302 12502 10319 12566
rect 10383 12502 10400 12566
rect 10464 12502 10481 12566
rect 10545 12502 10562 12566
rect 10626 12502 10643 12566
rect 10707 12502 10724 12566
rect 10788 12502 10805 12566
rect 10869 12502 10886 12566
rect 10950 12502 10967 12566
rect 11031 12502 11048 12566
rect 11112 12502 11129 12566
rect 11193 12502 11210 12566
rect 11274 12502 11291 12566
rect 11355 12502 11372 12566
rect 11436 12502 11453 12566
rect 11517 12502 11534 12566
rect 11598 12502 11615 12566
rect 11679 12502 11696 12566
rect 11760 12502 11777 12566
rect 11841 12502 11858 12566
rect 11922 12502 11939 12566
rect 12003 12502 12020 12566
rect 12084 12502 12101 12566
rect 12165 12502 12182 12566
rect 12246 12502 12263 12566
rect 12327 12502 12344 12566
rect 12408 12502 12425 12566
rect 12489 12502 12506 12566
rect 12570 12502 12587 12566
rect 12651 12502 12668 12566
rect 12732 12502 12749 12566
rect 12813 12502 12830 12566
rect 12894 12502 12911 12566
rect 12975 12502 12992 12566
rect 13056 12502 13073 12566
rect 13137 12502 13154 12566
rect 13218 12502 13235 12566
rect 13299 12502 13316 12566
rect 13380 12502 13397 12566
rect 13461 12502 13478 12566
rect 13542 12502 13559 12566
rect 13623 12502 13640 12566
rect 13704 12502 13721 12566
rect 13785 12502 13802 12566
rect 13866 12502 13883 12566
rect 13947 12502 13964 12566
rect 14028 12502 14045 12566
rect 14109 12502 14126 12566
rect 14190 12502 14207 12566
rect 14271 12502 14288 12566
rect 14352 12502 14369 12566
rect 14433 12502 14451 12566
rect 14515 12502 14533 12566
rect 14597 12502 14615 12566
rect 14679 12502 14697 12566
rect 14761 12502 14779 12566
rect 14843 12502 14861 12566
rect 14925 12502 14931 12566
rect 10151 12484 14931 12502
rect 10151 12420 10157 12484
rect 10221 12420 10238 12484
rect 10302 12420 10319 12484
rect 10383 12420 10400 12484
rect 10464 12420 10481 12484
rect 10545 12420 10562 12484
rect 10626 12420 10643 12484
rect 10707 12420 10724 12484
rect 10788 12420 10805 12484
rect 10869 12420 10886 12484
rect 10950 12420 10967 12484
rect 11031 12420 11048 12484
rect 11112 12420 11129 12484
rect 11193 12420 11210 12484
rect 11274 12420 11291 12484
rect 11355 12420 11372 12484
rect 11436 12420 11453 12484
rect 11517 12420 11534 12484
rect 11598 12420 11615 12484
rect 11679 12420 11696 12484
rect 11760 12420 11777 12484
rect 11841 12420 11858 12484
rect 11922 12420 11939 12484
rect 12003 12420 12020 12484
rect 12084 12420 12101 12484
rect 12165 12420 12182 12484
rect 12246 12420 12263 12484
rect 12327 12420 12344 12484
rect 12408 12420 12425 12484
rect 12489 12420 12506 12484
rect 12570 12420 12587 12484
rect 12651 12420 12668 12484
rect 12732 12420 12749 12484
rect 12813 12420 12830 12484
rect 12894 12420 12911 12484
rect 12975 12420 12992 12484
rect 13056 12420 13073 12484
rect 13137 12420 13154 12484
rect 13218 12420 13235 12484
rect 13299 12420 13316 12484
rect 13380 12420 13397 12484
rect 13461 12420 13478 12484
rect 13542 12420 13559 12484
rect 13623 12420 13640 12484
rect 13704 12420 13721 12484
rect 13785 12420 13802 12484
rect 13866 12420 13883 12484
rect 13947 12420 13964 12484
rect 14028 12420 14045 12484
rect 14109 12420 14126 12484
rect 14190 12420 14207 12484
rect 14271 12420 14288 12484
rect 14352 12420 14369 12484
rect 14433 12420 14451 12484
rect 14515 12420 14533 12484
rect 14597 12420 14615 12484
rect 14679 12420 14697 12484
rect 14761 12420 14779 12484
rect 14843 12420 14861 12484
rect 14925 12420 14931 12484
rect 10151 12418 14931 12420
rect 120 4484 4900 4486
rect 120 4420 126 4484
rect 190 4420 207 4484
rect 271 4420 288 4484
rect 352 4420 369 4484
rect 433 4420 450 4484
rect 514 4420 531 4484
rect 595 4420 612 4484
rect 676 4420 693 4484
rect 757 4420 774 4484
rect 838 4420 855 4484
rect 919 4420 936 4484
rect 1000 4420 1017 4484
rect 1081 4420 1098 4484
rect 1162 4420 1179 4484
rect 1243 4420 1260 4484
rect 1324 4420 1341 4484
rect 1405 4420 1422 4484
rect 1486 4420 1503 4484
rect 1567 4420 1584 4484
rect 1648 4420 1665 4484
rect 1729 4420 1746 4484
rect 1810 4420 1827 4484
rect 1891 4420 1908 4484
rect 1972 4420 1989 4484
rect 2053 4420 2070 4484
rect 2134 4420 2151 4484
rect 2215 4420 2232 4484
rect 2296 4420 2313 4484
rect 2377 4420 2394 4484
rect 2458 4420 2475 4484
rect 2539 4420 2556 4484
rect 2620 4420 2637 4484
rect 2701 4420 2718 4484
rect 2782 4420 2799 4484
rect 2863 4420 2880 4484
rect 2944 4420 2961 4484
rect 3025 4420 3042 4484
rect 3106 4420 3123 4484
rect 3187 4420 3204 4484
rect 3268 4420 3285 4484
rect 3349 4420 3366 4484
rect 3430 4420 3447 4484
rect 3511 4420 3528 4484
rect 3592 4420 3609 4484
rect 3673 4420 3690 4484
rect 3754 4420 3771 4484
rect 3835 4420 3852 4484
rect 3916 4420 3933 4484
rect 3997 4420 4014 4484
rect 4078 4420 4095 4484
rect 4159 4420 4176 4484
rect 4240 4420 4257 4484
rect 4321 4420 4338 4484
rect 4402 4420 4420 4484
rect 4484 4420 4502 4484
rect 4566 4420 4584 4484
rect 4648 4420 4666 4484
rect 4730 4420 4748 4484
rect 4812 4420 4830 4484
rect 4894 4420 4900 4484
rect 120 4398 4900 4420
rect 120 4334 126 4398
rect 190 4334 207 4398
rect 271 4334 288 4398
rect 352 4334 369 4398
rect 433 4334 450 4398
rect 514 4334 531 4398
rect 595 4334 612 4398
rect 676 4334 693 4398
rect 757 4334 774 4398
rect 838 4334 855 4398
rect 919 4334 936 4398
rect 1000 4334 1017 4398
rect 1081 4334 1098 4398
rect 1162 4334 1179 4398
rect 1243 4334 1260 4398
rect 1324 4334 1341 4398
rect 1405 4334 1422 4398
rect 1486 4334 1503 4398
rect 1567 4334 1584 4398
rect 1648 4334 1665 4398
rect 1729 4334 1746 4398
rect 1810 4334 1827 4398
rect 1891 4334 1908 4398
rect 1972 4334 1989 4398
rect 2053 4334 2070 4398
rect 2134 4334 2151 4398
rect 2215 4334 2232 4398
rect 2296 4334 2313 4398
rect 2377 4334 2394 4398
rect 2458 4334 2475 4398
rect 2539 4334 2556 4398
rect 2620 4334 2637 4398
rect 2701 4334 2718 4398
rect 2782 4334 2799 4398
rect 2863 4334 2880 4398
rect 2944 4334 2961 4398
rect 3025 4334 3042 4398
rect 3106 4334 3123 4398
rect 3187 4334 3204 4398
rect 3268 4334 3285 4398
rect 3349 4334 3366 4398
rect 3430 4334 3447 4398
rect 3511 4334 3528 4398
rect 3592 4334 3609 4398
rect 3673 4334 3690 4398
rect 3754 4334 3771 4398
rect 3835 4334 3852 4398
rect 3916 4334 3933 4398
rect 3997 4334 4014 4398
rect 4078 4334 4095 4398
rect 4159 4334 4176 4398
rect 4240 4334 4257 4398
rect 4321 4334 4338 4398
rect 4402 4334 4420 4398
rect 4484 4334 4502 4398
rect 4566 4334 4584 4398
rect 4648 4334 4666 4398
rect 4730 4334 4748 4398
rect 4812 4334 4830 4398
rect 4894 4334 4900 4398
rect 120 4312 4900 4334
rect 120 4248 126 4312
rect 190 4248 207 4312
rect 271 4248 288 4312
rect 352 4248 369 4312
rect 433 4248 450 4312
rect 514 4248 531 4312
rect 595 4248 612 4312
rect 676 4248 693 4312
rect 757 4248 774 4312
rect 838 4248 855 4312
rect 919 4248 936 4312
rect 1000 4248 1017 4312
rect 1081 4248 1098 4312
rect 1162 4248 1179 4312
rect 1243 4248 1260 4312
rect 1324 4248 1341 4312
rect 1405 4248 1422 4312
rect 1486 4248 1503 4312
rect 1567 4248 1584 4312
rect 1648 4248 1665 4312
rect 1729 4248 1746 4312
rect 1810 4248 1827 4312
rect 1891 4248 1908 4312
rect 1972 4248 1989 4312
rect 2053 4248 2070 4312
rect 2134 4248 2151 4312
rect 2215 4248 2232 4312
rect 2296 4248 2313 4312
rect 2377 4248 2394 4312
rect 2458 4248 2475 4312
rect 2539 4248 2556 4312
rect 2620 4248 2637 4312
rect 2701 4248 2718 4312
rect 2782 4248 2799 4312
rect 2863 4248 2880 4312
rect 2944 4248 2961 4312
rect 3025 4248 3042 4312
rect 3106 4248 3123 4312
rect 3187 4248 3204 4312
rect 3268 4248 3285 4312
rect 3349 4248 3366 4312
rect 3430 4248 3447 4312
rect 3511 4248 3528 4312
rect 3592 4248 3609 4312
rect 3673 4248 3690 4312
rect 3754 4248 3771 4312
rect 3835 4248 3852 4312
rect 3916 4248 3933 4312
rect 3997 4248 4014 4312
rect 4078 4248 4095 4312
rect 4159 4248 4176 4312
rect 4240 4248 4257 4312
rect 4321 4248 4338 4312
rect 4402 4248 4420 4312
rect 4484 4248 4502 4312
rect 4566 4248 4584 4312
rect 4648 4248 4666 4312
rect 4730 4248 4748 4312
rect 4812 4248 4830 4312
rect 4894 4248 4900 4312
rect 120 4226 4900 4248
rect 120 4162 126 4226
rect 190 4162 207 4226
rect 271 4162 288 4226
rect 352 4162 369 4226
rect 433 4162 450 4226
rect 514 4162 531 4226
rect 595 4162 612 4226
rect 676 4162 693 4226
rect 757 4162 774 4226
rect 838 4162 855 4226
rect 919 4162 936 4226
rect 1000 4162 1017 4226
rect 1081 4162 1098 4226
rect 1162 4162 1179 4226
rect 1243 4162 1260 4226
rect 1324 4162 1341 4226
rect 1405 4162 1422 4226
rect 1486 4162 1503 4226
rect 1567 4162 1584 4226
rect 1648 4162 1665 4226
rect 1729 4162 1746 4226
rect 1810 4162 1827 4226
rect 1891 4162 1908 4226
rect 1972 4162 1989 4226
rect 2053 4162 2070 4226
rect 2134 4162 2151 4226
rect 2215 4162 2232 4226
rect 2296 4162 2313 4226
rect 2377 4162 2394 4226
rect 2458 4162 2475 4226
rect 2539 4162 2556 4226
rect 2620 4162 2637 4226
rect 2701 4162 2718 4226
rect 2782 4162 2799 4226
rect 2863 4162 2880 4226
rect 2944 4162 2961 4226
rect 3025 4162 3042 4226
rect 3106 4162 3123 4226
rect 3187 4162 3204 4226
rect 3268 4162 3285 4226
rect 3349 4162 3366 4226
rect 3430 4162 3447 4226
rect 3511 4162 3528 4226
rect 3592 4162 3609 4226
rect 3673 4162 3690 4226
rect 3754 4162 3771 4226
rect 3835 4162 3852 4226
rect 3916 4162 3933 4226
rect 3997 4162 4014 4226
rect 4078 4162 4095 4226
rect 4159 4162 4176 4226
rect 4240 4162 4257 4226
rect 4321 4162 4338 4226
rect 4402 4162 4420 4226
rect 4484 4162 4502 4226
rect 4566 4162 4584 4226
rect 4648 4162 4666 4226
rect 4730 4162 4748 4226
rect 4812 4162 4830 4226
rect 4894 4162 4900 4226
rect 120 4140 4900 4162
rect 120 4076 126 4140
rect 190 4076 207 4140
rect 271 4076 288 4140
rect 352 4076 369 4140
rect 433 4076 450 4140
rect 514 4076 531 4140
rect 595 4076 612 4140
rect 676 4076 693 4140
rect 757 4076 774 4140
rect 838 4076 855 4140
rect 919 4076 936 4140
rect 1000 4076 1017 4140
rect 1081 4076 1098 4140
rect 1162 4076 1179 4140
rect 1243 4076 1260 4140
rect 1324 4076 1341 4140
rect 1405 4076 1422 4140
rect 1486 4076 1503 4140
rect 1567 4076 1584 4140
rect 1648 4076 1665 4140
rect 1729 4076 1746 4140
rect 1810 4076 1827 4140
rect 1891 4076 1908 4140
rect 1972 4076 1989 4140
rect 2053 4076 2070 4140
rect 2134 4076 2151 4140
rect 2215 4076 2232 4140
rect 2296 4076 2313 4140
rect 2377 4076 2394 4140
rect 2458 4076 2475 4140
rect 2539 4076 2556 4140
rect 2620 4076 2637 4140
rect 2701 4076 2718 4140
rect 2782 4076 2799 4140
rect 2863 4076 2880 4140
rect 2944 4076 2961 4140
rect 3025 4076 3042 4140
rect 3106 4076 3123 4140
rect 3187 4076 3204 4140
rect 3268 4076 3285 4140
rect 3349 4076 3366 4140
rect 3430 4076 3447 4140
rect 3511 4076 3528 4140
rect 3592 4076 3609 4140
rect 3673 4076 3690 4140
rect 3754 4076 3771 4140
rect 3835 4076 3852 4140
rect 3916 4076 3933 4140
rect 3997 4076 4014 4140
rect 4078 4076 4095 4140
rect 4159 4076 4176 4140
rect 4240 4076 4257 4140
rect 4321 4076 4338 4140
rect 4402 4076 4420 4140
rect 4484 4076 4502 4140
rect 4566 4076 4584 4140
rect 4648 4076 4666 4140
rect 4730 4076 4748 4140
rect 4812 4076 4830 4140
rect 4894 4076 4900 4140
rect 120 4054 4900 4076
rect 120 3990 126 4054
rect 190 3990 207 4054
rect 271 3990 288 4054
rect 352 3990 369 4054
rect 433 3990 450 4054
rect 514 3990 531 4054
rect 595 3990 612 4054
rect 676 3990 693 4054
rect 757 3990 774 4054
rect 838 3990 855 4054
rect 919 3990 936 4054
rect 1000 3990 1017 4054
rect 1081 3990 1098 4054
rect 1162 3990 1179 4054
rect 1243 3990 1260 4054
rect 1324 3990 1341 4054
rect 1405 3990 1422 4054
rect 1486 3990 1503 4054
rect 1567 3990 1584 4054
rect 1648 3990 1665 4054
rect 1729 3990 1746 4054
rect 1810 3990 1827 4054
rect 1891 3990 1908 4054
rect 1972 3990 1989 4054
rect 2053 3990 2070 4054
rect 2134 3990 2151 4054
rect 2215 3990 2232 4054
rect 2296 3990 2313 4054
rect 2377 3990 2394 4054
rect 2458 3990 2475 4054
rect 2539 3990 2556 4054
rect 2620 3990 2637 4054
rect 2701 3990 2718 4054
rect 2782 3990 2799 4054
rect 2863 3990 2880 4054
rect 2944 3990 2961 4054
rect 3025 3990 3042 4054
rect 3106 3990 3123 4054
rect 3187 3990 3204 4054
rect 3268 3990 3285 4054
rect 3349 3990 3366 4054
rect 3430 3990 3447 4054
rect 3511 3990 3528 4054
rect 3592 3990 3609 4054
rect 3673 3990 3690 4054
rect 3754 3990 3771 4054
rect 3835 3990 3852 4054
rect 3916 3990 3933 4054
rect 3997 3990 4014 4054
rect 4078 3990 4095 4054
rect 4159 3990 4176 4054
rect 4240 3990 4257 4054
rect 4321 3990 4338 4054
rect 4402 3990 4420 4054
rect 4484 3990 4502 4054
rect 4566 3990 4584 4054
rect 4648 3990 4666 4054
rect 4730 3990 4748 4054
rect 4812 3990 4830 4054
rect 4894 3990 4900 4054
rect 120 3968 4900 3990
rect 120 3904 126 3968
rect 190 3904 207 3968
rect 271 3904 288 3968
rect 352 3904 369 3968
rect 433 3904 450 3968
rect 514 3904 531 3968
rect 595 3904 612 3968
rect 676 3904 693 3968
rect 757 3904 774 3968
rect 838 3904 855 3968
rect 919 3904 936 3968
rect 1000 3904 1017 3968
rect 1081 3904 1098 3968
rect 1162 3904 1179 3968
rect 1243 3904 1260 3968
rect 1324 3904 1341 3968
rect 1405 3904 1422 3968
rect 1486 3904 1503 3968
rect 1567 3904 1584 3968
rect 1648 3904 1665 3968
rect 1729 3904 1746 3968
rect 1810 3904 1827 3968
rect 1891 3904 1908 3968
rect 1972 3904 1989 3968
rect 2053 3904 2070 3968
rect 2134 3904 2151 3968
rect 2215 3904 2232 3968
rect 2296 3904 2313 3968
rect 2377 3904 2394 3968
rect 2458 3904 2475 3968
rect 2539 3904 2556 3968
rect 2620 3904 2637 3968
rect 2701 3904 2718 3968
rect 2782 3904 2799 3968
rect 2863 3904 2880 3968
rect 2944 3904 2961 3968
rect 3025 3904 3042 3968
rect 3106 3904 3123 3968
rect 3187 3904 3204 3968
rect 3268 3904 3285 3968
rect 3349 3904 3366 3968
rect 3430 3904 3447 3968
rect 3511 3904 3528 3968
rect 3592 3904 3609 3968
rect 3673 3904 3690 3968
rect 3754 3904 3771 3968
rect 3835 3904 3852 3968
rect 3916 3904 3933 3968
rect 3997 3904 4014 3968
rect 4078 3904 4095 3968
rect 4159 3904 4176 3968
rect 4240 3904 4257 3968
rect 4321 3904 4338 3968
rect 4402 3904 4420 3968
rect 4484 3904 4502 3968
rect 4566 3904 4584 3968
rect 4648 3904 4666 3968
rect 4730 3904 4748 3968
rect 4812 3904 4830 3968
rect 4894 3904 4900 3968
rect 120 3882 4900 3904
rect 120 3818 126 3882
rect 190 3818 207 3882
rect 271 3818 288 3882
rect 352 3818 369 3882
rect 433 3818 450 3882
rect 514 3818 531 3882
rect 595 3818 612 3882
rect 676 3818 693 3882
rect 757 3818 774 3882
rect 838 3818 855 3882
rect 919 3818 936 3882
rect 1000 3818 1017 3882
rect 1081 3818 1098 3882
rect 1162 3818 1179 3882
rect 1243 3818 1260 3882
rect 1324 3818 1341 3882
rect 1405 3818 1422 3882
rect 1486 3818 1503 3882
rect 1567 3818 1584 3882
rect 1648 3818 1665 3882
rect 1729 3818 1746 3882
rect 1810 3818 1827 3882
rect 1891 3818 1908 3882
rect 1972 3818 1989 3882
rect 2053 3818 2070 3882
rect 2134 3818 2151 3882
rect 2215 3818 2232 3882
rect 2296 3818 2313 3882
rect 2377 3818 2394 3882
rect 2458 3818 2475 3882
rect 2539 3818 2556 3882
rect 2620 3818 2637 3882
rect 2701 3818 2718 3882
rect 2782 3818 2799 3882
rect 2863 3818 2880 3882
rect 2944 3818 2961 3882
rect 3025 3818 3042 3882
rect 3106 3818 3123 3882
rect 3187 3818 3204 3882
rect 3268 3818 3285 3882
rect 3349 3818 3366 3882
rect 3430 3818 3447 3882
rect 3511 3818 3528 3882
rect 3592 3818 3609 3882
rect 3673 3818 3690 3882
rect 3754 3818 3771 3882
rect 3835 3818 3852 3882
rect 3916 3818 3933 3882
rect 3997 3818 4014 3882
rect 4078 3818 4095 3882
rect 4159 3818 4176 3882
rect 4240 3818 4257 3882
rect 4321 3818 4338 3882
rect 4402 3818 4420 3882
rect 4484 3818 4502 3882
rect 4566 3818 4584 3882
rect 4648 3818 4666 3882
rect 4730 3818 4748 3882
rect 4812 3818 4830 3882
rect 4894 3818 4900 3882
rect 120 3796 4900 3818
rect 120 3732 126 3796
rect 190 3732 207 3796
rect 271 3732 288 3796
rect 352 3732 369 3796
rect 433 3732 450 3796
rect 514 3732 531 3796
rect 595 3732 612 3796
rect 676 3732 693 3796
rect 757 3732 774 3796
rect 838 3732 855 3796
rect 919 3732 936 3796
rect 1000 3732 1017 3796
rect 1081 3732 1098 3796
rect 1162 3732 1179 3796
rect 1243 3732 1260 3796
rect 1324 3732 1341 3796
rect 1405 3732 1422 3796
rect 1486 3732 1503 3796
rect 1567 3732 1584 3796
rect 1648 3732 1665 3796
rect 1729 3732 1746 3796
rect 1810 3732 1827 3796
rect 1891 3732 1908 3796
rect 1972 3732 1989 3796
rect 2053 3732 2070 3796
rect 2134 3732 2151 3796
rect 2215 3732 2232 3796
rect 2296 3732 2313 3796
rect 2377 3732 2394 3796
rect 2458 3732 2475 3796
rect 2539 3732 2556 3796
rect 2620 3732 2637 3796
rect 2701 3732 2718 3796
rect 2782 3732 2799 3796
rect 2863 3732 2880 3796
rect 2944 3732 2961 3796
rect 3025 3732 3042 3796
rect 3106 3732 3123 3796
rect 3187 3732 3204 3796
rect 3268 3732 3285 3796
rect 3349 3732 3366 3796
rect 3430 3732 3447 3796
rect 3511 3732 3528 3796
rect 3592 3732 3609 3796
rect 3673 3732 3690 3796
rect 3754 3732 3771 3796
rect 3835 3732 3852 3796
rect 3916 3732 3933 3796
rect 3997 3732 4014 3796
rect 4078 3732 4095 3796
rect 4159 3732 4176 3796
rect 4240 3732 4257 3796
rect 4321 3732 4338 3796
rect 4402 3732 4420 3796
rect 4484 3732 4502 3796
rect 4566 3732 4584 3796
rect 4648 3732 4666 3796
rect 4730 3732 4748 3796
rect 4812 3732 4830 3796
rect 4894 3732 4900 3796
rect 120 3710 4900 3732
rect 120 3646 126 3710
rect 190 3646 207 3710
rect 271 3646 288 3710
rect 352 3646 369 3710
rect 433 3646 450 3710
rect 514 3646 531 3710
rect 595 3646 612 3710
rect 676 3646 693 3710
rect 757 3646 774 3710
rect 838 3646 855 3710
rect 919 3646 936 3710
rect 1000 3646 1017 3710
rect 1081 3646 1098 3710
rect 1162 3646 1179 3710
rect 1243 3646 1260 3710
rect 1324 3646 1341 3710
rect 1405 3646 1422 3710
rect 1486 3646 1503 3710
rect 1567 3646 1584 3710
rect 1648 3646 1665 3710
rect 1729 3646 1746 3710
rect 1810 3646 1827 3710
rect 1891 3646 1908 3710
rect 1972 3646 1989 3710
rect 2053 3646 2070 3710
rect 2134 3646 2151 3710
rect 2215 3646 2232 3710
rect 2296 3646 2313 3710
rect 2377 3646 2394 3710
rect 2458 3646 2475 3710
rect 2539 3646 2556 3710
rect 2620 3646 2637 3710
rect 2701 3646 2718 3710
rect 2782 3646 2799 3710
rect 2863 3646 2880 3710
rect 2944 3646 2961 3710
rect 3025 3646 3042 3710
rect 3106 3646 3123 3710
rect 3187 3646 3204 3710
rect 3268 3646 3285 3710
rect 3349 3646 3366 3710
rect 3430 3646 3447 3710
rect 3511 3646 3528 3710
rect 3592 3646 3609 3710
rect 3673 3646 3690 3710
rect 3754 3646 3771 3710
rect 3835 3646 3852 3710
rect 3916 3646 3933 3710
rect 3997 3646 4014 3710
rect 4078 3646 4095 3710
rect 4159 3646 4176 3710
rect 4240 3646 4257 3710
rect 4321 3646 4338 3710
rect 4402 3646 4420 3710
rect 4484 3646 4502 3710
rect 4566 3646 4584 3710
rect 4648 3646 4666 3710
rect 4730 3646 4748 3710
rect 4812 3646 4830 3710
rect 4894 3646 4900 3710
rect 120 3624 4900 3646
rect 120 3560 126 3624
rect 190 3560 207 3624
rect 271 3560 288 3624
rect 352 3560 369 3624
rect 433 3560 450 3624
rect 514 3560 531 3624
rect 595 3560 612 3624
rect 676 3560 693 3624
rect 757 3560 774 3624
rect 838 3560 855 3624
rect 919 3560 936 3624
rect 1000 3560 1017 3624
rect 1081 3560 1098 3624
rect 1162 3560 1179 3624
rect 1243 3560 1260 3624
rect 1324 3560 1341 3624
rect 1405 3560 1422 3624
rect 1486 3560 1503 3624
rect 1567 3560 1584 3624
rect 1648 3560 1665 3624
rect 1729 3560 1746 3624
rect 1810 3560 1827 3624
rect 1891 3560 1908 3624
rect 1972 3560 1989 3624
rect 2053 3560 2070 3624
rect 2134 3560 2151 3624
rect 2215 3560 2232 3624
rect 2296 3560 2313 3624
rect 2377 3560 2394 3624
rect 2458 3560 2475 3624
rect 2539 3560 2556 3624
rect 2620 3560 2637 3624
rect 2701 3560 2718 3624
rect 2782 3560 2799 3624
rect 2863 3560 2880 3624
rect 2944 3560 2961 3624
rect 3025 3560 3042 3624
rect 3106 3560 3123 3624
rect 3187 3560 3204 3624
rect 3268 3560 3285 3624
rect 3349 3560 3366 3624
rect 3430 3560 3447 3624
rect 3511 3560 3528 3624
rect 3592 3560 3609 3624
rect 3673 3560 3690 3624
rect 3754 3560 3771 3624
rect 3835 3560 3852 3624
rect 3916 3560 3933 3624
rect 3997 3560 4014 3624
rect 4078 3560 4095 3624
rect 4159 3560 4176 3624
rect 4240 3560 4257 3624
rect 4321 3560 4338 3624
rect 4402 3560 4420 3624
rect 4484 3560 4502 3624
rect 4566 3560 4584 3624
rect 4648 3560 4666 3624
rect 4730 3560 4748 3624
rect 4812 3560 4830 3624
rect 4894 3560 4900 3624
rect 120 3558 4900 3560
rect 10151 4484 14931 4486
rect 10151 4420 10157 4484
rect 10221 4420 10238 4484
rect 10302 4420 10319 4484
rect 10383 4420 10400 4484
rect 10464 4420 10481 4484
rect 10545 4420 10562 4484
rect 10626 4420 10643 4484
rect 10707 4420 10724 4484
rect 10788 4420 10805 4484
rect 10869 4420 10886 4484
rect 10950 4420 10967 4484
rect 11031 4420 11048 4484
rect 11112 4420 11129 4484
rect 11193 4420 11210 4484
rect 11274 4420 11291 4484
rect 11355 4420 11372 4484
rect 11436 4420 11453 4484
rect 11517 4420 11534 4484
rect 11598 4420 11615 4484
rect 11679 4420 11696 4484
rect 11760 4420 11777 4484
rect 11841 4420 11858 4484
rect 11922 4420 11939 4484
rect 12003 4420 12020 4484
rect 12084 4420 12101 4484
rect 12165 4420 12182 4484
rect 12246 4420 12263 4484
rect 12327 4420 12344 4484
rect 12408 4420 12425 4484
rect 12489 4420 12506 4484
rect 12570 4420 12587 4484
rect 12651 4420 12668 4484
rect 12732 4420 12749 4484
rect 12813 4420 12830 4484
rect 12894 4420 12911 4484
rect 12975 4420 12992 4484
rect 13056 4420 13073 4484
rect 13137 4420 13154 4484
rect 13218 4420 13235 4484
rect 13299 4420 13316 4484
rect 13380 4420 13397 4484
rect 13461 4420 13478 4484
rect 13542 4420 13559 4484
rect 13623 4420 13640 4484
rect 13704 4420 13721 4484
rect 13785 4420 13802 4484
rect 13866 4420 13883 4484
rect 13947 4420 13964 4484
rect 14028 4420 14045 4484
rect 14109 4420 14126 4484
rect 14190 4420 14207 4484
rect 14271 4420 14288 4484
rect 14352 4420 14369 4484
rect 14433 4420 14451 4484
rect 14515 4420 14533 4484
rect 14597 4420 14615 4484
rect 14679 4420 14697 4484
rect 14761 4420 14779 4484
rect 14843 4420 14861 4484
rect 14925 4420 14931 4484
rect 10151 4398 14931 4420
rect 10151 4334 10157 4398
rect 10221 4334 10238 4398
rect 10302 4334 10319 4398
rect 10383 4334 10400 4398
rect 10464 4334 10481 4398
rect 10545 4334 10562 4398
rect 10626 4334 10643 4398
rect 10707 4334 10724 4398
rect 10788 4334 10805 4398
rect 10869 4334 10886 4398
rect 10950 4334 10967 4398
rect 11031 4334 11048 4398
rect 11112 4334 11129 4398
rect 11193 4334 11210 4398
rect 11274 4334 11291 4398
rect 11355 4334 11372 4398
rect 11436 4334 11453 4398
rect 11517 4334 11534 4398
rect 11598 4334 11615 4398
rect 11679 4334 11696 4398
rect 11760 4334 11777 4398
rect 11841 4334 11858 4398
rect 11922 4334 11939 4398
rect 12003 4334 12020 4398
rect 12084 4334 12101 4398
rect 12165 4334 12182 4398
rect 12246 4334 12263 4398
rect 12327 4334 12344 4398
rect 12408 4334 12425 4398
rect 12489 4334 12506 4398
rect 12570 4334 12587 4398
rect 12651 4334 12668 4398
rect 12732 4334 12749 4398
rect 12813 4334 12830 4398
rect 12894 4334 12911 4398
rect 12975 4334 12992 4398
rect 13056 4334 13073 4398
rect 13137 4334 13154 4398
rect 13218 4334 13235 4398
rect 13299 4334 13316 4398
rect 13380 4334 13397 4398
rect 13461 4334 13478 4398
rect 13542 4334 13559 4398
rect 13623 4334 13640 4398
rect 13704 4334 13721 4398
rect 13785 4334 13802 4398
rect 13866 4334 13883 4398
rect 13947 4334 13964 4398
rect 14028 4334 14045 4398
rect 14109 4334 14126 4398
rect 14190 4334 14207 4398
rect 14271 4334 14288 4398
rect 14352 4334 14369 4398
rect 14433 4334 14451 4398
rect 14515 4334 14533 4398
rect 14597 4334 14615 4398
rect 14679 4334 14697 4398
rect 14761 4334 14779 4398
rect 14843 4334 14861 4398
rect 14925 4334 14931 4398
rect 10151 4312 14931 4334
rect 10151 4248 10157 4312
rect 10221 4248 10238 4312
rect 10302 4248 10319 4312
rect 10383 4248 10400 4312
rect 10464 4248 10481 4312
rect 10545 4248 10562 4312
rect 10626 4248 10643 4312
rect 10707 4248 10724 4312
rect 10788 4248 10805 4312
rect 10869 4248 10886 4312
rect 10950 4248 10967 4312
rect 11031 4248 11048 4312
rect 11112 4248 11129 4312
rect 11193 4248 11210 4312
rect 11274 4248 11291 4312
rect 11355 4248 11372 4312
rect 11436 4248 11453 4312
rect 11517 4248 11534 4312
rect 11598 4248 11615 4312
rect 11679 4248 11696 4312
rect 11760 4248 11777 4312
rect 11841 4248 11858 4312
rect 11922 4248 11939 4312
rect 12003 4248 12020 4312
rect 12084 4248 12101 4312
rect 12165 4248 12182 4312
rect 12246 4248 12263 4312
rect 12327 4248 12344 4312
rect 12408 4248 12425 4312
rect 12489 4248 12506 4312
rect 12570 4248 12587 4312
rect 12651 4248 12668 4312
rect 12732 4248 12749 4312
rect 12813 4248 12830 4312
rect 12894 4248 12911 4312
rect 12975 4248 12992 4312
rect 13056 4248 13073 4312
rect 13137 4248 13154 4312
rect 13218 4248 13235 4312
rect 13299 4248 13316 4312
rect 13380 4248 13397 4312
rect 13461 4248 13478 4312
rect 13542 4248 13559 4312
rect 13623 4248 13640 4312
rect 13704 4248 13721 4312
rect 13785 4248 13802 4312
rect 13866 4248 13883 4312
rect 13947 4248 13964 4312
rect 14028 4248 14045 4312
rect 14109 4248 14126 4312
rect 14190 4248 14207 4312
rect 14271 4248 14288 4312
rect 14352 4248 14369 4312
rect 14433 4248 14451 4312
rect 14515 4248 14533 4312
rect 14597 4248 14615 4312
rect 14679 4248 14697 4312
rect 14761 4248 14779 4312
rect 14843 4248 14861 4312
rect 14925 4248 14931 4312
rect 10151 4226 14931 4248
rect 10151 4162 10157 4226
rect 10221 4162 10238 4226
rect 10302 4162 10319 4226
rect 10383 4162 10400 4226
rect 10464 4162 10481 4226
rect 10545 4162 10562 4226
rect 10626 4162 10643 4226
rect 10707 4162 10724 4226
rect 10788 4162 10805 4226
rect 10869 4162 10886 4226
rect 10950 4162 10967 4226
rect 11031 4162 11048 4226
rect 11112 4162 11129 4226
rect 11193 4162 11210 4226
rect 11274 4162 11291 4226
rect 11355 4162 11372 4226
rect 11436 4162 11453 4226
rect 11517 4162 11534 4226
rect 11598 4162 11615 4226
rect 11679 4162 11696 4226
rect 11760 4162 11777 4226
rect 11841 4162 11858 4226
rect 11922 4162 11939 4226
rect 12003 4162 12020 4226
rect 12084 4162 12101 4226
rect 12165 4162 12182 4226
rect 12246 4162 12263 4226
rect 12327 4162 12344 4226
rect 12408 4162 12425 4226
rect 12489 4162 12506 4226
rect 12570 4162 12587 4226
rect 12651 4162 12668 4226
rect 12732 4162 12749 4226
rect 12813 4162 12830 4226
rect 12894 4162 12911 4226
rect 12975 4162 12992 4226
rect 13056 4162 13073 4226
rect 13137 4162 13154 4226
rect 13218 4162 13235 4226
rect 13299 4162 13316 4226
rect 13380 4162 13397 4226
rect 13461 4162 13478 4226
rect 13542 4162 13559 4226
rect 13623 4162 13640 4226
rect 13704 4162 13721 4226
rect 13785 4162 13802 4226
rect 13866 4162 13883 4226
rect 13947 4162 13964 4226
rect 14028 4162 14045 4226
rect 14109 4162 14126 4226
rect 14190 4162 14207 4226
rect 14271 4162 14288 4226
rect 14352 4162 14369 4226
rect 14433 4162 14451 4226
rect 14515 4162 14533 4226
rect 14597 4162 14615 4226
rect 14679 4162 14697 4226
rect 14761 4162 14779 4226
rect 14843 4162 14861 4226
rect 14925 4162 14931 4226
rect 10151 4140 14931 4162
rect 10151 4076 10157 4140
rect 10221 4076 10238 4140
rect 10302 4076 10319 4140
rect 10383 4076 10400 4140
rect 10464 4076 10481 4140
rect 10545 4076 10562 4140
rect 10626 4076 10643 4140
rect 10707 4076 10724 4140
rect 10788 4076 10805 4140
rect 10869 4076 10886 4140
rect 10950 4076 10967 4140
rect 11031 4076 11048 4140
rect 11112 4076 11129 4140
rect 11193 4076 11210 4140
rect 11274 4076 11291 4140
rect 11355 4076 11372 4140
rect 11436 4076 11453 4140
rect 11517 4076 11534 4140
rect 11598 4076 11615 4140
rect 11679 4076 11696 4140
rect 11760 4076 11777 4140
rect 11841 4076 11858 4140
rect 11922 4076 11939 4140
rect 12003 4076 12020 4140
rect 12084 4076 12101 4140
rect 12165 4076 12182 4140
rect 12246 4076 12263 4140
rect 12327 4076 12344 4140
rect 12408 4076 12425 4140
rect 12489 4076 12506 4140
rect 12570 4076 12587 4140
rect 12651 4076 12668 4140
rect 12732 4076 12749 4140
rect 12813 4076 12830 4140
rect 12894 4076 12911 4140
rect 12975 4076 12992 4140
rect 13056 4076 13073 4140
rect 13137 4076 13154 4140
rect 13218 4076 13235 4140
rect 13299 4076 13316 4140
rect 13380 4076 13397 4140
rect 13461 4076 13478 4140
rect 13542 4076 13559 4140
rect 13623 4076 13640 4140
rect 13704 4076 13721 4140
rect 13785 4076 13802 4140
rect 13866 4076 13883 4140
rect 13947 4076 13964 4140
rect 14028 4076 14045 4140
rect 14109 4076 14126 4140
rect 14190 4076 14207 4140
rect 14271 4076 14288 4140
rect 14352 4076 14369 4140
rect 14433 4076 14451 4140
rect 14515 4076 14533 4140
rect 14597 4076 14615 4140
rect 14679 4076 14697 4140
rect 14761 4076 14779 4140
rect 14843 4076 14861 4140
rect 14925 4076 14931 4140
rect 10151 4054 14931 4076
rect 10151 3990 10157 4054
rect 10221 3990 10238 4054
rect 10302 3990 10319 4054
rect 10383 3990 10400 4054
rect 10464 3990 10481 4054
rect 10545 3990 10562 4054
rect 10626 3990 10643 4054
rect 10707 3990 10724 4054
rect 10788 3990 10805 4054
rect 10869 3990 10886 4054
rect 10950 3990 10967 4054
rect 11031 3990 11048 4054
rect 11112 3990 11129 4054
rect 11193 3990 11210 4054
rect 11274 3990 11291 4054
rect 11355 3990 11372 4054
rect 11436 3990 11453 4054
rect 11517 3990 11534 4054
rect 11598 3990 11615 4054
rect 11679 3990 11696 4054
rect 11760 3990 11777 4054
rect 11841 3990 11858 4054
rect 11922 3990 11939 4054
rect 12003 3990 12020 4054
rect 12084 3990 12101 4054
rect 12165 3990 12182 4054
rect 12246 3990 12263 4054
rect 12327 3990 12344 4054
rect 12408 3990 12425 4054
rect 12489 3990 12506 4054
rect 12570 3990 12587 4054
rect 12651 3990 12668 4054
rect 12732 3990 12749 4054
rect 12813 3990 12830 4054
rect 12894 3990 12911 4054
rect 12975 3990 12992 4054
rect 13056 3990 13073 4054
rect 13137 3990 13154 4054
rect 13218 3990 13235 4054
rect 13299 3990 13316 4054
rect 13380 3990 13397 4054
rect 13461 3990 13478 4054
rect 13542 3990 13559 4054
rect 13623 3990 13640 4054
rect 13704 3990 13721 4054
rect 13785 3990 13802 4054
rect 13866 3990 13883 4054
rect 13947 3990 13964 4054
rect 14028 3990 14045 4054
rect 14109 3990 14126 4054
rect 14190 3990 14207 4054
rect 14271 3990 14288 4054
rect 14352 3990 14369 4054
rect 14433 3990 14451 4054
rect 14515 3990 14533 4054
rect 14597 3990 14615 4054
rect 14679 3990 14697 4054
rect 14761 3990 14779 4054
rect 14843 3990 14861 4054
rect 14925 3990 14931 4054
rect 10151 3968 14931 3990
rect 10151 3904 10157 3968
rect 10221 3904 10238 3968
rect 10302 3904 10319 3968
rect 10383 3904 10400 3968
rect 10464 3904 10481 3968
rect 10545 3904 10562 3968
rect 10626 3904 10643 3968
rect 10707 3904 10724 3968
rect 10788 3904 10805 3968
rect 10869 3904 10886 3968
rect 10950 3904 10967 3968
rect 11031 3904 11048 3968
rect 11112 3904 11129 3968
rect 11193 3904 11210 3968
rect 11274 3904 11291 3968
rect 11355 3904 11372 3968
rect 11436 3904 11453 3968
rect 11517 3904 11534 3968
rect 11598 3904 11615 3968
rect 11679 3904 11696 3968
rect 11760 3904 11777 3968
rect 11841 3904 11858 3968
rect 11922 3904 11939 3968
rect 12003 3904 12020 3968
rect 12084 3904 12101 3968
rect 12165 3904 12182 3968
rect 12246 3904 12263 3968
rect 12327 3904 12344 3968
rect 12408 3904 12425 3968
rect 12489 3904 12506 3968
rect 12570 3904 12587 3968
rect 12651 3904 12668 3968
rect 12732 3904 12749 3968
rect 12813 3904 12830 3968
rect 12894 3904 12911 3968
rect 12975 3904 12992 3968
rect 13056 3904 13073 3968
rect 13137 3904 13154 3968
rect 13218 3904 13235 3968
rect 13299 3904 13316 3968
rect 13380 3904 13397 3968
rect 13461 3904 13478 3968
rect 13542 3904 13559 3968
rect 13623 3904 13640 3968
rect 13704 3904 13721 3968
rect 13785 3904 13802 3968
rect 13866 3904 13883 3968
rect 13947 3904 13964 3968
rect 14028 3904 14045 3968
rect 14109 3904 14126 3968
rect 14190 3904 14207 3968
rect 14271 3904 14288 3968
rect 14352 3904 14369 3968
rect 14433 3904 14451 3968
rect 14515 3904 14533 3968
rect 14597 3904 14615 3968
rect 14679 3904 14697 3968
rect 14761 3904 14779 3968
rect 14843 3904 14861 3968
rect 14925 3904 14931 3968
rect 10151 3882 14931 3904
rect 10151 3818 10157 3882
rect 10221 3818 10238 3882
rect 10302 3818 10319 3882
rect 10383 3818 10400 3882
rect 10464 3818 10481 3882
rect 10545 3818 10562 3882
rect 10626 3818 10643 3882
rect 10707 3818 10724 3882
rect 10788 3818 10805 3882
rect 10869 3818 10886 3882
rect 10950 3818 10967 3882
rect 11031 3818 11048 3882
rect 11112 3818 11129 3882
rect 11193 3818 11210 3882
rect 11274 3818 11291 3882
rect 11355 3818 11372 3882
rect 11436 3818 11453 3882
rect 11517 3818 11534 3882
rect 11598 3818 11615 3882
rect 11679 3818 11696 3882
rect 11760 3818 11777 3882
rect 11841 3818 11858 3882
rect 11922 3818 11939 3882
rect 12003 3818 12020 3882
rect 12084 3818 12101 3882
rect 12165 3818 12182 3882
rect 12246 3818 12263 3882
rect 12327 3818 12344 3882
rect 12408 3818 12425 3882
rect 12489 3818 12506 3882
rect 12570 3818 12587 3882
rect 12651 3818 12668 3882
rect 12732 3818 12749 3882
rect 12813 3818 12830 3882
rect 12894 3818 12911 3882
rect 12975 3818 12992 3882
rect 13056 3818 13073 3882
rect 13137 3818 13154 3882
rect 13218 3818 13235 3882
rect 13299 3818 13316 3882
rect 13380 3818 13397 3882
rect 13461 3818 13478 3882
rect 13542 3818 13559 3882
rect 13623 3818 13640 3882
rect 13704 3818 13721 3882
rect 13785 3818 13802 3882
rect 13866 3818 13883 3882
rect 13947 3818 13964 3882
rect 14028 3818 14045 3882
rect 14109 3818 14126 3882
rect 14190 3818 14207 3882
rect 14271 3818 14288 3882
rect 14352 3818 14369 3882
rect 14433 3818 14451 3882
rect 14515 3818 14533 3882
rect 14597 3818 14615 3882
rect 14679 3818 14697 3882
rect 14761 3818 14779 3882
rect 14843 3818 14861 3882
rect 14925 3818 14931 3882
rect 10151 3796 14931 3818
rect 10151 3732 10157 3796
rect 10221 3732 10238 3796
rect 10302 3732 10319 3796
rect 10383 3732 10400 3796
rect 10464 3732 10481 3796
rect 10545 3732 10562 3796
rect 10626 3732 10643 3796
rect 10707 3732 10724 3796
rect 10788 3732 10805 3796
rect 10869 3732 10886 3796
rect 10950 3732 10967 3796
rect 11031 3732 11048 3796
rect 11112 3732 11129 3796
rect 11193 3732 11210 3796
rect 11274 3732 11291 3796
rect 11355 3732 11372 3796
rect 11436 3732 11453 3796
rect 11517 3732 11534 3796
rect 11598 3732 11615 3796
rect 11679 3732 11696 3796
rect 11760 3732 11777 3796
rect 11841 3732 11858 3796
rect 11922 3732 11939 3796
rect 12003 3732 12020 3796
rect 12084 3732 12101 3796
rect 12165 3732 12182 3796
rect 12246 3732 12263 3796
rect 12327 3732 12344 3796
rect 12408 3732 12425 3796
rect 12489 3732 12506 3796
rect 12570 3732 12587 3796
rect 12651 3732 12668 3796
rect 12732 3732 12749 3796
rect 12813 3732 12830 3796
rect 12894 3732 12911 3796
rect 12975 3732 12992 3796
rect 13056 3732 13073 3796
rect 13137 3732 13154 3796
rect 13218 3732 13235 3796
rect 13299 3732 13316 3796
rect 13380 3732 13397 3796
rect 13461 3732 13478 3796
rect 13542 3732 13559 3796
rect 13623 3732 13640 3796
rect 13704 3732 13721 3796
rect 13785 3732 13802 3796
rect 13866 3732 13883 3796
rect 13947 3732 13964 3796
rect 14028 3732 14045 3796
rect 14109 3732 14126 3796
rect 14190 3732 14207 3796
rect 14271 3732 14288 3796
rect 14352 3732 14369 3796
rect 14433 3732 14451 3796
rect 14515 3732 14533 3796
rect 14597 3732 14615 3796
rect 14679 3732 14697 3796
rect 14761 3732 14779 3796
rect 14843 3732 14861 3796
rect 14925 3732 14931 3796
rect 10151 3710 14931 3732
rect 10151 3646 10157 3710
rect 10221 3646 10238 3710
rect 10302 3646 10319 3710
rect 10383 3646 10400 3710
rect 10464 3646 10481 3710
rect 10545 3646 10562 3710
rect 10626 3646 10643 3710
rect 10707 3646 10724 3710
rect 10788 3646 10805 3710
rect 10869 3646 10886 3710
rect 10950 3646 10967 3710
rect 11031 3646 11048 3710
rect 11112 3646 11129 3710
rect 11193 3646 11210 3710
rect 11274 3646 11291 3710
rect 11355 3646 11372 3710
rect 11436 3646 11453 3710
rect 11517 3646 11534 3710
rect 11598 3646 11615 3710
rect 11679 3646 11696 3710
rect 11760 3646 11777 3710
rect 11841 3646 11858 3710
rect 11922 3646 11939 3710
rect 12003 3646 12020 3710
rect 12084 3646 12101 3710
rect 12165 3646 12182 3710
rect 12246 3646 12263 3710
rect 12327 3646 12344 3710
rect 12408 3646 12425 3710
rect 12489 3646 12506 3710
rect 12570 3646 12587 3710
rect 12651 3646 12668 3710
rect 12732 3646 12749 3710
rect 12813 3646 12830 3710
rect 12894 3646 12911 3710
rect 12975 3646 12992 3710
rect 13056 3646 13073 3710
rect 13137 3646 13154 3710
rect 13218 3646 13235 3710
rect 13299 3646 13316 3710
rect 13380 3646 13397 3710
rect 13461 3646 13478 3710
rect 13542 3646 13559 3710
rect 13623 3646 13640 3710
rect 13704 3646 13721 3710
rect 13785 3646 13802 3710
rect 13866 3646 13883 3710
rect 13947 3646 13964 3710
rect 14028 3646 14045 3710
rect 14109 3646 14126 3710
rect 14190 3646 14207 3710
rect 14271 3646 14288 3710
rect 14352 3646 14369 3710
rect 14433 3646 14451 3710
rect 14515 3646 14533 3710
rect 14597 3646 14615 3710
rect 14679 3646 14697 3710
rect 14761 3646 14779 3710
rect 14843 3646 14861 3710
rect 14925 3646 14931 3710
rect 10151 3624 14931 3646
rect 10151 3560 10157 3624
rect 10221 3560 10238 3624
rect 10302 3560 10319 3624
rect 10383 3560 10400 3624
rect 10464 3560 10481 3624
rect 10545 3560 10562 3624
rect 10626 3560 10643 3624
rect 10707 3560 10724 3624
rect 10788 3560 10805 3624
rect 10869 3560 10886 3624
rect 10950 3560 10967 3624
rect 11031 3560 11048 3624
rect 11112 3560 11129 3624
rect 11193 3560 11210 3624
rect 11274 3560 11291 3624
rect 11355 3560 11372 3624
rect 11436 3560 11453 3624
rect 11517 3560 11534 3624
rect 11598 3560 11615 3624
rect 11679 3560 11696 3624
rect 11760 3560 11777 3624
rect 11841 3560 11858 3624
rect 11922 3560 11939 3624
rect 12003 3560 12020 3624
rect 12084 3560 12101 3624
rect 12165 3560 12182 3624
rect 12246 3560 12263 3624
rect 12327 3560 12344 3624
rect 12408 3560 12425 3624
rect 12489 3560 12506 3624
rect 12570 3560 12587 3624
rect 12651 3560 12668 3624
rect 12732 3560 12749 3624
rect 12813 3560 12830 3624
rect 12894 3560 12911 3624
rect 12975 3560 12992 3624
rect 13056 3560 13073 3624
rect 13137 3560 13154 3624
rect 13218 3560 13235 3624
rect 13299 3560 13316 3624
rect 13380 3560 13397 3624
rect 13461 3560 13478 3624
rect 13542 3560 13559 3624
rect 13623 3560 13640 3624
rect 13704 3560 13721 3624
rect 13785 3560 13802 3624
rect 13866 3560 13883 3624
rect 13947 3560 13964 3624
rect 14028 3560 14045 3624
rect 14109 3560 14126 3624
rect 14190 3560 14207 3624
rect 14271 3560 14288 3624
rect 14352 3560 14369 3624
rect 14433 3560 14451 3624
rect 14515 3560 14533 3624
rect 14597 3560 14615 3624
rect 14679 3560 14697 3624
rect 14761 3560 14779 3624
rect 14843 3560 14861 3624
rect 14925 3560 14931 3624
rect 10151 3558 14931 3560
<< via3 >>
rect 135 18527 199 18591
rect 217 18527 281 18591
rect 299 18527 363 18591
rect 381 18527 445 18591
rect 463 18527 527 18591
rect 545 18527 609 18591
rect 627 18527 691 18591
rect 709 18527 773 18591
rect 791 18527 855 18591
rect 873 18527 937 18591
rect 955 18527 1019 18591
rect 1037 18527 1101 18591
rect 1119 18527 1183 18591
rect 1201 18527 1265 18591
rect 1283 18527 1347 18591
rect 1365 18527 1429 18591
rect 1447 18527 1511 18591
rect 1529 18527 1593 18591
rect 1611 18527 1675 18591
rect 1693 18527 1757 18591
rect 1775 18527 1839 18591
rect 1857 18527 1921 18591
rect 1939 18527 2003 18591
rect 2021 18527 2085 18591
rect 2103 18527 2167 18591
rect 2185 18527 2249 18591
rect 2267 18527 2331 18591
rect 2349 18527 2413 18591
rect 2431 18527 2495 18591
rect 2513 18527 2577 18591
rect 2594 18527 2658 18591
rect 2675 18527 2739 18591
rect 2756 18527 2820 18591
rect 135 18445 199 18509
rect 217 18445 281 18509
rect 299 18445 363 18509
rect 381 18445 445 18509
rect 463 18445 527 18509
rect 545 18445 609 18509
rect 627 18445 691 18509
rect 709 18445 773 18509
rect 791 18445 855 18509
rect 873 18445 937 18509
rect 955 18445 1019 18509
rect 1037 18445 1101 18509
rect 1119 18445 1183 18509
rect 1201 18445 1265 18509
rect 1283 18445 1347 18509
rect 1365 18445 1429 18509
rect 1447 18445 1511 18509
rect 1529 18445 1593 18509
rect 1611 18445 1675 18509
rect 1693 18445 1757 18509
rect 1775 18445 1839 18509
rect 1857 18445 1921 18509
rect 1939 18445 2003 18509
rect 2021 18445 2085 18509
rect 2103 18445 2167 18509
rect 2185 18445 2249 18509
rect 2267 18445 2331 18509
rect 2349 18445 2413 18509
rect 2431 18445 2495 18509
rect 2513 18445 2577 18509
rect 2594 18445 2658 18509
rect 2675 18445 2739 18509
rect 2756 18445 2820 18509
rect 135 18363 199 18427
rect 217 18363 281 18427
rect 299 18363 363 18427
rect 381 18363 445 18427
rect 463 18363 527 18427
rect 545 18363 609 18427
rect 627 18363 691 18427
rect 709 18363 773 18427
rect 791 18363 855 18427
rect 873 18363 937 18427
rect 955 18363 1019 18427
rect 1037 18363 1101 18427
rect 1119 18363 1183 18427
rect 1201 18363 1265 18427
rect 1283 18363 1347 18427
rect 1365 18363 1429 18427
rect 1447 18363 1511 18427
rect 1529 18363 1593 18427
rect 1611 18363 1675 18427
rect 1693 18363 1757 18427
rect 1775 18363 1839 18427
rect 1857 18363 1921 18427
rect 1939 18363 2003 18427
rect 2021 18363 2085 18427
rect 2103 18363 2167 18427
rect 2185 18363 2249 18427
rect 2267 18363 2331 18427
rect 2349 18363 2413 18427
rect 2431 18363 2495 18427
rect 2513 18363 2577 18427
rect 2594 18363 2658 18427
rect 2675 18363 2739 18427
rect 2756 18363 2820 18427
rect 12231 18527 12295 18591
rect 12312 18527 12376 18591
rect 12393 18527 12457 18591
rect 12474 18527 12538 18591
rect 12556 18527 12620 18591
rect 12638 18527 12702 18591
rect 12720 18527 12784 18591
rect 12802 18527 12866 18591
rect 12884 18527 12948 18591
rect 12966 18527 13030 18591
rect 13048 18527 13112 18591
rect 13130 18527 13194 18591
rect 13212 18527 13276 18591
rect 13294 18527 13358 18591
rect 13376 18527 13440 18591
rect 13458 18527 13522 18591
rect 13540 18527 13604 18591
rect 13622 18527 13686 18591
rect 13704 18527 13768 18591
rect 13786 18527 13850 18591
rect 13868 18527 13932 18591
rect 13950 18527 14014 18591
rect 14032 18527 14096 18591
rect 14114 18527 14178 18591
rect 14196 18527 14260 18591
rect 14278 18527 14342 18591
rect 14360 18527 14424 18591
rect 14442 18527 14506 18591
rect 14524 18527 14588 18591
rect 14606 18527 14670 18591
rect 14688 18527 14752 18591
rect 14770 18527 14834 18591
rect 14852 18527 14916 18591
rect 12231 18445 12295 18509
rect 12312 18445 12376 18509
rect 12393 18445 12457 18509
rect 12474 18445 12538 18509
rect 12556 18445 12620 18509
rect 12638 18445 12702 18509
rect 12720 18445 12784 18509
rect 12802 18445 12866 18509
rect 12884 18445 12948 18509
rect 12966 18445 13030 18509
rect 13048 18445 13112 18509
rect 13130 18445 13194 18509
rect 13212 18445 13276 18509
rect 13294 18445 13358 18509
rect 13376 18445 13440 18509
rect 13458 18445 13522 18509
rect 13540 18445 13604 18509
rect 13622 18445 13686 18509
rect 13704 18445 13768 18509
rect 13786 18445 13850 18509
rect 13868 18445 13932 18509
rect 13950 18445 14014 18509
rect 14032 18445 14096 18509
rect 14114 18445 14178 18509
rect 14196 18445 14260 18509
rect 14278 18445 14342 18509
rect 14360 18445 14424 18509
rect 14442 18445 14506 18509
rect 14524 18445 14588 18509
rect 14606 18445 14670 18509
rect 14688 18445 14752 18509
rect 14770 18445 14834 18509
rect 14852 18445 14916 18509
rect 12231 18363 12295 18427
rect 12312 18363 12376 18427
rect 12393 18363 12457 18427
rect 12474 18363 12538 18427
rect 12556 18363 12620 18427
rect 12638 18363 12702 18427
rect 12720 18363 12784 18427
rect 12802 18363 12866 18427
rect 12884 18363 12948 18427
rect 12966 18363 13030 18427
rect 13048 18363 13112 18427
rect 13130 18363 13194 18427
rect 13212 18363 13276 18427
rect 13294 18363 13358 18427
rect 13376 18363 13440 18427
rect 13458 18363 13522 18427
rect 13540 18363 13604 18427
rect 13622 18363 13686 18427
rect 13704 18363 13768 18427
rect 13786 18363 13850 18427
rect 13868 18363 13932 18427
rect 13950 18363 14014 18427
rect 14032 18363 14096 18427
rect 14114 18363 14178 18427
rect 14196 18363 14260 18427
rect 14278 18363 14342 18427
rect 14360 18363 14424 18427
rect 14442 18363 14506 18427
rect 14524 18363 14588 18427
rect 14606 18363 14670 18427
rect 14688 18363 14752 18427
rect 14770 18363 14834 18427
rect 14852 18363 14916 18427
rect 135 18281 199 18345
rect 217 18281 281 18345
rect 299 18281 363 18345
rect 381 18281 445 18345
rect 463 18281 527 18345
rect 545 18281 609 18345
rect 627 18281 691 18345
rect 709 18281 773 18345
rect 791 18281 855 18345
rect 873 18281 937 18345
rect 955 18281 1019 18345
rect 1037 18281 1101 18345
rect 1119 18281 1183 18345
rect 1201 18281 1265 18345
rect 1283 18281 1347 18345
rect 1365 18281 1429 18345
rect 1447 18281 1511 18345
rect 1529 18281 1593 18345
rect 1611 18281 1675 18345
rect 1693 18281 1757 18345
rect 1775 18281 1839 18345
rect 1857 18281 1921 18345
rect 1939 18281 2003 18345
rect 2021 18281 2085 18345
rect 2103 18281 2167 18345
rect 2185 18281 2249 18345
rect 2267 18281 2331 18345
rect 2349 18281 2413 18345
rect 2431 18281 2495 18345
rect 2513 18281 2577 18345
rect 2594 18281 2658 18345
rect 2675 18281 2739 18345
rect 2756 18281 2820 18345
rect 2852 18277 2916 18341
rect 3008 18277 3072 18341
rect 135 18199 199 18263
rect 217 18199 281 18263
rect 299 18199 363 18263
rect 381 18199 445 18263
rect 463 18199 527 18263
rect 545 18199 609 18263
rect 627 18199 691 18263
rect 709 18199 773 18263
rect 791 18199 855 18263
rect 873 18199 937 18263
rect 955 18199 1019 18263
rect 1037 18199 1101 18263
rect 1119 18199 1183 18263
rect 1201 18199 1265 18263
rect 1283 18199 1347 18263
rect 1365 18199 1429 18263
rect 1447 18199 1511 18263
rect 1529 18199 1593 18263
rect 1611 18199 1675 18263
rect 1693 18199 1757 18263
rect 1775 18199 1839 18263
rect 1857 18199 1921 18263
rect 1939 18199 2003 18263
rect 2021 18199 2085 18263
rect 2103 18199 2167 18263
rect 2185 18199 2249 18263
rect 2267 18199 2331 18263
rect 2349 18199 2413 18263
rect 2431 18199 2495 18263
rect 2513 18199 2577 18263
rect 2594 18199 2658 18263
rect 2675 18199 2739 18263
rect 2756 18199 2820 18263
rect 2852 18191 2916 18255
rect 3008 18191 3072 18255
rect 11979 18277 12043 18341
rect 12135 18277 12199 18341
rect 12231 18281 12295 18345
rect 12312 18281 12376 18345
rect 12393 18281 12457 18345
rect 12474 18281 12538 18345
rect 12556 18281 12620 18345
rect 12638 18281 12702 18345
rect 12720 18281 12784 18345
rect 12802 18281 12866 18345
rect 12884 18281 12948 18345
rect 12966 18281 13030 18345
rect 13048 18281 13112 18345
rect 13130 18281 13194 18345
rect 13212 18281 13276 18345
rect 13294 18281 13358 18345
rect 13376 18281 13440 18345
rect 13458 18281 13522 18345
rect 13540 18281 13604 18345
rect 13622 18281 13686 18345
rect 13704 18281 13768 18345
rect 13786 18281 13850 18345
rect 13868 18281 13932 18345
rect 13950 18281 14014 18345
rect 14032 18281 14096 18345
rect 14114 18281 14178 18345
rect 14196 18281 14260 18345
rect 14278 18281 14342 18345
rect 14360 18281 14424 18345
rect 14442 18281 14506 18345
rect 14524 18281 14588 18345
rect 14606 18281 14670 18345
rect 14688 18281 14752 18345
rect 14770 18281 14834 18345
rect 14852 18281 14916 18345
rect 11979 18191 12043 18255
rect 12135 18191 12199 18255
rect 12231 18199 12295 18263
rect 12312 18199 12376 18263
rect 12393 18199 12457 18263
rect 12474 18199 12538 18263
rect 12556 18199 12620 18263
rect 12638 18199 12702 18263
rect 12720 18199 12784 18263
rect 12802 18199 12866 18263
rect 12884 18199 12948 18263
rect 12966 18199 13030 18263
rect 13048 18199 13112 18263
rect 13130 18199 13194 18263
rect 13212 18199 13276 18263
rect 13294 18199 13358 18263
rect 13376 18199 13440 18263
rect 13458 18199 13522 18263
rect 13540 18199 13604 18263
rect 13622 18199 13686 18263
rect 13704 18199 13768 18263
rect 13786 18199 13850 18263
rect 13868 18199 13932 18263
rect 13950 18199 14014 18263
rect 14032 18199 14096 18263
rect 14114 18199 14178 18263
rect 14196 18199 14260 18263
rect 14278 18199 14342 18263
rect 14360 18199 14424 18263
rect 14442 18199 14506 18263
rect 14524 18199 14588 18263
rect 14606 18199 14670 18263
rect 14688 18199 14752 18263
rect 14770 18199 14834 18263
rect 14852 18199 14916 18263
rect 135 18117 199 18181
rect 217 18117 281 18181
rect 299 18117 363 18181
rect 381 18117 445 18181
rect 463 18117 527 18181
rect 545 18117 609 18181
rect 627 18117 691 18181
rect 709 18117 773 18181
rect 791 18117 855 18181
rect 873 18117 937 18181
rect 955 18117 1019 18181
rect 1037 18117 1101 18181
rect 1119 18117 1183 18181
rect 1201 18117 1265 18181
rect 1283 18117 1347 18181
rect 1365 18117 1429 18181
rect 1447 18117 1511 18181
rect 1529 18117 1593 18181
rect 1611 18117 1675 18181
rect 1693 18117 1757 18181
rect 1775 18117 1839 18181
rect 1857 18117 1921 18181
rect 1939 18117 2003 18181
rect 2021 18117 2085 18181
rect 2103 18117 2167 18181
rect 2185 18117 2249 18181
rect 2267 18117 2331 18181
rect 2349 18117 2413 18181
rect 2431 18117 2495 18181
rect 2513 18117 2577 18181
rect 2594 18117 2658 18181
rect 2675 18117 2739 18181
rect 2756 18117 2820 18181
rect 2856 18099 2920 18163
rect 2938 18099 3002 18163
rect 3020 18099 3084 18163
rect 3102 18099 3166 18163
rect 3184 18099 3248 18163
rect 135 18035 199 18099
rect 217 18035 281 18099
rect 299 18035 363 18099
rect 381 18035 445 18099
rect 463 18035 527 18099
rect 545 18035 609 18099
rect 627 18035 691 18099
rect 709 18035 773 18099
rect 791 18035 855 18099
rect 873 18035 937 18099
rect 955 18035 1019 18099
rect 1037 18035 1101 18099
rect 1119 18035 1183 18099
rect 1201 18035 1265 18099
rect 1283 18035 1347 18099
rect 1365 18035 1429 18099
rect 1447 18035 1511 18099
rect 1529 18035 1593 18099
rect 1611 18035 1675 18099
rect 1693 18035 1757 18099
rect 1775 18035 1839 18099
rect 1857 18035 1921 18099
rect 1939 18035 2003 18099
rect 2021 18035 2085 18099
rect 2103 18035 2167 18099
rect 2185 18035 2249 18099
rect 2267 18035 2331 18099
rect 2349 18035 2413 18099
rect 2431 18035 2495 18099
rect 2513 18035 2577 18099
rect 2594 18035 2658 18099
rect 2675 18035 2739 18099
rect 2756 18035 2820 18099
rect 135 17953 199 18017
rect 217 17953 281 18017
rect 299 17953 363 18017
rect 381 17953 445 18017
rect 463 17953 527 18017
rect 545 17953 609 18017
rect 627 17953 691 18017
rect 709 17953 773 18017
rect 791 17953 855 18017
rect 873 17953 937 18017
rect 955 17953 1019 18017
rect 1037 17953 1101 18017
rect 1119 17953 1183 18017
rect 1201 17953 1265 18017
rect 1283 17953 1347 18017
rect 1365 17953 1429 18017
rect 1447 17953 1511 18017
rect 1529 17953 1593 18017
rect 1611 17953 1675 18017
rect 1693 17953 1757 18017
rect 1775 17953 1839 18017
rect 1857 17953 1921 18017
rect 1939 17953 2003 18017
rect 2021 17953 2085 18017
rect 2103 17953 2167 18017
rect 2185 17953 2249 18017
rect 2267 17953 2331 18017
rect 2349 17953 2413 18017
rect 2431 17953 2495 18017
rect 2513 17953 2577 18017
rect 2594 17953 2658 18017
rect 2675 17953 2739 18017
rect 2756 17953 2820 18017
rect 2856 18013 2920 18077
rect 2938 18013 3002 18077
rect 3020 18013 3084 18077
rect 3102 18013 3166 18077
rect 3184 18013 3248 18077
rect 135 17871 199 17935
rect 217 17871 281 17935
rect 299 17871 363 17935
rect 381 17871 445 17935
rect 463 17871 527 17935
rect 545 17871 609 17935
rect 627 17871 691 17935
rect 709 17871 773 17935
rect 791 17871 855 17935
rect 873 17871 937 17935
rect 955 17871 1019 17935
rect 1037 17871 1101 17935
rect 1119 17871 1183 17935
rect 1201 17871 1265 17935
rect 1283 17871 1347 17935
rect 1365 17871 1429 17935
rect 1447 17871 1511 17935
rect 1529 17871 1593 17935
rect 1611 17871 1675 17935
rect 1693 17871 1757 17935
rect 1775 17871 1839 17935
rect 1857 17871 1921 17935
rect 1939 17871 2003 17935
rect 2021 17871 2085 17935
rect 2103 17871 2167 17935
rect 2185 17871 2249 17935
rect 2267 17871 2331 17935
rect 2349 17871 2413 17935
rect 2431 17871 2495 17935
rect 2513 17871 2577 17935
rect 2594 17871 2658 17935
rect 2675 17871 2739 17935
rect 2756 17871 2820 17935
rect 2856 17927 2920 17991
rect 2938 17927 3002 17991
rect 3020 17927 3084 17991
rect 3102 17927 3166 17991
rect 3184 17927 3248 17991
rect 11803 18099 11867 18163
rect 11885 18099 11949 18163
rect 11967 18099 12031 18163
rect 12049 18099 12113 18163
rect 12131 18099 12195 18163
rect 12231 18117 12295 18181
rect 12312 18117 12376 18181
rect 12393 18117 12457 18181
rect 12474 18117 12538 18181
rect 12556 18117 12620 18181
rect 12638 18117 12702 18181
rect 12720 18117 12784 18181
rect 12802 18117 12866 18181
rect 12884 18117 12948 18181
rect 12966 18117 13030 18181
rect 13048 18117 13112 18181
rect 13130 18117 13194 18181
rect 13212 18117 13276 18181
rect 13294 18117 13358 18181
rect 13376 18117 13440 18181
rect 13458 18117 13522 18181
rect 13540 18117 13604 18181
rect 13622 18117 13686 18181
rect 13704 18117 13768 18181
rect 13786 18117 13850 18181
rect 13868 18117 13932 18181
rect 13950 18117 14014 18181
rect 14032 18117 14096 18181
rect 14114 18117 14178 18181
rect 14196 18117 14260 18181
rect 14278 18117 14342 18181
rect 14360 18117 14424 18181
rect 14442 18117 14506 18181
rect 14524 18117 14588 18181
rect 14606 18117 14670 18181
rect 14688 18117 14752 18181
rect 14770 18117 14834 18181
rect 14852 18117 14916 18181
rect 11803 18013 11867 18077
rect 11885 18013 11949 18077
rect 11967 18013 12031 18077
rect 12049 18013 12113 18077
rect 12131 18013 12195 18077
rect 12231 18035 12295 18099
rect 12312 18035 12376 18099
rect 12393 18035 12457 18099
rect 12474 18035 12538 18099
rect 12556 18035 12620 18099
rect 12638 18035 12702 18099
rect 12720 18035 12784 18099
rect 12802 18035 12866 18099
rect 12884 18035 12948 18099
rect 12966 18035 13030 18099
rect 13048 18035 13112 18099
rect 13130 18035 13194 18099
rect 13212 18035 13276 18099
rect 13294 18035 13358 18099
rect 13376 18035 13440 18099
rect 13458 18035 13522 18099
rect 13540 18035 13604 18099
rect 13622 18035 13686 18099
rect 13704 18035 13768 18099
rect 13786 18035 13850 18099
rect 13868 18035 13932 18099
rect 13950 18035 14014 18099
rect 14032 18035 14096 18099
rect 14114 18035 14178 18099
rect 14196 18035 14260 18099
rect 14278 18035 14342 18099
rect 14360 18035 14424 18099
rect 14442 18035 14506 18099
rect 14524 18035 14588 18099
rect 14606 18035 14670 18099
rect 14688 18035 14752 18099
rect 14770 18035 14834 18099
rect 14852 18035 14916 18099
rect 11803 17927 11867 17991
rect 11885 17927 11949 17991
rect 11967 17927 12031 17991
rect 12049 17927 12113 17991
rect 12131 17927 12195 17991
rect 12231 17953 12295 18017
rect 12312 17953 12376 18017
rect 12393 17953 12457 18017
rect 12474 17953 12538 18017
rect 12556 17953 12620 18017
rect 12638 17953 12702 18017
rect 12720 17953 12784 18017
rect 12802 17953 12866 18017
rect 12884 17953 12948 18017
rect 12966 17953 13030 18017
rect 13048 17953 13112 18017
rect 13130 17953 13194 18017
rect 13212 17953 13276 18017
rect 13294 17953 13358 18017
rect 13376 17953 13440 18017
rect 13458 17953 13522 18017
rect 13540 17953 13604 18017
rect 13622 17953 13686 18017
rect 13704 17953 13768 18017
rect 13786 17953 13850 18017
rect 13868 17953 13932 18017
rect 13950 17953 14014 18017
rect 14032 17953 14096 18017
rect 14114 17953 14178 18017
rect 14196 17953 14260 18017
rect 14278 17953 14342 18017
rect 14360 17953 14424 18017
rect 14442 17953 14506 18017
rect 14524 17953 14588 18017
rect 14606 17953 14670 18017
rect 14688 17953 14752 18017
rect 14770 17953 14834 18017
rect 14852 17953 14916 18017
rect 135 17789 199 17853
rect 217 17789 281 17853
rect 299 17789 363 17853
rect 381 17789 445 17853
rect 463 17789 527 17853
rect 545 17789 609 17853
rect 627 17789 691 17853
rect 709 17789 773 17853
rect 791 17789 855 17853
rect 873 17789 937 17853
rect 955 17789 1019 17853
rect 1037 17789 1101 17853
rect 1119 17789 1183 17853
rect 1201 17789 1265 17853
rect 1283 17789 1347 17853
rect 1365 17789 1429 17853
rect 1447 17789 1511 17853
rect 1529 17789 1593 17853
rect 1611 17789 1675 17853
rect 1693 17789 1757 17853
rect 1775 17789 1839 17853
rect 1857 17789 1921 17853
rect 1939 17789 2003 17853
rect 2021 17789 2085 17853
rect 2103 17789 2167 17853
rect 2185 17789 2249 17853
rect 2267 17789 2331 17853
rect 2349 17789 2413 17853
rect 2431 17789 2495 17853
rect 2513 17789 2577 17853
rect 2594 17789 2658 17853
rect 2675 17789 2739 17853
rect 2756 17789 2820 17853
rect 2856 17841 2920 17905
rect 2938 17841 3002 17905
rect 3020 17841 3084 17905
rect 3102 17841 3166 17905
rect 3184 17841 3248 17905
rect 3284 17841 3348 17905
rect 3440 17841 3504 17905
rect 135 17707 199 17771
rect 217 17707 281 17771
rect 299 17707 363 17771
rect 381 17707 445 17771
rect 463 17707 527 17771
rect 545 17707 609 17771
rect 627 17707 691 17771
rect 709 17707 773 17771
rect 791 17707 855 17771
rect 873 17707 937 17771
rect 955 17707 1019 17771
rect 1037 17707 1101 17771
rect 1119 17707 1183 17771
rect 1201 17707 1265 17771
rect 1283 17707 1347 17771
rect 1365 17707 1429 17771
rect 1447 17707 1511 17771
rect 1529 17707 1593 17771
rect 1611 17707 1675 17771
rect 1693 17707 1757 17771
rect 1775 17707 1839 17771
rect 1857 17707 1921 17771
rect 1939 17707 2003 17771
rect 2021 17707 2085 17771
rect 2103 17707 2167 17771
rect 2185 17707 2249 17771
rect 2267 17707 2331 17771
rect 2349 17707 2413 17771
rect 2431 17707 2495 17771
rect 2513 17707 2577 17771
rect 2594 17707 2658 17771
rect 2675 17707 2739 17771
rect 2756 17707 2820 17771
rect 2856 17755 2920 17819
rect 2938 17755 3002 17819
rect 3020 17755 3084 17819
rect 3102 17755 3166 17819
rect 3184 17755 3248 17819
rect 3284 17757 3348 17821
rect 3440 17757 3504 17821
rect 135 17625 199 17689
rect 217 17625 281 17689
rect 299 17625 363 17689
rect 381 17625 445 17689
rect 463 17625 527 17689
rect 545 17625 609 17689
rect 627 17625 691 17689
rect 709 17625 773 17689
rect 791 17625 855 17689
rect 873 17625 937 17689
rect 955 17625 1019 17689
rect 1037 17625 1101 17689
rect 1119 17625 1183 17689
rect 1201 17625 1265 17689
rect 1283 17625 1347 17689
rect 1365 17625 1429 17689
rect 1447 17625 1511 17689
rect 1529 17625 1593 17689
rect 1611 17625 1675 17689
rect 1693 17625 1757 17689
rect 1775 17625 1839 17689
rect 1857 17625 1921 17689
rect 1939 17625 2003 17689
rect 2021 17625 2085 17689
rect 2103 17625 2167 17689
rect 2185 17625 2249 17689
rect 2267 17625 2331 17689
rect 2349 17625 2413 17689
rect 2431 17625 2495 17689
rect 2513 17625 2577 17689
rect 2594 17625 2658 17689
rect 2675 17625 2739 17689
rect 2756 17625 2820 17689
rect 2856 17670 2920 17734
rect 2938 17670 3002 17734
rect 3020 17670 3084 17734
rect 3102 17670 3166 17734
rect 3184 17670 3248 17734
rect 3284 17674 3348 17738
rect 3440 17674 3504 17738
rect 11547 17841 11611 17905
rect 11703 17841 11767 17905
rect 11803 17841 11867 17905
rect 11885 17841 11949 17905
rect 11967 17841 12031 17905
rect 12049 17841 12113 17905
rect 12131 17841 12195 17905
rect 12231 17871 12295 17935
rect 12312 17871 12376 17935
rect 12393 17871 12457 17935
rect 12474 17871 12538 17935
rect 12556 17871 12620 17935
rect 12638 17871 12702 17935
rect 12720 17871 12784 17935
rect 12802 17871 12866 17935
rect 12884 17871 12948 17935
rect 12966 17871 13030 17935
rect 13048 17871 13112 17935
rect 13130 17871 13194 17935
rect 13212 17871 13276 17935
rect 13294 17871 13358 17935
rect 13376 17871 13440 17935
rect 13458 17871 13522 17935
rect 13540 17871 13604 17935
rect 13622 17871 13686 17935
rect 13704 17871 13768 17935
rect 13786 17871 13850 17935
rect 13868 17871 13932 17935
rect 13950 17871 14014 17935
rect 14032 17871 14096 17935
rect 14114 17871 14178 17935
rect 14196 17871 14260 17935
rect 14278 17871 14342 17935
rect 14360 17871 14424 17935
rect 14442 17871 14506 17935
rect 14524 17871 14588 17935
rect 14606 17871 14670 17935
rect 14688 17871 14752 17935
rect 14770 17871 14834 17935
rect 14852 17871 14916 17935
rect 11547 17757 11611 17821
rect 11703 17757 11767 17821
rect 11803 17755 11867 17819
rect 11885 17755 11949 17819
rect 11967 17755 12031 17819
rect 12049 17755 12113 17819
rect 12131 17755 12195 17819
rect 12231 17789 12295 17853
rect 12312 17789 12376 17853
rect 12393 17789 12457 17853
rect 12474 17789 12538 17853
rect 12556 17789 12620 17853
rect 12638 17789 12702 17853
rect 12720 17789 12784 17853
rect 12802 17789 12866 17853
rect 12884 17789 12948 17853
rect 12966 17789 13030 17853
rect 13048 17789 13112 17853
rect 13130 17789 13194 17853
rect 13212 17789 13276 17853
rect 13294 17789 13358 17853
rect 13376 17789 13440 17853
rect 13458 17789 13522 17853
rect 13540 17789 13604 17853
rect 13622 17789 13686 17853
rect 13704 17789 13768 17853
rect 13786 17789 13850 17853
rect 13868 17789 13932 17853
rect 13950 17789 14014 17853
rect 14032 17789 14096 17853
rect 14114 17789 14178 17853
rect 14196 17789 14260 17853
rect 14278 17789 14342 17853
rect 14360 17789 14424 17853
rect 14442 17789 14506 17853
rect 14524 17789 14588 17853
rect 14606 17789 14670 17853
rect 14688 17789 14752 17853
rect 14770 17789 14834 17853
rect 14852 17789 14916 17853
rect 11547 17674 11611 17738
rect 11703 17674 11767 17738
rect 11803 17670 11867 17734
rect 11885 17670 11949 17734
rect 11967 17670 12031 17734
rect 12049 17670 12113 17734
rect 12131 17670 12195 17734
rect 12231 17707 12295 17771
rect 12312 17707 12376 17771
rect 12393 17707 12457 17771
rect 12474 17707 12538 17771
rect 12556 17707 12620 17771
rect 12638 17707 12702 17771
rect 12720 17707 12784 17771
rect 12802 17707 12866 17771
rect 12884 17707 12948 17771
rect 12966 17707 13030 17771
rect 13048 17707 13112 17771
rect 13130 17707 13194 17771
rect 13212 17707 13276 17771
rect 13294 17707 13358 17771
rect 13376 17707 13440 17771
rect 13458 17707 13522 17771
rect 13540 17707 13604 17771
rect 13622 17707 13686 17771
rect 13704 17707 13768 17771
rect 13786 17707 13850 17771
rect 13868 17707 13932 17771
rect 13950 17707 14014 17771
rect 14032 17707 14096 17771
rect 14114 17707 14178 17771
rect 14196 17707 14260 17771
rect 14278 17707 14342 17771
rect 14360 17707 14424 17771
rect 14442 17707 14506 17771
rect 14524 17707 14588 17771
rect 14606 17707 14670 17771
rect 14688 17707 14752 17771
rect 14770 17707 14834 17771
rect 14852 17707 14916 17771
rect 135 17543 199 17607
rect 217 17543 281 17607
rect 299 17543 363 17607
rect 381 17543 445 17607
rect 463 17543 527 17607
rect 545 17543 609 17607
rect 627 17543 691 17607
rect 709 17543 773 17607
rect 791 17543 855 17607
rect 873 17543 937 17607
rect 955 17543 1019 17607
rect 1037 17543 1101 17607
rect 1119 17543 1183 17607
rect 1201 17543 1265 17607
rect 1283 17543 1347 17607
rect 1365 17543 1429 17607
rect 1447 17543 1511 17607
rect 1529 17543 1593 17607
rect 1611 17543 1675 17607
rect 1693 17543 1757 17607
rect 1775 17543 1839 17607
rect 1857 17543 1921 17607
rect 1939 17543 2003 17607
rect 2021 17543 2085 17607
rect 2103 17543 2167 17607
rect 2185 17543 2249 17607
rect 2267 17543 2331 17607
rect 2349 17543 2413 17607
rect 2431 17543 2495 17607
rect 2513 17543 2577 17607
rect 2594 17543 2658 17607
rect 2675 17543 2739 17607
rect 2756 17543 2820 17607
rect 2881 17563 2945 17627
rect 2963 17563 3027 17627
rect 3045 17563 3109 17627
rect 3127 17563 3191 17627
rect 3209 17563 3273 17627
rect 3291 17563 3355 17627
rect 3373 17563 3437 17627
rect 3455 17563 3519 17627
rect 3537 17563 3601 17627
rect 3619 17563 3683 17627
rect 3701 17563 3765 17627
rect 135 17461 199 17525
rect 217 17461 281 17525
rect 299 17461 363 17525
rect 381 17461 445 17525
rect 463 17461 527 17525
rect 545 17461 609 17525
rect 627 17461 691 17525
rect 709 17461 773 17525
rect 791 17461 855 17525
rect 873 17461 937 17525
rect 955 17461 1019 17525
rect 1037 17461 1101 17525
rect 1119 17461 1183 17525
rect 1201 17461 1265 17525
rect 1283 17461 1347 17525
rect 1365 17461 1429 17525
rect 1447 17461 1511 17525
rect 1529 17461 1593 17525
rect 1611 17461 1675 17525
rect 1693 17461 1757 17525
rect 1775 17461 1839 17525
rect 1857 17461 1921 17525
rect 1939 17461 2003 17525
rect 2021 17461 2085 17525
rect 2103 17461 2167 17525
rect 2185 17461 2249 17525
rect 2267 17461 2331 17525
rect 2349 17461 2413 17525
rect 2431 17461 2495 17525
rect 2513 17461 2577 17525
rect 2594 17461 2658 17525
rect 2675 17461 2739 17525
rect 2756 17461 2820 17525
rect 2881 17482 2945 17546
rect 2963 17482 3027 17546
rect 3045 17482 3109 17546
rect 3127 17482 3191 17546
rect 3209 17482 3273 17546
rect 3291 17482 3355 17546
rect 3373 17482 3437 17546
rect 3455 17482 3519 17546
rect 3537 17482 3601 17546
rect 3619 17482 3683 17546
rect 3701 17482 3765 17546
rect 135 17379 199 17443
rect 217 17379 281 17443
rect 299 17379 363 17443
rect 381 17379 445 17443
rect 463 17379 527 17443
rect 545 17379 609 17443
rect 627 17379 691 17443
rect 709 17379 773 17443
rect 791 17379 855 17443
rect 873 17379 937 17443
rect 955 17379 1019 17443
rect 1037 17379 1101 17443
rect 1119 17379 1183 17443
rect 1201 17379 1265 17443
rect 1283 17379 1347 17443
rect 1365 17379 1429 17443
rect 1447 17379 1511 17443
rect 1529 17379 1593 17443
rect 1611 17379 1675 17443
rect 1693 17379 1757 17443
rect 1775 17379 1839 17443
rect 1857 17379 1921 17443
rect 1939 17379 2003 17443
rect 2021 17379 2085 17443
rect 2103 17379 2167 17443
rect 2185 17379 2249 17443
rect 2267 17379 2331 17443
rect 2349 17379 2413 17443
rect 2431 17379 2495 17443
rect 2513 17379 2577 17443
rect 2594 17379 2658 17443
rect 2675 17379 2739 17443
rect 2756 17379 2820 17443
rect 2881 17401 2945 17465
rect 2963 17401 3027 17465
rect 3045 17401 3109 17465
rect 3127 17401 3191 17465
rect 3209 17401 3273 17465
rect 3291 17401 3355 17465
rect 3373 17401 3437 17465
rect 3455 17401 3519 17465
rect 3537 17401 3601 17465
rect 3619 17401 3683 17465
rect 3701 17401 3765 17465
rect 11286 17563 11350 17627
rect 11368 17563 11432 17627
rect 11450 17563 11514 17627
rect 11532 17563 11596 17627
rect 11614 17563 11678 17627
rect 11696 17563 11760 17627
rect 11778 17563 11842 17627
rect 11860 17563 11924 17627
rect 11942 17563 12006 17627
rect 12024 17563 12088 17627
rect 12106 17563 12170 17627
rect 12231 17625 12295 17689
rect 12312 17625 12376 17689
rect 12393 17625 12457 17689
rect 12474 17625 12538 17689
rect 12556 17625 12620 17689
rect 12638 17625 12702 17689
rect 12720 17625 12784 17689
rect 12802 17625 12866 17689
rect 12884 17625 12948 17689
rect 12966 17625 13030 17689
rect 13048 17625 13112 17689
rect 13130 17625 13194 17689
rect 13212 17625 13276 17689
rect 13294 17625 13358 17689
rect 13376 17625 13440 17689
rect 13458 17625 13522 17689
rect 13540 17625 13604 17689
rect 13622 17625 13686 17689
rect 13704 17625 13768 17689
rect 13786 17625 13850 17689
rect 13868 17625 13932 17689
rect 13950 17625 14014 17689
rect 14032 17625 14096 17689
rect 14114 17625 14178 17689
rect 14196 17625 14260 17689
rect 14278 17625 14342 17689
rect 14360 17625 14424 17689
rect 14442 17625 14506 17689
rect 14524 17625 14588 17689
rect 14606 17625 14670 17689
rect 14688 17625 14752 17689
rect 14770 17625 14834 17689
rect 14852 17625 14916 17689
rect 11286 17482 11350 17546
rect 11368 17482 11432 17546
rect 11450 17482 11514 17546
rect 11532 17482 11596 17546
rect 11614 17482 11678 17546
rect 11696 17482 11760 17546
rect 11778 17482 11842 17546
rect 11860 17482 11924 17546
rect 11942 17482 12006 17546
rect 12024 17482 12088 17546
rect 12106 17482 12170 17546
rect 12231 17543 12295 17607
rect 12312 17543 12376 17607
rect 12393 17543 12457 17607
rect 12474 17543 12538 17607
rect 12556 17543 12620 17607
rect 12638 17543 12702 17607
rect 12720 17543 12784 17607
rect 12802 17543 12866 17607
rect 12884 17543 12948 17607
rect 12966 17543 13030 17607
rect 13048 17543 13112 17607
rect 13130 17543 13194 17607
rect 13212 17543 13276 17607
rect 13294 17543 13358 17607
rect 13376 17543 13440 17607
rect 13458 17543 13522 17607
rect 13540 17543 13604 17607
rect 13622 17543 13686 17607
rect 13704 17543 13768 17607
rect 13786 17543 13850 17607
rect 13868 17543 13932 17607
rect 13950 17543 14014 17607
rect 14032 17543 14096 17607
rect 14114 17543 14178 17607
rect 14196 17543 14260 17607
rect 14278 17543 14342 17607
rect 14360 17543 14424 17607
rect 14442 17543 14506 17607
rect 14524 17543 14588 17607
rect 14606 17543 14670 17607
rect 14688 17543 14752 17607
rect 14770 17543 14834 17607
rect 14852 17543 14916 17607
rect 135 17297 199 17361
rect 217 17297 281 17361
rect 299 17297 363 17361
rect 381 17297 445 17361
rect 463 17297 527 17361
rect 545 17297 609 17361
rect 627 17297 691 17361
rect 709 17297 773 17361
rect 791 17297 855 17361
rect 873 17297 937 17361
rect 955 17297 1019 17361
rect 1037 17297 1101 17361
rect 1119 17297 1183 17361
rect 1201 17297 1265 17361
rect 1283 17297 1347 17361
rect 1365 17297 1429 17361
rect 1447 17297 1511 17361
rect 1529 17297 1593 17361
rect 1611 17297 1675 17361
rect 1693 17297 1757 17361
rect 1775 17297 1839 17361
rect 1857 17297 1921 17361
rect 1939 17297 2003 17361
rect 2021 17297 2085 17361
rect 2103 17297 2167 17361
rect 2185 17297 2249 17361
rect 2267 17297 2331 17361
rect 2349 17297 2413 17361
rect 2431 17297 2495 17361
rect 2513 17297 2577 17361
rect 2594 17297 2658 17361
rect 2675 17297 2739 17361
rect 2756 17297 2820 17361
rect 2881 17320 2945 17384
rect 2963 17320 3027 17384
rect 3045 17320 3109 17384
rect 3127 17320 3191 17384
rect 3209 17320 3273 17384
rect 3291 17320 3355 17384
rect 3373 17320 3437 17384
rect 3455 17320 3519 17384
rect 3537 17320 3601 17384
rect 3619 17320 3683 17384
rect 3701 17320 3765 17384
rect 3800 17338 3864 17402
rect 3948 17338 4012 17402
rect 135 17215 199 17279
rect 217 17215 281 17279
rect 299 17215 363 17279
rect 381 17215 445 17279
rect 463 17215 527 17279
rect 545 17215 609 17279
rect 627 17215 691 17279
rect 709 17215 773 17279
rect 791 17215 855 17279
rect 873 17215 937 17279
rect 955 17215 1019 17279
rect 1037 17215 1101 17279
rect 1119 17215 1183 17279
rect 1201 17215 1265 17279
rect 1283 17215 1347 17279
rect 1365 17215 1429 17279
rect 1447 17215 1511 17279
rect 1529 17215 1593 17279
rect 1611 17215 1675 17279
rect 1693 17215 1757 17279
rect 1775 17215 1839 17279
rect 1857 17215 1921 17279
rect 1939 17215 2003 17279
rect 2021 17215 2085 17279
rect 2103 17215 2167 17279
rect 2185 17215 2249 17279
rect 2267 17215 2331 17279
rect 2349 17215 2413 17279
rect 2431 17215 2495 17279
rect 2513 17215 2577 17279
rect 2594 17215 2658 17279
rect 2675 17215 2739 17279
rect 2756 17215 2820 17279
rect 2881 17239 2945 17303
rect 2963 17239 3027 17303
rect 3045 17239 3109 17303
rect 3127 17239 3191 17303
rect 3209 17239 3273 17303
rect 3291 17239 3355 17303
rect 3373 17239 3437 17303
rect 3455 17239 3519 17303
rect 3537 17239 3601 17303
rect 3619 17239 3683 17303
rect 3701 17239 3765 17303
rect 3800 17250 3864 17314
rect 3948 17250 4012 17314
rect 135 17133 199 17197
rect 217 17133 281 17197
rect 299 17133 363 17197
rect 381 17133 445 17197
rect 463 17133 527 17197
rect 545 17133 609 17197
rect 627 17133 691 17197
rect 709 17133 773 17197
rect 791 17133 855 17197
rect 873 17133 937 17197
rect 955 17133 1019 17197
rect 1037 17133 1101 17197
rect 1119 17133 1183 17197
rect 1201 17133 1265 17197
rect 1283 17133 1347 17197
rect 1365 17133 1429 17197
rect 1447 17133 1511 17197
rect 1529 17133 1593 17197
rect 1611 17133 1675 17197
rect 1693 17133 1757 17197
rect 1775 17133 1839 17197
rect 1857 17133 1921 17197
rect 1939 17133 2003 17197
rect 2021 17133 2085 17197
rect 2103 17133 2167 17197
rect 2185 17133 2249 17197
rect 2267 17133 2331 17197
rect 2349 17133 2413 17197
rect 2431 17133 2495 17197
rect 2513 17133 2577 17197
rect 2594 17133 2658 17197
rect 2675 17133 2739 17197
rect 2756 17133 2820 17197
rect 2881 17159 2945 17223
rect 2963 17159 3027 17223
rect 3045 17159 3109 17223
rect 3127 17159 3191 17223
rect 3209 17159 3273 17223
rect 3291 17159 3355 17223
rect 3373 17159 3437 17223
rect 3455 17159 3519 17223
rect 3537 17159 3601 17223
rect 3619 17159 3683 17223
rect 3701 17159 3765 17223
rect 3800 17163 3864 17227
rect 3948 17163 4012 17227
rect 11039 17338 11103 17402
rect 11187 17338 11251 17402
rect 11286 17401 11350 17465
rect 11368 17401 11432 17465
rect 11450 17401 11514 17465
rect 11532 17401 11596 17465
rect 11614 17401 11678 17465
rect 11696 17401 11760 17465
rect 11778 17401 11842 17465
rect 11860 17401 11924 17465
rect 11942 17401 12006 17465
rect 12024 17401 12088 17465
rect 12106 17401 12170 17465
rect 12231 17461 12295 17525
rect 12312 17461 12376 17525
rect 12393 17461 12457 17525
rect 12474 17461 12538 17525
rect 12556 17461 12620 17525
rect 12638 17461 12702 17525
rect 12720 17461 12784 17525
rect 12802 17461 12866 17525
rect 12884 17461 12948 17525
rect 12966 17461 13030 17525
rect 13048 17461 13112 17525
rect 13130 17461 13194 17525
rect 13212 17461 13276 17525
rect 13294 17461 13358 17525
rect 13376 17461 13440 17525
rect 13458 17461 13522 17525
rect 13540 17461 13604 17525
rect 13622 17461 13686 17525
rect 13704 17461 13768 17525
rect 13786 17461 13850 17525
rect 13868 17461 13932 17525
rect 13950 17461 14014 17525
rect 14032 17461 14096 17525
rect 14114 17461 14178 17525
rect 14196 17461 14260 17525
rect 14278 17461 14342 17525
rect 14360 17461 14424 17525
rect 14442 17461 14506 17525
rect 14524 17461 14588 17525
rect 14606 17461 14670 17525
rect 14688 17461 14752 17525
rect 14770 17461 14834 17525
rect 14852 17461 14916 17525
rect 11286 17320 11350 17384
rect 11368 17320 11432 17384
rect 11450 17320 11514 17384
rect 11532 17320 11596 17384
rect 11614 17320 11678 17384
rect 11696 17320 11760 17384
rect 11778 17320 11842 17384
rect 11860 17320 11924 17384
rect 11942 17320 12006 17384
rect 12024 17320 12088 17384
rect 12106 17320 12170 17384
rect 12231 17379 12295 17443
rect 12312 17379 12376 17443
rect 12393 17379 12457 17443
rect 12474 17379 12538 17443
rect 12556 17379 12620 17443
rect 12638 17379 12702 17443
rect 12720 17379 12784 17443
rect 12802 17379 12866 17443
rect 12884 17379 12948 17443
rect 12966 17379 13030 17443
rect 13048 17379 13112 17443
rect 13130 17379 13194 17443
rect 13212 17379 13276 17443
rect 13294 17379 13358 17443
rect 13376 17379 13440 17443
rect 13458 17379 13522 17443
rect 13540 17379 13604 17443
rect 13622 17379 13686 17443
rect 13704 17379 13768 17443
rect 13786 17379 13850 17443
rect 13868 17379 13932 17443
rect 13950 17379 14014 17443
rect 14032 17379 14096 17443
rect 14114 17379 14178 17443
rect 14196 17379 14260 17443
rect 14278 17379 14342 17443
rect 14360 17379 14424 17443
rect 14442 17379 14506 17443
rect 14524 17379 14588 17443
rect 14606 17379 14670 17443
rect 14688 17379 14752 17443
rect 14770 17379 14834 17443
rect 14852 17379 14916 17443
rect 11039 17250 11103 17314
rect 11187 17250 11251 17314
rect 11286 17239 11350 17303
rect 11368 17239 11432 17303
rect 11450 17239 11514 17303
rect 11532 17239 11596 17303
rect 11614 17239 11678 17303
rect 11696 17239 11760 17303
rect 11778 17239 11842 17303
rect 11860 17239 11924 17303
rect 11942 17239 12006 17303
rect 12024 17239 12088 17303
rect 12106 17239 12170 17303
rect 12231 17297 12295 17361
rect 12312 17297 12376 17361
rect 12393 17297 12457 17361
rect 12474 17297 12538 17361
rect 12556 17297 12620 17361
rect 12638 17297 12702 17361
rect 12720 17297 12784 17361
rect 12802 17297 12866 17361
rect 12884 17297 12948 17361
rect 12966 17297 13030 17361
rect 13048 17297 13112 17361
rect 13130 17297 13194 17361
rect 13212 17297 13276 17361
rect 13294 17297 13358 17361
rect 13376 17297 13440 17361
rect 13458 17297 13522 17361
rect 13540 17297 13604 17361
rect 13622 17297 13686 17361
rect 13704 17297 13768 17361
rect 13786 17297 13850 17361
rect 13868 17297 13932 17361
rect 13950 17297 14014 17361
rect 14032 17297 14096 17361
rect 14114 17297 14178 17361
rect 14196 17297 14260 17361
rect 14278 17297 14342 17361
rect 14360 17297 14424 17361
rect 14442 17297 14506 17361
rect 14524 17297 14588 17361
rect 14606 17297 14670 17361
rect 14688 17297 14752 17361
rect 14770 17297 14834 17361
rect 14852 17297 14916 17361
rect 11039 17163 11103 17227
rect 11187 17163 11251 17227
rect 11286 17159 11350 17223
rect 11368 17159 11432 17223
rect 11450 17159 11514 17223
rect 11532 17159 11596 17223
rect 11614 17159 11678 17223
rect 11696 17159 11760 17223
rect 11778 17159 11842 17223
rect 11860 17159 11924 17223
rect 11942 17159 12006 17223
rect 12024 17159 12088 17223
rect 12106 17159 12170 17223
rect 12231 17215 12295 17279
rect 12312 17215 12376 17279
rect 12393 17215 12457 17279
rect 12474 17215 12538 17279
rect 12556 17215 12620 17279
rect 12638 17215 12702 17279
rect 12720 17215 12784 17279
rect 12802 17215 12866 17279
rect 12884 17215 12948 17279
rect 12966 17215 13030 17279
rect 13048 17215 13112 17279
rect 13130 17215 13194 17279
rect 13212 17215 13276 17279
rect 13294 17215 13358 17279
rect 13376 17215 13440 17279
rect 13458 17215 13522 17279
rect 13540 17215 13604 17279
rect 13622 17215 13686 17279
rect 13704 17215 13768 17279
rect 13786 17215 13850 17279
rect 13868 17215 13932 17279
rect 13950 17215 14014 17279
rect 14032 17215 14096 17279
rect 14114 17215 14178 17279
rect 14196 17215 14260 17279
rect 14278 17215 14342 17279
rect 14360 17215 14424 17279
rect 14442 17215 14506 17279
rect 14524 17215 14588 17279
rect 14606 17215 14670 17279
rect 14688 17215 14752 17279
rect 14770 17215 14834 17279
rect 14852 17215 14916 17279
rect 135 17051 199 17115
rect 217 17051 281 17115
rect 299 17051 363 17115
rect 381 17051 445 17115
rect 463 17051 527 17115
rect 545 17051 609 17115
rect 627 17051 691 17115
rect 709 17051 773 17115
rect 791 17051 855 17115
rect 873 17051 937 17115
rect 955 17051 1019 17115
rect 1037 17051 1101 17115
rect 1119 17051 1183 17115
rect 1201 17051 1265 17115
rect 1283 17051 1347 17115
rect 1365 17051 1429 17115
rect 1447 17051 1511 17115
rect 1529 17051 1593 17115
rect 1611 17051 1675 17115
rect 1693 17051 1757 17115
rect 1775 17051 1839 17115
rect 1857 17051 1921 17115
rect 1939 17051 2003 17115
rect 2021 17051 2085 17115
rect 2103 17051 2167 17115
rect 2185 17051 2249 17115
rect 2267 17051 2331 17115
rect 2349 17051 2413 17115
rect 2431 17051 2495 17115
rect 2513 17051 2577 17115
rect 2594 17051 2658 17115
rect 2675 17051 2739 17115
rect 2756 17051 2820 17115
rect 2881 17079 2945 17143
rect 2963 17079 3027 17143
rect 3045 17079 3109 17143
rect 3127 17079 3191 17143
rect 3209 17079 3273 17143
rect 3291 17079 3355 17143
rect 3373 17079 3437 17143
rect 3455 17079 3519 17143
rect 3537 17079 3601 17143
rect 3619 17079 3683 17143
rect 3701 17079 3765 17143
rect 135 16969 199 17033
rect 217 16969 281 17033
rect 299 16969 363 17033
rect 381 16969 445 17033
rect 463 16969 527 17033
rect 545 16969 609 17033
rect 627 16969 691 17033
rect 709 16969 773 17033
rect 791 16969 855 17033
rect 873 16969 937 17033
rect 955 16969 1019 17033
rect 1037 16969 1101 17033
rect 1119 16969 1183 17033
rect 1201 16969 1265 17033
rect 1283 16969 1347 17033
rect 1365 16969 1429 17033
rect 1447 16969 1511 17033
rect 1529 16969 1593 17033
rect 1611 16969 1675 17033
rect 1693 16969 1757 17033
rect 1775 16969 1839 17033
rect 1857 16969 1921 17033
rect 1939 16969 2003 17033
rect 2021 16969 2085 17033
rect 2103 16969 2167 17033
rect 2185 16969 2249 17033
rect 2267 16969 2331 17033
rect 2349 16969 2413 17033
rect 2431 16969 2495 17033
rect 2513 16969 2577 17033
rect 2594 16969 2658 17033
rect 2675 16969 2739 17033
rect 2756 16969 2820 17033
rect 2881 16999 2945 17063
rect 2963 16999 3027 17063
rect 3045 16999 3109 17063
rect 3127 16999 3191 17063
rect 3209 16999 3273 17063
rect 3291 16999 3355 17063
rect 3373 16999 3437 17063
rect 3455 16999 3519 17063
rect 3537 16999 3601 17063
rect 3619 16999 3683 17063
rect 3701 16999 3765 17063
rect 3838 17053 3902 17117
rect 3934 17053 3998 17117
rect 4030 17053 4094 17117
rect 4126 17053 4190 17117
rect 4222 17053 4286 17117
rect 135 16887 199 16951
rect 217 16887 281 16951
rect 299 16887 363 16951
rect 381 16887 445 16951
rect 463 16887 527 16951
rect 545 16887 609 16951
rect 627 16887 691 16951
rect 709 16887 773 16951
rect 791 16887 855 16951
rect 873 16887 937 16951
rect 955 16887 1019 16951
rect 1037 16887 1101 16951
rect 1119 16887 1183 16951
rect 1201 16887 1265 16951
rect 1283 16887 1347 16951
rect 1365 16887 1429 16951
rect 1447 16887 1511 16951
rect 1529 16887 1593 16951
rect 1611 16887 1675 16951
rect 1693 16887 1757 16951
rect 1775 16887 1839 16951
rect 1857 16887 1921 16951
rect 1939 16887 2003 16951
rect 2021 16887 2085 16951
rect 2103 16887 2167 16951
rect 2185 16887 2249 16951
rect 2267 16887 2331 16951
rect 2349 16887 2413 16951
rect 2431 16887 2495 16951
rect 2513 16887 2577 16951
rect 2594 16887 2658 16951
rect 2675 16887 2739 16951
rect 2756 16887 2820 16951
rect 2881 16919 2945 16983
rect 2963 16919 3027 16983
rect 3045 16919 3109 16983
rect 3127 16919 3191 16983
rect 3209 16919 3273 16983
rect 3291 16919 3355 16983
rect 3373 16919 3437 16983
rect 3455 16919 3519 16983
rect 3537 16919 3601 16983
rect 3619 16919 3683 16983
rect 3701 16919 3765 16983
rect 3838 16960 3902 17024
rect 3934 16960 3998 17024
rect 4030 16960 4094 17024
rect 4126 16960 4190 17024
rect 4222 16960 4286 17024
rect 135 16805 199 16869
rect 217 16805 281 16869
rect 299 16805 363 16869
rect 381 16805 445 16869
rect 463 16805 527 16869
rect 545 16805 609 16869
rect 627 16805 691 16869
rect 709 16805 773 16869
rect 791 16805 855 16869
rect 873 16805 937 16869
rect 955 16805 1019 16869
rect 1037 16805 1101 16869
rect 1119 16805 1183 16869
rect 1201 16805 1265 16869
rect 1283 16805 1347 16869
rect 1365 16805 1429 16869
rect 1447 16805 1511 16869
rect 1529 16805 1593 16869
rect 1611 16805 1675 16869
rect 1693 16805 1757 16869
rect 1775 16805 1839 16869
rect 1857 16805 1921 16869
rect 1939 16805 2003 16869
rect 2021 16805 2085 16869
rect 2103 16805 2167 16869
rect 2185 16805 2249 16869
rect 2267 16805 2331 16869
rect 2349 16805 2413 16869
rect 2431 16805 2495 16869
rect 2513 16805 2577 16869
rect 2594 16805 2658 16869
rect 2675 16805 2739 16869
rect 2756 16805 2820 16869
rect 2881 16839 2945 16903
rect 2963 16839 3027 16903
rect 3045 16839 3109 16903
rect 3127 16839 3191 16903
rect 3209 16839 3273 16903
rect 3291 16839 3355 16903
rect 3373 16839 3437 16903
rect 3455 16839 3519 16903
rect 3537 16839 3601 16903
rect 3619 16839 3683 16903
rect 3701 16839 3765 16903
rect 3838 16867 3902 16931
rect 3934 16867 3998 16931
rect 4030 16867 4094 16931
rect 4126 16867 4190 16931
rect 4222 16867 4286 16931
rect 10765 17053 10829 17117
rect 10861 17053 10925 17117
rect 10957 17053 11021 17117
rect 11053 17053 11117 17117
rect 11149 17053 11213 17117
rect 11286 17079 11350 17143
rect 11368 17079 11432 17143
rect 11450 17079 11514 17143
rect 11532 17079 11596 17143
rect 11614 17079 11678 17143
rect 11696 17079 11760 17143
rect 11778 17079 11842 17143
rect 11860 17079 11924 17143
rect 11942 17079 12006 17143
rect 12024 17079 12088 17143
rect 12106 17079 12170 17143
rect 12231 17133 12295 17197
rect 12312 17133 12376 17197
rect 12393 17133 12457 17197
rect 12474 17133 12538 17197
rect 12556 17133 12620 17197
rect 12638 17133 12702 17197
rect 12720 17133 12784 17197
rect 12802 17133 12866 17197
rect 12884 17133 12948 17197
rect 12966 17133 13030 17197
rect 13048 17133 13112 17197
rect 13130 17133 13194 17197
rect 13212 17133 13276 17197
rect 13294 17133 13358 17197
rect 13376 17133 13440 17197
rect 13458 17133 13522 17197
rect 13540 17133 13604 17197
rect 13622 17133 13686 17197
rect 13704 17133 13768 17197
rect 13786 17133 13850 17197
rect 13868 17133 13932 17197
rect 13950 17133 14014 17197
rect 14032 17133 14096 17197
rect 14114 17133 14178 17197
rect 14196 17133 14260 17197
rect 14278 17133 14342 17197
rect 14360 17133 14424 17197
rect 14442 17133 14506 17197
rect 14524 17133 14588 17197
rect 14606 17133 14670 17197
rect 14688 17133 14752 17197
rect 14770 17133 14834 17197
rect 14852 17133 14916 17197
rect 10765 16960 10829 17024
rect 10861 16960 10925 17024
rect 10957 16960 11021 17024
rect 11053 16960 11117 17024
rect 11149 16960 11213 17024
rect 11286 16999 11350 17063
rect 11368 16999 11432 17063
rect 11450 16999 11514 17063
rect 11532 16999 11596 17063
rect 11614 16999 11678 17063
rect 11696 16999 11760 17063
rect 11778 16999 11842 17063
rect 11860 16999 11924 17063
rect 11942 16999 12006 17063
rect 12024 16999 12088 17063
rect 12106 16999 12170 17063
rect 12231 17051 12295 17115
rect 12312 17051 12376 17115
rect 12393 17051 12457 17115
rect 12474 17051 12538 17115
rect 12556 17051 12620 17115
rect 12638 17051 12702 17115
rect 12720 17051 12784 17115
rect 12802 17051 12866 17115
rect 12884 17051 12948 17115
rect 12966 17051 13030 17115
rect 13048 17051 13112 17115
rect 13130 17051 13194 17115
rect 13212 17051 13276 17115
rect 13294 17051 13358 17115
rect 13376 17051 13440 17115
rect 13458 17051 13522 17115
rect 13540 17051 13604 17115
rect 13622 17051 13686 17115
rect 13704 17051 13768 17115
rect 13786 17051 13850 17115
rect 13868 17051 13932 17115
rect 13950 17051 14014 17115
rect 14032 17051 14096 17115
rect 14114 17051 14178 17115
rect 14196 17051 14260 17115
rect 14278 17051 14342 17115
rect 14360 17051 14424 17115
rect 14442 17051 14506 17115
rect 14524 17051 14588 17115
rect 14606 17051 14670 17115
rect 14688 17051 14752 17115
rect 14770 17051 14834 17115
rect 14852 17051 14916 17115
rect 10765 16867 10829 16931
rect 10861 16867 10925 16931
rect 10957 16867 11021 16931
rect 11053 16867 11117 16931
rect 11149 16867 11213 16931
rect 11286 16919 11350 16983
rect 11368 16919 11432 16983
rect 11450 16919 11514 16983
rect 11532 16919 11596 16983
rect 11614 16919 11678 16983
rect 11696 16919 11760 16983
rect 11778 16919 11842 16983
rect 11860 16919 11924 16983
rect 11942 16919 12006 16983
rect 12024 16919 12088 16983
rect 12106 16919 12170 16983
rect 12231 16969 12295 17033
rect 12312 16969 12376 17033
rect 12393 16969 12457 17033
rect 12474 16969 12538 17033
rect 12556 16969 12620 17033
rect 12638 16969 12702 17033
rect 12720 16969 12784 17033
rect 12802 16969 12866 17033
rect 12884 16969 12948 17033
rect 12966 16969 13030 17033
rect 13048 16969 13112 17033
rect 13130 16969 13194 17033
rect 13212 16969 13276 17033
rect 13294 16969 13358 17033
rect 13376 16969 13440 17033
rect 13458 16969 13522 17033
rect 13540 16969 13604 17033
rect 13622 16969 13686 17033
rect 13704 16969 13768 17033
rect 13786 16969 13850 17033
rect 13868 16969 13932 17033
rect 13950 16969 14014 17033
rect 14032 16969 14096 17033
rect 14114 16969 14178 17033
rect 14196 16969 14260 17033
rect 14278 16969 14342 17033
rect 14360 16969 14424 17033
rect 14442 16969 14506 17033
rect 14524 16969 14588 17033
rect 14606 16969 14670 17033
rect 14688 16969 14752 17033
rect 14770 16969 14834 17033
rect 14852 16969 14916 17033
rect 135 16723 199 16787
rect 217 16723 281 16787
rect 299 16723 363 16787
rect 381 16723 445 16787
rect 463 16723 527 16787
rect 545 16723 609 16787
rect 627 16723 691 16787
rect 709 16723 773 16787
rect 791 16723 855 16787
rect 873 16723 937 16787
rect 955 16723 1019 16787
rect 1037 16723 1101 16787
rect 1119 16723 1183 16787
rect 1201 16723 1265 16787
rect 1283 16723 1347 16787
rect 1365 16723 1429 16787
rect 1447 16723 1511 16787
rect 1529 16723 1593 16787
rect 1611 16723 1675 16787
rect 1693 16723 1757 16787
rect 1775 16723 1839 16787
rect 1857 16723 1921 16787
rect 1939 16723 2003 16787
rect 2021 16723 2085 16787
rect 2103 16723 2167 16787
rect 2185 16723 2249 16787
rect 2267 16723 2331 16787
rect 2349 16723 2413 16787
rect 2431 16723 2495 16787
rect 2513 16723 2577 16787
rect 2594 16723 2658 16787
rect 2675 16723 2739 16787
rect 2756 16723 2820 16787
rect 2881 16759 2945 16823
rect 2963 16759 3027 16823
rect 3045 16759 3109 16823
rect 3127 16759 3191 16823
rect 3209 16759 3273 16823
rect 3291 16759 3355 16823
rect 3373 16759 3437 16823
rect 3455 16759 3519 16823
rect 3537 16759 3601 16823
rect 3619 16759 3683 16823
rect 3701 16759 3765 16823
rect 3838 16774 3902 16838
rect 3934 16774 3998 16838
rect 4030 16774 4094 16838
rect 4126 16774 4190 16838
rect 4222 16774 4286 16838
rect 4331 16792 4395 16856
rect 4489 16792 4553 16856
rect 135 16641 199 16705
rect 217 16641 281 16705
rect 299 16641 363 16705
rect 381 16641 445 16705
rect 463 16641 527 16705
rect 545 16641 609 16705
rect 627 16641 691 16705
rect 709 16641 773 16705
rect 791 16641 855 16705
rect 873 16641 937 16705
rect 955 16641 1019 16705
rect 1037 16641 1101 16705
rect 1119 16641 1183 16705
rect 1201 16641 1265 16705
rect 1283 16641 1347 16705
rect 1365 16641 1429 16705
rect 1447 16641 1511 16705
rect 1529 16641 1593 16705
rect 1611 16641 1675 16705
rect 1693 16641 1757 16705
rect 1775 16641 1839 16705
rect 1857 16641 1921 16705
rect 1939 16641 2003 16705
rect 2021 16641 2085 16705
rect 2103 16641 2167 16705
rect 2185 16641 2249 16705
rect 2267 16641 2331 16705
rect 2349 16641 2413 16705
rect 2431 16641 2495 16705
rect 2513 16641 2577 16705
rect 2594 16641 2658 16705
rect 2675 16641 2739 16705
rect 2756 16641 2820 16705
rect 2881 16679 2945 16743
rect 2963 16679 3027 16743
rect 3045 16679 3109 16743
rect 3127 16679 3191 16743
rect 3209 16679 3273 16743
rect 3291 16679 3355 16743
rect 3373 16679 3437 16743
rect 3455 16679 3519 16743
rect 3537 16679 3601 16743
rect 3619 16679 3683 16743
rect 3701 16679 3765 16743
rect 3838 16682 3902 16746
rect 3934 16682 3998 16746
rect 4030 16682 4094 16746
rect 4126 16682 4190 16746
rect 4222 16682 4286 16746
rect 4331 16682 4395 16746
rect 4489 16682 4553 16746
rect 135 16559 199 16623
rect 217 16559 281 16623
rect 299 16559 363 16623
rect 381 16559 445 16623
rect 463 16559 527 16623
rect 545 16559 609 16623
rect 627 16559 691 16623
rect 709 16559 773 16623
rect 791 16559 855 16623
rect 873 16559 937 16623
rect 955 16559 1019 16623
rect 1037 16559 1101 16623
rect 1119 16559 1183 16623
rect 1201 16559 1265 16623
rect 1283 16559 1347 16623
rect 1365 16559 1429 16623
rect 1447 16559 1511 16623
rect 1529 16559 1593 16623
rect 1611 16559 1675 16623
rect 1693 16559 1757 16623
rect 1775 16559 1839 16623
rect 1857 16559 1921 16623
rect 1939 16559 2003 16623
rect 2021 16559 2085 16623
rect 2103 16559 2167 16623
rect 2185 16559 2249 16623
rect 2267 16559 2331 16623
rect 2349 16559 2413 16623
rect 2431 16559 2495 16623
rect 2513 16559 2577 16623
rect 2594 16559 2658 16623
rect 2675 16559 2739 16623
rect 2756 16559 2820 16623
rect 2881 16599 2945 16663
rect 2963 16599 3027 16663
rect 3045 16599 3109 16663
rect 3127 16599 3191 16663
rect 3209 16599 3273 16663
rect 3291 16599 3355 16663
rect 3373 16599 3437 16663
rect 3455 16599 3519 16663
rect 3537 16599 3601 16663
rect 3619 16599 3683 16663
rect 3701 16599 3765 16663
rect 3838 16590 3902 16654
rect 3934 16590 3998 16654
rect 4030 16590 4094 16654
rect 4126 16590 4190 16654
rect 4222 16590 4286 16654
rect 4331 16572 4395 16636
rect 4489 16572 4553 16636
rect 10498 16792 10562 16856
rect 10656 16792 10720 16856
rect 11286 16839 11350 16903
rect 11368 16839 11432 16903
rect 11450 16839 11514 16903
rect 11532 16839 11596 16903
rect 11614 16839 11678 16903
rect 11696 16839 11760 16903
rect 11778 16839 11842 16903
rect 11860 16839 11924 16903
rect 11942 16839 12006 16903
rect 12024 16839 12088 16903
rect 12106 16839 12170 16903
rect 12231 16887 12295 16951
rect 12312 16887 12376 16951
rect 12393 16887 12457 16951
rect 12474 16887 12538 16951
rect 12556 16887 12620 16951
rect 12638 16887 12702 16951
rect 12720 16887 12784 16951
rect 12802 16887 12866 16951
rect 12884 16887 12948 16951
rect 12966 16887 13030 16951
rect 13048 16887 13112 16951
rect 13130 16887 13194 16951
rect 13212 16887 13276 16951
rect 13294 16887 13358 16951
rect 13376 16887 13440 16951
rect 13458 16887 13522 16951
rect 13540 16887 13604 16951
rect 13622 16887 13686 16951
rect 13704 16887 13768 16951
rect 13786 16887 13850 16951
rect 13868 16887 13932 16951
rect 13950 16887 14014 16951
rect 14032 16887 14096 16951
rect 14114 16887 14178 16951
rect 14196 16887 14260 16951
rect 14278 16887 14342 16951
rect 14360 16887 14424 16951
rect 14442 16887 14506 16951
rect 14524 16887 14588 16951
rect 14606 16887 14670 16951
rect 14688 16887 14752 16951
rect 14770 16887 14834 16951
rect 14852 16887 14916 16951
rect 10765 16774 10829 16838
rect 10861 16774 10925 16838
rect 10957 16774 11021 16838
rect 11053 16774 11117 16838
rect 11149 16774 11213 16838
rect 11286 16759 11350 16823
rect 11368 16759 11432 16823
rect 11450 16759 11514 16823
rect 11532 16759 11596 16823
rect 11614 16759 11678 16823
rect 11696 16759 11760 16823
rect 11778 16759 11842 16823
rect 11860 16759 11924 16823
rect 11942 16759 12006 16823
rect 12024 16759 12088 16823
rect 12106 16759 12170 16823
rect 12231 16805 12295 16869
rect 12312 16805 12376 16869
rect 12393 16805 12457 16869
rect 12474 16805 12538 16869
rect 12556 16805 12620 16869
rect 12638 16805 12702 16869
rect 12720 16805 12784 16869
rect 12802 16805 12866 16869
rect 12884 16805 12948 16869
rect 12966 16805 13030 16869
rect 13048 16805 13112 16869
rect 13130 16805 13194 16869
rect 13212 16805 13276 16869
rect 13294 16805 13358 16869
rect 13376 16805 13440 16869
rect 13458 16805 13522 16869
rect 13540 16805 13604 16869
rect 13622 16805 13686 16869
rect 13704 16805 13768 16869
rect 13786 16805 13850 16869
rect 13868 16805 13932 16869
rect 13950 16805 14014 16869
rect 14032 16805 14096 16869
rect 14114 16805 14178 16869
rect 14196 16805 14260 16869
rect 14278 16805 14342 16869
rect 14360 16805 14424 16869
rect 14442 16805 14506 16869
rect 14524 16805 14588 16869
rect 14606 16805 14670 16869
rect 14688 16805 14752 16869
rect 14770 16805 14834 16869
rect 14852 16805 14916 16869
rect 10498 16682 10562 16746
rect 10656 16682 10720 16746
rect 10765 16682 10829 16746
rect 10861 16682 10925 16746
rect 10957 16682 11021 16746
rect 11053 16682 11117 16746
rect 11149 16682 11213 16746
rect 11286 16679 11350 16743
rect 11368 16679 11432 16743
rect 11450 16679 11514 16743
rect 11532 16679 11596 16743
rect 11614 16679 11678 16743
rect 11696 16679 11760 16743
rect 11778 16679 11842 16743
rect 11860 16679 11924 16743
rect 11942 16679 12006 16743
rect 12024 16679 12088 16743
rect 12106 16679 12170 16743
rect 12231 16723 12295 16787
rect 12312 16723 12376 16787
rect 12393 16723 12457 16787
rect 12474 16723 12538 16787
rect 12556 16723 12620 16787
rect 12638 16723 12702 16787
rect 12720 16723 12784 16787
rect 12802 16723 12866 16787
rect 12884 16723 12948 16787
rect 12966 16723 13030 16787
rect 13048 16723 13112 16787
rect 13130 16723 13194 16787
rect 13212 16723 13276 16787
rect 13294 16723 13358 16787
rect 13376 16723 13440 16787
rect 13458 16723 13522 16787
rect 13540 16723 13604 16787
rect 13622 16723 13686 16787
rect 13704 16723 13768 16787
rect 13786 16723 13850 16787
rect 13868 16723 13932 16787
rect 13950 16723 14014 16787
rect 14032 16723 14096 16787
rect 14114 16723 14178 16787
rect 14196 16723 14260 16787
rect 14278 16723 14342 16787
rect 14360 16723 14424 16787
rect 14442 16723 14506 16787
rect 14524 16723 14588 16787
rect 14606 16723 14670 16787
rect 14688 16723 14752 16787
rect 14770 16723 14834 16787
rect 14852 16723 14916 16787
rect 10498 16572 10562 16636
rect 10656 16572 10720 16636
rect 10765 16590 10829 16654
rect 10861 16590 10925 16654
rect 10957 16590 11021 16654
rect 11053 16590 11117 16654
rect 11149 16590 11213 16654
rect 11286 16599 11350 16663
rect 11368 16599 11432 16663
rect 11450 16599 11514 16663
rect 11532 16599 11596 16663
rect 11614 16599 11678 16663
rect 11696 16599 11760 16663
rect 11778 16599 11842 16663
rect 11860 16599 11924 16663
rect 11942 16599 12006 16663
rect 12024 16599 12088 16663
rect 12106 16599 12170 16663
rect 12231 16641 12295 16705
rect 12312 16641 12376 16705
rect 12393 16641 12457 16705
rect 12474 16641 12538 16705
rect 12556 16641 12620 16705
rect 12638 16641 12702 16705
rect 12720 16641 12784 16705
rect 12802 16641 12866 16705
rect 12884 16641 12948 16705
rect 12966 16641 13030 16705
rect 13048 16641 13112 16705
rect 13130 16641 13194 16705
rect 13212 16641 13276 16705
rect 13294 16641 13358 16705
rect 13376 16641 13440 16705
rect 13458 16641 13522 16705
rect 13540 16641 13604 16705
rect 13622 16641 13686 16705
rect 13704 16641 13768 16705
rect 13786 16641 13850 16705
rect 13868 16641 13932 16705
rect 13950 16641 14014 16705
rect 14032 16641 14096 16705
rect 14114 16641 14178 16705
rect 14196 16641 14260 16705
rect 14278 16641 14342 16705
rect 14360 16641 14424 16705
rect 14442 16641 14506 16705
rect 14524 16641 14588 16705
rect 14606 16641 14670 16705
rect 14688 16641 14752 16705
rect 14770 16641 14834 16705
rect 14852 16641 14916 16705
rect 12231 16559 12295 16623
rect 12312 16559 12376 16623
rect 12393 16559 12457 16623
rect 12474 16559 12538 16623
rect 12556 16559 12620 16623
rect 12638 16559 12702 16623
rect 12720 16559 12784 16623
rect 12802 16559 12866 16623
rect 12884 16559 12948 16623
rect 12966 16559 13030 16623
rect 13048 16559 13112 16623
rect 13130 16559 13194 16623
rect 13212 16559 13276 16623
rect 13294 16559 13358 16623
rect 13376 16559 13440 16623
rect 13458 16559 13522 16623
rect 13540 16559 13604 16623
rect 13622 16559 13686 16623
rect 13704 16559 13768 16623
rect 13786 16559 13850 16623
rect 13868 16559 13932 16623
rect 13950 16559 14014 16623
rect 14032 16559 14096 16623
rect 14114 16559 14178 16623
rect 14196 16559 14260 16623
rect 14278 16559 14342 16623
rect 14360 16559 14424 16623
rect 14442 16559 14506 16623
rect 14524 16559 14588 16623
rect 14606 16559 14670 16623
rect 14688 16559 14752 16623
rect 14770 16559 14834 16623
rect 14852 16559 14916 16623
rect 157 16460 221 16524
rect 237 16460 301 16524
rect 317 16460 381 16524
rect 397 16460 461 16524
rect 477 16460 541 16524
rect 557 16460 621 16524
rect 637 16460 701 16524
rect 717 16460 781 16524
rect 797 16460 861 16524
rect 877 16460 941 16524
rect 957 16460 1021 16524
rect 1037 16460 1101 16524
rect 1117 16460 1181 16524
rect 1197 16460 1261 16524
rect 1277 16460 1341 16524
rect 1357 16460 1421 16524
rect 1437 16460 1501 16524
rect 1517 16460 1581 16524
rect 1597 16460 1661 16524
rect 1677 16460 1741 16524
rect 1757 16460 1821 16524
rect 1837 16460 1901 16524
rect 1917 16460 1981 16524
rect 1997 16460 2061 16524
rect 2077 16460 2141 16524
rect 2157 16460 2221 16524
rect 2237 16460 2301 16524
rect 2317 16460 2381 16524
rect 2397 16460 2461 16524
rect 2477 16460 2541 16524
rect 2557 16460 2621 16524
rect 2637 16460 2701 16524
rect 2717 16460 2781 16524
rect 2797 16460 2861 16524
rect 2877 16460 2941 16524
rect 2957 16460 3021 16524
rect 3037 16460 3101 16524
rect 3117 16460 3181 16524
rect 3197 16460 3261 16524
rect 3277 16460 3341 16524
rect 3357 16460 3421 16524
rect 3437 16460 3501 16524
rect 3517 16460 3581 16524
rect 3597 16460 3661 16524
rect 3677 16460 3741 16524
rect 3757 16460 3821 16524
rect 3837 16460 3901 16524
rect 3917 16460 3981 16524
rect 3997 16460 4061 16524
rect 4077 16460 4141 16524
rect 4157 16460 4221 16524
rect 4237 16460 4301 16524
rect 4317 16460 4381 16524
rect 4397 16460 4461 16524
rect 4477 16460 4541 16524
rect 4557 16460 4621 16524
rect 4637 16460 4701 16524
rect 4717 16460 4781 16524
rect 4797 16460 4861 16524
rect 157 16379 221 16443
rect 237 16379 301 16443
rect 317 16379 381 16443
rect 397 16379 461 16443
rect 477 16379 541 16443
rect 557 16379 621 16443
rect 637 16379 701 16443
rect 717 16379 781 16443
rect 797 16379 861 16443
rect 877 16379 941 16443
rect 957 16379 1021 16443
rect 1037 16379 1101 16443
rect 1117 16379 1181 16443
rect 1197 16379 1261 16443
rect 1277 16379 1341 16443
rect 1357 16379 1421 16443
rect 1437 16379 1501 16443
rect 1517 16379 1581 16443
rect 1597 16379 1661 16443
rect 1677 16379 1741 16443
rect 1757 16379 1821 16443
rect 1837 16379 1901 16443
rect 1917 16379 1981 16443
rect 1997 16379 2061 16443
rect 2077 16379 2141 16443
rect 2157 16379 2221 16443
rect 2237 16379 2301 16443
rect 2317 16379 2381 16443
rect 2397 16379 2461 16443
rect 2477 16379 2541 16443
rect 2557 16379 2621 16443
rect 2637 16379 2701 16443
rect 2717 16379 2781 16443
rect 2797 16379 2861 16443
rect 2877 16379 2941 16443
rect 2957 16379 3021 16443
rect 3037 16379 3101 16443
rect 3117 16379 3181 16443
rect 3197 16379 3261 16443
rect 3277 16379 3341 16443
rect 3357 16379 3421 16443
rect 3437 16379 3501 16443
rect 3517 16379 3581 16443
rect 3597 16379 3661 16443
rect 3677 16379 3741 16443
rect 3757 16379 3821 16443
rect 3837 16379 3901 16443
rect 3917 16379 3981 16443
rect 3997 16379 4061 16443
rect 4077 16379 4141 16443
rect 4157 16379 4221 16443
rect 4237 16379 4301 16443
rect 4317 16379 4381 16443
rect 4397 16379 4461 16443
rect 4477 16379 4541 16443
rect 4557 16379 4621 16443
rect 4637 16379 4701 16443
rect 4717 16379 4781 16443
rect 4797 16379 4861 16443
rect 157 16298 221 16362
rect 237 16298 301 16362
rect 317 16298 381 16362
rect 397 16298 461 16362
rect 477 16298 541 16362
rect 557 16298 621 16362
rect 637 16298 701 16362
rect 717 16298 781 16362
rect 797 16298 861 16362
rect 877 16298 941 16362
rect 957 16298 1021 16362
rect 1037 16298 1101 16362
rect 1117 16298 1181 16362
rect 1197 16298 1261 16362
rect 1277 16298 1341 16362
rect 1357 16298 1421 16362
rect 1437 16298 1501 16362
rect 1517 16298 1581 16362
rect 1597 16298 1661 16362
rect 1677 16298 1741 16362
rect 1757 16298 1821 16362
rect 1837 16298 1901 16362
rect 1917 16298 1981 16362
rect 1997 16298 2061 16362
rect 2077 16298 2141 16362
rect 2157 16298 2221 16362
rect 2237 16298 2301 16362
rect 2317 16298 2381 16362
rect 2397 16298 2461 16362
rect 2477 16298 2541 16362
rect 2557 16298 2621 16362
rect 2637 16298 2701 16362
rect 2717 16298 2781 16362
rect 2797 16298 2861 16362
rect 2877 16298 2941 16362
rect 2957 16298 3021 16362
rect 3037 16298 3101 16362
rect 3117 16298 3181 16362
rect 3197 16298 3261 16362
rect 3277 16298 3341 16362
rect 3357 16298 3421 16362
rect 3437 16298 3501 16362
rect 3517 16298 3581 16362
rect 3597 16298 3661 16362
rect 3677 16298 3741 16362
rect 3757 16298 3821 16362
rect 3837 16298 3901 16362
rect 3917 16298 3981 16362
rect 3997 16298 4061 16362
rect 4077 16298 4141 16362
rect 4157 16298 4221 16362
rect 4237 16298 4301 16362
rect 4317 16298 4381 16362
rect 4397 16298 4461 16362
rect 4477 16298 4541 16362
rect 4557 16298 4621 16362
rect 4637 16298 4701 16362
rect 4717 16298 4781 16362
rect 4797 16298 4861 16362
rect 157 16217 221 16281
rect 237 16217 301 16281
rect 317 16217 381 16281
rect 397 16217 461 16281
rect 477 16217 541 16281
rect 557 16217 621 16281
rect 637 16217 701 16281
rect 717 16217 781 16281
rect 797 16217 861 16281
rect 877 16217 941 16281
rect 957 16217 1021 16281
rect 1037 16217 1101 16281
rect 1117 16217 1181 16281
rect 1197 16217 1261 16281
rect 1277 16217 1341 16281
rect 1357 16217 1421 16281
rect 1437 16217 1501 16281
rect 1517 16217 1581 16281
rect 1597 16217 1661 16281
rect 1677 16217 1741 16281
rect 1757 16217 1821 16281
rect 1837 16217 1901 16281
rect 1917 16217 1981 16281
rect 1997 16217 2061 16281
rect 2077 16217 2141 16281
rect 2157 16217 2221 16281
rect 2237 16217 2301 16281
rect 2317 16217 2381 16281
rect 2397 16217 2461 16281
rect 2477 16217 2541 16281
rect 2557 16217 2621 16281
rect 2637 16217 2701 16281
rect 2717 16217 2781 16281
rect 2797 16217 2861 16281
rect 2877 16217 2941 16281
rect 2957 16217 3021 16281
rect 3037 16217 3101 16281
rect 3117 16217 3181 16281
rect 3197 16217 3261 16281
rect 3277 16217 3341 16281
rect 3357 16217 3421 16281
rect 3437 16217 3501 16281
rect 3517 16217 3581 16281
rect 3597 16217 3661 16281
rect 3677 16217 3741 16281
rect 3757 16217 3821 16281
rect 3837 16217 3901 16281
rect 3917 16217 3981 16281
rect 3997 16217 4061 16281
rect 4077 16217 4141 16281
rect 4157 16217 4221 16281
rect 4237 16217 4301 16281
rect 4317 16217 4381 16281
rect 4397 16217 4461 16281
rect 4477 16217 4541 16281
rect 4557 16217 4621 16281
rect 4637 16217 4701 16281
rect 4717 16217 4781 16281
rect 4797 16217 4861 16281
rect 157 16136 221 16200
rect 237 16136 301 16200
rect 317 16136 381 16200
rect 397 16136 461 16200
rect 477 16136 541 16200
rect 557 16136 621 16200
rect 637 16136 701 16200
rect 717 16136 781 16200
rect 797 16136 861 16200
rect 877 16136 941 16200
rect 957 16136 1021 16200
rect 1037 16136 1101 16200
rect 1117 16136 1181 16200
rect 1197 16136 1261 16200
rect 1277 16136 1341 16200
rect 1357 16136 1421 16200
rect 1437 16136 1501 16200
rect 1517 16136 1581 16200
rect 1597 16136 1661 16200
rect 1677 16136 1741 16200
rect 1757 16136 1821 16200
rect 1837 16136 1901 16200
rect 1917 16136 1981 16200
rect 1997 16136 2061 16200
rect 2077 16136 2141 16200
rect 2157 16136 2221 16200
rect 2237 16136 2301 16200
rect 2317 16136 2381 16200
rect 2397 16136 2461 16200
rect 2477 16136 2541 16200
rect 2557 16136 2621 16200
rect 2637 16136 2701 16200
rect 2717 16136 2781 16200
rect 2797 16136 2861 16200
rect 2877 16136 2941 16200
rect 2957 16136 3021 16200
rect 3037 16136 3101 16200
rect 3117 16136 3181 16200
rect 3197 16136 3261 16200
rect 3277 16136 3341 16200
rect 3357 16136 3421 16200
rect 3437 16136 3501 16200
rect 3517 16136 3581 16200
rect 3597 16136 3661 16200
rect 3677 16136 3741 16200
rect 3757 16136 3821 16200
rect 3837 16136 3901 16200
rect 3917 16136 3981 16200
rect 3997 16136 4061 16200
rect 4077 16136 4141 16200
rect 4157 16136 4221 16200
rect 4237 16136 4301 16200
rect 4317 16136 4381 16200
rect 4397 16136 4461 16200
rect 4477 16136 4541 16200
rect 4557 16136 4621 16200
rect 4637 16136 4701 16200
rect 4717 16136 4781 16200
rect 4797 16136 4861 16200
rect 157 16055 221 16119
rect 237 16055 301 16119
rect 317 16055 381 16119
rect 397 16055 461 16119
rect 477 16055 541 16119
rect 557 16055 621 16119
rect 637 16055 701 16119
rect 717 16055 781 16119
rect 797 16055 861 16119
rect 877 16055 941 16119
rect 957 16055 1021 16119
rect 1037 16055 1101 16119
rect 1117 16055 1181 16119
rect 1197 16055 1261 16119
rect 1277 16055 1341 16119
rect 1357 16055 1421 16119
rect 1437 16055 1501 16119
rect 1517 16055 1581 16119
rect 1597 16055 1661 16119
rect 1677 16055 1741 16119
rect 1757 16055 1821 16119
rect 1837 16055 1901 16119
rect 1917 16055 1981 16119
rect 1997 16055 2061 16119
rect 2077 16055 2141 16119
rect 2157 16055 2221 16119
rect 2237 16055 2301 16119
rect 2317 16055 2381 16119
rect 2397 16055 2461 16119
rect 2477 16055 2541 16119
rect 2557 16055 2621 16119
rect 2637 16055 2701 16119
rect 2717 16055 2781 16119
rect 2797 16055 2861 16119
rect 2877 16055 2941 16119
rect 2957 16055 3021 16119
rect 3037 16055 3101 16119
rect 3117 16055 3181 16119
rect 3197 16055 3261 16119
rect 3277 16055 3341 16119
rect 3357 16055 3421 16119
rect 3437 16055 3501 16119
rect 3517 16055 3581 16119
rect 3597 16055 3661 16119
rect 3677 16055 3741 16119
rect 3757 16055 3821 16119
rect 3837 16055 3901 16119
rect 3917 16055 3981 16119
rect 3997 16055 4061 16119
rect 4077 16055 4141 16119
rect 4157 16055 4221 16119
rect 4237 16055 4301 16119
rect 4317 16055 4381 16119
rect 4397 16055 4461 16119
rect 4477 16055 4541 16119
rect 4557 16055 4621 16119
rect 4637 16055 4701 16119
rect 4717 16055 4781 16119
rect 4797 16055 4861 16119
rect 157 15974 221 16038
rect 237 15974 301 16038
rect 317 15974 381 16038
rect 397 15974 461 16038
rect 477 15974 541 16038
rect 557 15974 621 16038
rect 637 15974 701 16038
rect 717 15974 781 16038
rect 797 15974 861 16038
rect 877 15974 941 16038
rect 957 15974 1021 16038
rect 1037 15974 1101 16038
rect 1117 15974 1181 16038
rect 1197 15974 1261 16038
rect 1277 15974 1341 16038
rect 1357 15974 1421 16038
rect 1437 15974 1501 16038
rect 1517 15974 1581 16038
rect 1597 15974 1661 16038
rect 1677 15974 1741 16038
rect 1757 15974 1821 16038
rect 1837 15974 1901 16038
rect 1917 15974 1981 16038
rect 1997 15974 2061 16038
rect 2077 15974 2141 16038
rect 2157 15974 2221 16038
rect 2237 15974 2301 16038
rect 2317 15974 2381 16038
rect 2397 15974 2461 16038
rect 2477 15974 2541 16038
rect 2557 15974 2621 16038
rect 2637 15974 2701 16038
rect 2717 15974 2781 16038
rect 2797 15974 2861 16038
rect 2877 15974 2941 16038
rect 2957 15974 3021 16038
rect 3037 15974 3101 16038
rect 3117 15974 3181 16038
rect 3197 15974 3261 16038
rect 3277 15974 3341 16038
rect 3357 15974 3421 16038
rect 3437 15974 3501 16038
rect 3517 15974 3581 16038
rect 3597 15974 3661 16038
rect 3677 15974 3741 16038
rect 3757 15974 3821 16038
rect 3837 15974 3901 16038
rect 3917 15974 3981 16038
rect 3997 15974 4061 16038
rect 4077 15974 4141 16038
rect 4157 15974 4221 16038
rect 4237 15974 4301 16038
rect 4317 15974 4381 16038
rect 4397 15974 4461 16038
rect 4477 15974 4541 16038
rect 4557 15974 4621 16038
rect 4637 15974 4701 16038
rect 4717 15974 4781 16038
rect 4797 15974 4861 16038
rect 157 15893 221 15957
rect 237 15893 301 15957
rect 317 15893 381 15957
rect 397 15893 461 15957
rect 477 15893 541 15957
rect 557 15893 621 15957
rect 637 15893 701 15957
rect 717 15893 781 15957
rect 797 15893 861 15957
rect 877 15893 941 15957
rect 957 15893 1021 15957
rect 1037 15893 1101 15957
rect 1117 15893 1181 15957
rect 1197 15893 1261 15957
rect 1277 15893 1341 15957
rect 1357 15893 1421 15957
rect 1437 15893 1501 15957
rect 1517 15893 1581 15957
rect 1597 15893 1661 15957
rect 1677 15893 1741 15957
rect 1757 15893 1821 15957
rect 1837 15893 1901 15957
rect 1917 15893 1981 15957
rect 1997 15893 2061 15957
rect 2077 15893 2141 15957
rect 2157 15893 2221 15957
rect 2237 15893 2301 15957
rect 2317 15893 2381 15957
rect 2397 15893 2461 15957
rect 2477 15893 2541 15957
rect 2557 15893 2621 15957
rect 2637 15893 2701 15957
rect 2717 15893 2781 15957
rect 2797 15893 2861 15957
rect 2877 15893 2941 15957
rect 2957 15893 3021 15957
rect 3037 15893 3101 15957
rect 3117 15893 3181 15957
rect 3197 15893 3261 15957
rect 3277 15893 3341 15957
rect 3357 15893 3421 15957
rect 3437 15893 3501 15957
rect 3517 15893 3581 15957
rect 3597 15893 3661 15957
rect 3677 15893 3741 15957
rect 3757 15893 3821 15957
rect 3837 15893 3901 15957
rect 3917 15893 3981 15957
rect 3997 15893 4061 15957
rect 4077 15893 4141 15957
rect 4157 15893 4221 15957
rect 4237 15893 4301 15957
rect 4317 15893 4381 15957
rect 4397 15893 4461 15957
rect 4477 15893 4541 15957
rect 4557 15893 4621 15957
rect 4637 15893 4701 15957
rect 4717 15893 4781 15957
rect 4797 15893 4861 15957
rect 157 15812 221 15876
rect 237 15812 301 15876
rect 317 15812 381 15876
rect 397 15812 461 15876
rect 477 15812 541 15876
rect 557 15812 621 15876
rect 637 15812 701 15876
rect 717 15812 781 15876
rect 797 15812 861 15876
rect 877 15812 941 15876
rect 957 15812 1021 15876
rect 1037 15812 1101 15876
rect 1117 15812 1181 15876
rect 1197 15812 1261 15876
rect 1277 15812 1341 15876
rect 1357 15812 1421 15876
rect 1437 15812 1501 15876
rect 1517 15812 1581 15876
rect 1597 15812 1661 15876
rect 1677 15812 1741 15876
rect 1757 15812 1821 15876
rect 1837 15812 1901 15876
rect 1917 15812 1981 15876
rect 1997 15812 2061 15876
rect 2077 15812 2141 15876
rect 2157 15812 2221 15876
rect 2237 15812 2301 15876
rect 2317 15812 2381 15876
rect 2397 15812 2461 15876
rect 2477 15812 2541 15876
rect 2557 15812 2621 15876
rect 2637 15812 2701 15876
rect 2717 15812 2781 15876
rect 2797 15812 2861 15876
rect 2877 15812 2941 15876
rect 2957 15812 3021 15876
rect 3037 15812 3101 15876
rect 3117 15812 3181 15876
rect 3197 15812 3261 15876
rect 3277 15812 3341 15876
rect 3357 15812 3421 15876
rect 3437 15812 3501 15876
rect 3517 15812 3581 15876
rect 3597 15812 3661 15876
rect 3677 15812 3741 15876
rect 3757 15812 3821 15876
rect 3837 15812 3901 15876
rect 3917 15812 3981 15876
rect 3997 15812 4061 15876
rect 4077 15812 4141 15876
rect 4157 15812 4221 15876
rect 4237 15812 4301 15876
rect 4317 15812 4381 15876
rect 4397 15812 4461 15876
rect 4477 15812 4541 15876
rect 4557 15812 4621 15876
rect 4637 15812 4701 15876
rect 4717 15812 4781 15876
rect 4797 15812 4861 15876
rect 157 15731 221 15795
rect 237 15731 301 15795
rect 317 15731 381 15795
rect 397 15731 461 15795
rect 477 15731 541 15795
rect 557 15731 621 15795
rect 637 15731 701 15795
rect 717 15731 781 15795
rect 797 15731 861 15795
rect 877 15731 941 15795
rect 957 15731 1021 15795
rect 1037 15731 1101 15795
rect 1117 15731 1181 15795
rect 1197 15731 1261 15795
rect 1277 15731 1341 15795
rect 1357 15731 1421 15795
rect 1437 15731 1501 15795
rect 1517 15731 1581 15795
rect 1597 15731 1661 15795
rect 1677 15731 1741 15795
rect 1757 15731 1821 15795
rect 1837 15731 1901 15795
rect 1917 15731 1981 15795
rect 1997 15731 2061 15795
rect 2077 15731 2141 15795
rect 2157 15731 2221 15795
rect 2237 15731 2301 15795
rect 2317 15731 2381 15795
rect 2397 15731 2461 15795
rect 2477 15731 2541 15795
rect 2557 15731 2621 15795
rect 2637 15731 2701 15795
rect 2717 15731 2781 15795
rect 2797 15731 2861 15795
rect 2877 15731 2941 15795
rect 2957 15731 3021 15795
rect 3037 15731 3101 15795
rect 3117 15731 3181 15795
rect 3197 15731 3261 15795
rect 3277 15731 3341 15795
rect 3357 15731 3421 15795
rect 3437 15731 3501 15795
rect 3517 15731 3581 15795
rect 3597 15731 3661 15795
rect 3677 15731 3741 15795
rect 3757 15731 3821 15795
rect 3837 15731 3901 15795
rect 3917 15731 3981 15795
rect 3997 15731 4061 15795
rect 4077 15731 4141 15795
rect 4157 15731 4221 15795
rect 4237 15731 4301 15795
rect 4317 15731 4381 15795
rect 4397 15731 4461 15795
rect 4477 15731 4541 15795
rect 4557 15731 4621 15795
rect 4637 15731 4701 15795
rect 4717 15731 4781 15795
rect 4797 15731 4861 15795
rect 157 15650 221 15714
rect 237 15650 301 15714
rect 317 15650 381 15714
rect 397 15650 461 15714
rect 477 15650 541 15714
rect 557 15650 621 15714
rect 637 15650 701 15714
rect 717 15650 781 15714
rect 797 15650 861 15714
rect 877 15650 941 15714
rect 957 15650 1021 15714
rect 1037 15650 1101 15714
rect 1117 15650 1181 15714
rect 1197 15650 1261 15714
rect 1277 15650 1341 15714
rect 1357 15650 1421 15714
rect 1437 15650 1501 15714
rect 1517 15650 1581 15714
rect 1597 15650 1661 15714
rect 1677 15650 1741 15714
rect 1757 15650 1821 15714
rect 1837 15650 1901 15714
rect 1917 15650 1981 15714
rect 1997 15650 2061 15714
rect 2077 15650 2141 15714
rect 2157 15650 2221 15714
rect 2237 15650 2301 15714
rect 2317 15650 2381 15714
rect 2397 15650 2461 15714
rect 2477 15650 2541 15714
rect 2557 15650 2621 15714
rect 2637 15650 2701 15714
rect 2717 15650 2781 15714
rect 2797 15650 2861 15714
rect 2877 15650 2941 15714
rect 2957 15650 3021 15714
rect 3037 15650 3101 15714
rect 3117 15650 3181 15714
rect 3197 15650 3261 15714
rect 3277 15650 3341 15714
rect 3357 15650 3421 15714
rect 3437 15650 3501 15714
rect 3517 15650 3581 15714
rect 3597 15650 3661 15714
rect 3677 15650 3741 15714
rect 3757 15650 3821 15714
rect 3837 15650 3901 15714
rect 3917 15650 3981 15714
rect 3997 15650 4061 15714
rect 4077 15650 4141 15714
rect 4157 15650 4221 15714
rect 4237 15650 4301 15714
rect 4317 15650 4381 15714
rect 4397 15650 4461 15714
rect 4477 15650 4541 15714
rect 4557 15650 4621 15714
rect 4637 15650 4701 15714
rect 4717 15650 4781 15714
rect 4797 15650 4861 15714
rect 157 15569 221 15633
rect 237 15569 301 15633
rect 317 15569 381 15633
rect 397 15569 461 15633
rect 477 15569 541 15633
rect 557 15569 621 15633
rect 637 15569 701 15633
rect 717 15569 781 15633
rect 797 15569 861 15633
rect 877 15569 941 15633
rect 957 15569 1021 15633
rect 1037 15569 1101 15633
rect 1117 15569 1181 15633
rect 1197 15569 1261 15633
rect 1277 15569 1341 15633
rect 1357 15569 1421 15633
rect 1437 15569 1501 15633
rect 1517 15569 1581 15633
rect 1597 15569 1661 15633
rect 1677 15569 1741 15633
rect 1757 15569 1821 15633
rect 1837 15569 1901 15633
rect 1917 15569 1981 15633
rect 1997 15569 2061 15633
rect 2077 15569 2141 15633
rect 2157 15569 2221 15633
rect 2237 15569 2301 15633
rect 2317 15569 2381 15633
rect 2397 15569 2461 15633
rect 2477 15569 2541 15633
rect 2557 15569 2621 15633
rect 2637 15569 2701 15633
rect 2717 15569 2781 15633
rect 2797 15569 2861 15633
rect 2877 15569 2941 15633
rect 2957 15569 3021 15633
rect 3037 15569 3101 15633
rect 3117 15569 3181 15633
rect 3197 15569 3261 15633
rect 3277 15569 3341 15633
rect 3357 15569 3421 15633
rect 3437 15569 3501 15633
rect 3517 15569 3581 15633
rect 3597 15569 3661 15633
rect 3677 15569 3741 15633
rect 3757 15569 3821 15633
rect 3837 15569 3901 15633
rect 3917 15569 3981 15633
rect 3997 15569 4061 15633
rect 4077 15569 4141 15633
rect 4157 15569 4221 15633
rect 4237 15569 4301 15633
rect 4317 15569 4381 15633
rect 4397 15569 4461 15633
rect 4477 15569 4541 15633
rect 4557 15569 4621 15633
rect 4637 15569 4701 15633
rect 4717 15569 4781 15633
rect 4797 15569 4861 15633
rect 157 15488 221 15552
rect 237 15488 301 15552
rect 317 15488 381 15552
rect 397 15488 461 15552
rect 477 15488 541 15552
rect 557 15488 621 15552
rect 637 15488 701 15552
rect 717 15488 781 15552
rect 797 15488 861 15552
rect 877 15488 941 15552
rect 957 15488 1021 15552
rect 1037 15488 1101 15552
rect 1117 15488 1181 15552
rect 1197 15488 1261 15552
rect 1277 15488 1341 15552
rect 1357 15488 1421 15552
rect 1437 15488 1501 15552
rect 1517 15488 1581 15552
rect 1597 15488 1661 15552
rect 1677 15488 1741 15552
rect 1757 15488 1821 15552
rect 1837 15488 1901 15552
rect 1917 15488 1981 15552
rect 1997 15488 2061 15552
rect 2077 15488 2141 15552
rect 2157 15488 2221 15552
rect 2237 15488 2301 15552
rect 2317 15488 2381 15552
rect 2397 15488 2461 15552
rect 2477 15488 2541 15552
rect 2557 15488 2621 15552
rect 2637 15488 2701 15552
rect 2717 15488 2781 15552
rect 2797 15488 2861 15552
rect 2877 15488 2941 15552
rect 2957 15488 3021 15552
rect 3037 15488 3101 15552
rect 3117 15488 3181 15552
rect 3197 15488 3261 15552
rect 3277 15488 3341 15552
rect 3357 15488 3421 15552
rect 3437 15488 3501 15552
rect 3517 15488 3581 15552
rect 3597 15488 3661 15552
rect 3677 15488 3741 15552
rect 3757 15488 3821 15552
rect 3837 15488 3901 15552
rect 3917 15488 3981 15552
rect 3997 15488 4061 15552
rect 4077 15488 4141 15552
rect 4157 15488 4221 15552
rect 4237 15488 4301 15552
rect 4317 15488 4381 15552
rect 4397 15488 4461 15552
rect 4477 15488 4541 15552
rect 4557 15488 4621 15552
rect 4637 15488 4701 15552
rect 4717 15488 4781 15552
rect 4797 15488 4861 15552
rect 157 15407 221 15471
rect 237 15407 301 15471
rect 317 15407 381 15471
rect 397 15407 461 15471
rect 477 15407 541 15471
rect 557 15407 621 15471
rect 637 15407 701 15471
rect 717 15407 781 15471
rect 797 15407 861 15471
rect 877 15407 941 15471
rect 957 15407 1021 15471
rect 1037 15407 1101 15471
rect 1117 15407 1181 15471
rect 1197 15407 1261 15471
rect 1277 15407 1341 15471
rect 1357 15407 1421 15471
rect 1437 15407 1501 15471
rect 1517 15407 1581 15471
rect 1597 15407 1661 15471
rect 1677 15407 1741 15471
rect 1757 15407 1821 15471
rect 1837 15407 1901 15471
rect 1917 15407 1981 15471
rect 1997 15407 2061 15471
rect 2077 15407 2141 15471
rect 2157 15407 2221 15471
rect 2237 15407 2301 15471
rect 2317 15407 2381 15471
rect 2397 15407 2461 15471
rect 2477 15407 2541 15471
rect 2557 15407 2621 15471
rect 2637 15407 2701 15471
rect 2717 15407 2781 15471
rect 2797 15407 2861 15471
rect 2877 15407 2941 15471
rect 2957 15407 3021 15471
rect 3037 15407 3101 15471
rect 3117 15407 3181 15471
rect 3197 15407 3261 15471
rect 3277 15407 3341 15471
rect 3357 15407 3421 15471
rect 3437 15407 3501 15471
rect 3517 15407 3581 15471
rect 3597 15407 3661 15471
rect 3677 15407 3741 15471
rect 3757 15407 3821 15471
rect 3837 15407 3901 15471
rect 3917 15407 3981 15471
rect 3997 15407 4061 15471
rect 4077 15407 4141 15471
rect 4157 15407 4221 15471
rect 4237 15407 4301 15471
rect 4317 15407 4381 15471
rect 4397 15407 4461 15471
rect 4477 15407 4541 15471
rect 4557 15407 4621 15471
rect 4637 15407 4701 15471
rect 4717 15407 4781 15471
rect 4797 15407 4861 15471
rect 157 15326 221 15390
rect 237 15326 301 15390
rect 317 15326 381 15390
rect 397 15326 461 15390
rect 477 15326 541 15390
rect 557 15326 621 15390
rect 637 15326 701 15390
rect 717 15326 781 15390
rect 797 15326 861 15390
rect 877 15326 941 15390
rect 957 15326 1021 15390
rect 1037 15326 1101 15390
rect 1117 15326 1181 15390
rect 1197 15326 1261 15390
rect 1277 15326 1341 15390
rect 1357 15326 1421 15390
rect 1437 15326 1501 15390
rect 1517 15326 1581 15390
rect 1597 15326 1661 15390
rect 1677 15326 1741 15390
rect 1757 15326 1821 15390
rect 1837 15326 1901 15390
rect 1917 15326 1981 15390
rect 1997 15326 2061 15390
rect 2077 15326 2141 15390
rect 2157 15326 2221 15390
rect 2237 15326 2301 15390
rect 2317 15326 2381 15390
rect 2397 15326 2461 15390
rect 2477 15326 2541 15390
rect 2557 15326 2621 15390
rect 2637 15326 2701 15390
rect 2717 15326 2781 15390
rect 2797 15326 2861 15390
rect 2877 15326 2941 15390
rect 2957 15326 3021 15390
rect 3037 15326 3101 15390
rect 3117 15326 3181 15390
rect 3197 15326 3261 15390
rect 3277 15326 3341 15390
rect 3357 15326 3421 15390
rect 3437 15326 3501 15390
rect 3517 15326 3581 15390
rect 3597 15326 3661 15390
rect 3677 15326 3741 15390
rect 3757 15326 3821 15390
rect 3837 15326 3901 15390
rect 3917 15326 3981 15390
rect 3997 15326 4061 15390
rect 4077 15326 4141 15390
rect 4157 15326 4221 15390
rect 4237 15326 4301 15390
rect 4317 15326 4381 15390
rect 4397 15326 4461 15390
rect 4477 15326 4541 15390
rect 4557 15326 4621 15390
rect 4637 15326 4701 15390
rect 4717 15326 4781 15390
rect 4797 15326 4861 15390
rect 157 15245 221 15309
rect 237 15245 301 15309
rect 317 15245 381 15309
rect 397 15245 461 15309
rect 477 15245 541 15309
rect 557 15245 621 15309
rect 637 15245 701 15309
rect 717 15245 781 15309
rect 797 15245 861 15309
rect 877 15245 941 15309
rect 957 15245 1021 15309
rect 1037 15245 1101 15309
rect 1117 15245 1181 15309
rect 1197 15245 1261 15309
rect 1277 15245 1341 15309
rect 1357 15245 1421 15309
rect 1437 15245 1501 15309
rect 1517 15245 1581 15309
rect 1597 15245 1661 15309
rect 1677 15245 1741 15309
rect 1757 15245 1821 15309
rect 1837 15245 1901 15309
rect 1917 15245 1981 15309
rect 1997 15245 2061 15309
rect 2077 15245 2141 15309
rect 2157 15245 2221 15309
rect 2237 15245 2301 15309
rect 2317 15245 2381 15309
rect 2397 15245 2461 15309
rect 2477 15245 2541 15309
rect 2557 15245 2621 15309
rect 2637 15245 2701 15309
rect 2717 15245 2781 15309
rect 2797 15245 2861 15309
rect 2877 15245 2941 15309
rect 2957 15245 3021 15309
rect 3037 15245 3101 15309
rect 3117 15245 3181 15309
rect 3197 15245 3261 15309
rect 3277 15245 3341 15309
rect 3357 15245 3421 15309
rect 3437 15245 3501 15309
rect 3517 15245 3581 15309
rect 3597 15245 3661 15309
rect 3677 15245 3741 15309
rect 3757 15245 3821 15309
rect 3837 15245 3901 15309
rect 3917 15245 3981 15309
rect 3997 15245 4061 15309
rect 4077 15245 4141 15309
rect 4157 15245 4221 15309
rect 4237 15245 4301 15309
rect 4317 15245 4381 15309
rect 4397 15245 4461 15309
rect 4477 15245 4541 15309
rect 4557 15245 4621 15309
rect 4637 15245 4701 15309
rect 4717 15245 4781 15309
rect 4797 15245 4861 15309
rect 157 15164 221 15228
rect 237 15164 301 15228
rect 317 15164 381 15228
rect 397 15164 461 15228
rect 477 15164 541 15228
rect 557 15164 621 15228
rect 637 15164 701 15228
rect 717 15164 781 15228
rect 797 15164 861 15228
rect 877 15164 941 15228
rect 957 15164 1021 15228
rect 1037 15164 1101 15228
rect 1117 15164 1181 15228
rect 1197 15164 1261 15228
rect 1277 15164 1341 15228
rect 1357 15164 1421 15228
rect 1437 15164 1501 15228
rect 1517 15164 1581 15228
rect 1597 15164 1661 15228
rect 1677 15164 1741 15228
rect 1757 15164 1821 15228
rect 1837 15164 1901 15228
rect 1917 15164 1981 15228
rect 1997 15164 2061 15228
rect 2077 15164 2141 15228
rect 2157 15164 2221 15228
rect 2237 15164 2301 15228
rect 2317 15164 2381 15228
rect 2397 15164 2461 15228
rect 2477 15164 2541 15228
rect 2557 15164 2621 15228
rect 2637 15164 2701 15228
rect 2717 15164 2781 15228
rect 2797 15164 2861 15228
rect 2877 15164 2941 15228
rect 2957 15164 3021 15228
rect 3037 15164 3101 15228
rect 3117 15164 3181 15228
rect 3197 15164 3261 15228
rect 3277 15164 3341 15228
rect 3357 15164 3421 15228
rect 3437 15164 3501 15228
rect 3517 15164 3581 15228
rect 3597 15164 3661 15228
rect 3677 15164 3741 15228
rect 3757 15164 3821 15228
rect 3837 15164 3901 15228
rect 3917 15164 3981 15228
rect 3997 15164 4061 15228
rect 4077 15164 4141 15228
rect 4157 15164 4221 15228
rect 4237 15164 4301 15228
rect 4317 15164 4381 15228
rect 4397 15164 4461 15228
rect 4477 15164 4541 15228
rect 4557 15164 4621 15228
rect 4637 15164 4701 15228
rect 4717 15164 4781 15228
rect 4797 15164 4861 15228
rect 157 15083 221 15147
rect 237 15083 301 15147
rect 317 15083 381 15147
rect 397 15083 461 15147
rect 477 15083 541 15147
rect 557 15083 621 15147
rect 637 15083 701 15147
rect 717 15083 781 15147
rect 797 15083 861 15147
rect 877 15083 941 15147
rect 957 15083 1021 15147
rect 1037 15083 1101 15147
rect 1117 15083 1181 15147
rect 1197 15083 1261 15147
rect 1277 15083 1341 15147
rect 1357 15083 1421 15147
rect 1437 15083 1501 15147
rect 1517 15083 1581 15147
rect 1597 15083 1661 15147
rect 1677 15083 1741 15147
rect 1757 15083 1821 15147
rect 1837 15083 1901 15147
rect 1917 15083 1981 15147
rect 1997 15083 2061 15147
rect 2077 15083 2141 15147
rect 2157 15083 2221 15147
rect 2237 15083 2301 15147
rect 2317 15083 2381 15147
rect 2397 15083 2461 15147
rect 2477 15083 2541 15147
rect 2557 15083 2621 15147
rect 2637 15083 2701 15147
rect 2717 15083 2781 15147
rect 2797 15083 2861 15147
rect 2877 15083 2941 15147
rect 2957 15083 3021 15147
rect 3037 15083 3101 15147
rect 3117 15083 3181 15147
rect 3197 15083 3261 15147
rect 3277 15083 3341 15147
rect 3357 15083 3421 15147
rect 3437 15083 3501 15147
rect 3517 15083 3581 15147
rect 3597 15083 3661 15147
rect 3677 15083 3741 15147
rect 3757 15083 3821 15147
rect 3837 15083 3901 15147
rect 3917 15083 3981 15147
rect 3997 15083 4061 15147
rect 4077 15083 4141 15147
rect 4157 15083 4221 15147
rect 4237 15083 4301 15147
rect 4317 15083 4381 15147
rect 4397 15083 4461 15147
rect 4477 15083 4541 15147
rect 4557 15083 4621 15147
rect 4637 15083 4701 15147
rect 4717 15083 4781 15147
rect 4797 15083 4861 15147
rect 157 15002 221 15066
rect 237 15002 301 15066
rect 317 15002 381 15066
rect 397 15002 461 15066
rect 477 15002 541 15066
rect 557 15002 621 15066
rect 637 15002 701 15066
rect 717 15002 781 15066
rect 797 15002 861 15066
rect 877 15002 941 15066
rect 957 15002 1021 15066
rect 1037 15002 1101 15066
rect 1117 15002 1181 15066
rect 1197 15002 1261 15066
rect 1277 15002 1341 15066
rect 1357 15002 1421 15066
rect 1437 15002 1501 15066
rect 1517 15002 1581 15066
rect 1597 15002 1661 15066
rect 1677 15002 1741 15066
rect 1757 15002 1821 15066
rect 1837 15002 1901 15066
rect 1917 15002 1981 15066
rect 1997 15002 2061 15066
rect 2077 15002 2141 15066
rect 2157 15002 2221 15066
rect 2237 15002 2301 15066
rect 2317 15002 2381 15066
rect 2397 15002 2461 15066
rect 2477 15002 2541 15066
rect 2557 15002 2621 15066
rect 2637 15002 2701 15066
rect 2717 15002 2781 15066
rect 2797 15002 2861 15066
rect 2877 15002 2941 15066
rect 2957 15002 3021 15066
rect 3037 15002 3101 15066
rect 3117 15002 3181 15066
rect 3197 15002 3261 15066
rect 3277 15002 3341 15066
rect 3357 15002 3421 15066
rect 3437 15002 3501 15066
rect 3517 15002 3581 15066
rect 3597 15002 3661 15066
rect 3677 15002 3741 15066
rect 3757 15002 3821 15066
rect 3837 15002 3901 15066
rect 3917 15002 3981 15066
rect 3997 15002 4061 15066
rect 4077 15002 4141 15066
rect 4157 15002 4221 15066
rect 4237 15002 4301 15066
rect 4317 15002 4381 15066
rect 4397 15002 4461 15066
rect 4477 15002 4541 15066
rect 4557 15002 4621 15066
rect 4637 15002 4701 15066
rect 4717 15002 4781 15066
rect 4797 15002 4861 15066
rect 157 14921 221 14985
rect 237 14921 301 14985
rect 317 14921 381 14985
rect 397 14921 461 14985
rect 477 14921 541 14985
rect 557 14921 621 14985
rect 637 14921 701 14985
rect 717 14921 781 14985
rect 797 14921 861 14985
rect 877 14921 941 14985
rect 957 14921 1021 14985
rect 1037 14921 1101 14985
rect 1117 14921 1181 14985
rect 1197 14921 1261 14985
rect 1277 14921 1341 14985
rect 1357 14921 1421 14985
rect 1437 14921 1501 14985
rect 1517 14921 1581 14985
rect 1597 14921 1661 14985
rect 1677 14921 1741 14985
rect 1757 14921 1821 14985
rect 1837 14921 1901 14985
rect 1917 14921 1981 14985
rect 1997 14921 2061 14985
rect 2077 14921 2141 14985
rect 2157 14921 2221 14985
rect 2237 14921 2301 14985
rect 2317 14921 2381 14985
rect 2397 14921 2461 14985
rect 2477 14921 2541 14985
rect 2557 14921 2621 14985
rect 2637 14921 2701 14985
rect 2717 14921 2781 14985
rect 2797 14921 2861 14985
rect 2877 14921 2941 14985
rect 2957 14921 3021 14985
rect 3037 14921 3101 14985
rect 3117 14921 3181 14985
rect 3197 14921 3261 14985
rect 3277 14921 3341 14985
rect 3357 14921 3421 14985
rect 3437 14921 3501 14985
rect 3517 14921 3581 14985
rect 3597 14921 3661 14985
rect 3677 14921 3741 14985
rect 3757 14921 3821 14985
rect 3837 14921 3901 14985
rect 3917 14921 3981 14985
rect 3997 14921 4061 14985
rect 4077 14921 4141 14985
rect 4157 14921 4221 14985
rect 4237 14921 4301 14985
rect 4317 14921 4381 14985
rect 4397 14921 4461 14985
rect 4477 14921 4541 14985
rect 4557 14921 4621 14985
rect 4637 14921 4701 14985
rect 4717 14921 4781 14985
rect 4797 14921 4861 14985
rect 157 14840 221 14904
rect 237 14840 301 14904
rect 317 14840 381 14904
rect 397 14840 461 14904
rect 477 14840 541 14904
rect 557 14840 621 14904
rect 637 14840 701 14904
rect 717 14840 781 14904
rect 797 14840 861 14904
rect 877 14840 941 14904
rect 957 14840 1021 14904
rect 1037 14840 1101 14904
rect 1117 14840 1181 14904
rect 1197 14840 1261 14904
rect 1277 14840 1341 14904
rect 1357 14840 1421 14904
rect 1437 14840 1501 14904
rect 1517 14840 1581 14904
rect 1597 14840 1661 14904
rect 1677 14840 1741 14904
rect 1757 14840 1821 14904
rect 1837 14840 1901 14904
rect 1917 14840 1981 14904
rect 1997 14840 2061 14904
rect 2077 14840 2141 14904
rect 2157 14840 2221 14904
rect 2237 14840 2301 14904
rect 2317 14840 2381 14904
rect 2397 14840 2461 14904
rect 2477 14840 2541 14904
rect 2557 14840 2621 14904
rect 2637 14840 2701 14904
rect 2717 14840 2781 14904
rect 2797 14840 2861 14904
rect 2877 14840 2941 14904
rect 2957 14840 3021 14904
rect 3037 14840 3101 14904
rect 3117 14840 3181 14904
rect 3197 14840 3261 14904
rect 3277 14840 3341 14904
rect 3357 14840 3421 14904
rect 3437 14840 3501 14904
rect 3517 14840 3581 14904
rect 3597 14840 3661 14904
rect 3677 14840 3741 14904
rect 3757 14840 3821 14904
rect 3837 14840 3901 14904
rect 3917 14840 3981 14904
rect 3997 14840 4061 14904
rect 4077 14840 4141 14904
rect 4157 14840 4221 14904
rect 4237 14840 4301 14904
rect 4317 14840 4381 14904
rect 4397 14840 4461 14904
rect 4477 14840 4541 14904
rect 4557 14840 4621 14904
rect 4637 14840 4701 14904
rect 4717 14840 4781 14904
rect 4797 14840 4861 14904
rect 157 14759 221 14823
rect 237 14759 301 14823
rect 317 14759 381 14823
rect 397 14759 461 14823
rect 477 14759 541 14823
rect 557 14759 621 14823
rect 637 14759 701 14823
rect 717 14759 781 14823
rect 797 14759 861 14823
rect 877 14759 941 14823
rect 957 14759 1021 14823
rect 1037 14759 1101 14823
rect 1117 14759 1181 14823
rect 1197 14759 1261 14823
rect 1277 14759 1341 14823
rect 1357 14759 1421 14823
rect 1437 14759 1501 14823
rect 1517 14759 1581 14823
rect 1597 14759 1661 14823
rect 1677 14759 1741 14823
rect 1757 14759 1821 14823
rect 1837 14759 1901 14823
rect 1917 14759 1981 14823
rect 1997 14759 2061 14823
rect 2077 14759 2141 14823
rect 2157 14759 2221 14823
rect 2237 14759 2301 14823
rect 2317 14759 2381 14823
rect 2397 14759 2461 14823
rect 2477 14759 2541 14823
rect 2557 14759 2621 14823
rect 2637 14759 2701 14823
rect 2717 14759 2781 14823
rect 2797 14759 2861 14823
rect 2877 14759 2941 14823
rect 2957 14759 3021 14823
rect 3037 14759 3101 14823
rect 3117 14759 3181 14823
rect 3197 14759 3261 14823
rect 3277 14759 3341 14823
rect 3357 14759 3421 14823
rect 3437 14759 3501 14823
rect 3517 14759 3581 14823
rect 3597 14759 3661 14823
rect 3677 14759 3741 14823
rect 3757 14759 3821 14823
rect 3837 14759 3901 14823
rect 3917 14759 3981 14823
rect 3997 14759 4061 14823
rect 4077 14759 4141 14823
rect 4157 14759 4221 14823
rect 4237 14759 4301 14823
rect 4317 14759 4381 14823
rect 4397 14759 4461 14823
rect 4477 14759 4541 14823
rect 4557 14759 4621 14823
rect 4637 14759 4701 14823
rect 4717 14759 4781 14823
rect 4797 14759 4861 14823
rect 157 14678 221 14742
rect 237 14678 301 14742
rect 317 14678 381 14742
rect 397 14678 461 14742
rect 477 14678 541 14742
rect 557 14678 621 14742
rect 637 14678 701 14742
rect 717 14678 781 14742
rect 797 14678 861 14742
rect 877 14678 941 14742
rect 957 14678 1021 14742
rect 1037 14678 1101 14742
rect 1117 14678 1181 14742
rect 1197 14678 1261 14742
rect 1277 14678 1341 14742
rect 1357 14678 1421 14742
rect 1437 14678 1501 14742
rect 1517 14678 1581 14742
rect 1597 14678 1661 14742
rect 1677 14678 1741 14742
rect 1757 14678 1821 14742
rect 1837 14678 1901 14742
rect 1917 14678 1981 14742
rect 1997 14678 2061 14742
rect 2077 14678 2141 14742
rect 2157 14678 2221 14742
rect 2237 14678 2301 14742
rect 2317 14678 2381 14742
rect 2397 14678 2461 14742
rect 2477 14678 2541 14742
rect 2557 14678 2621 14742
rect 2637 14678 2701 14742
rect 2717 14678 2781 14742
rect 2797 14678 2861 14742
rect 2877 14678 2941 14742
rect 2957 14678 3021 14742
rect 3037 14678 3101 14742
rect 3117 14678 3181 14742
rect 3197 14678 3261 14742
rect 3277 14678 3341 14742
rect 3357 14678 3421 14742
rect 3437 14678 3501 14742
rect 3517 14678 3581 14742
rect 3597 14678 3661 14742
rect 3677 14678 3741 14742
rect 3757 14678 3821 14742
rect 3837 14678 3901 14742
rect 3917 14678 3981 14742
rect 3997 14678 4061 14742
rect 4077 14678 4141 14742
rect 4157 14678 4221 14742
rect 4237 14678 4301 14742
rect 4317 14678 4381 14742
rect 4397 14678 4461 14742
rect 4477 14678 4541 14742
rect 4557 14678 4621 14742
rect 4637 14678 4701 14742
rect 4717 14678 4781 14742
rect 4797 14678 4861 14742
rect 157 14597 221 14661
rect 237 14597 301 14661
rect 317 14597 381 14661
rect 397 14597 461 14661
rect 477 14597 541 14661
rect 557 14597 621 14661
rect 637 14597 701 14661
rect 717 14597 781 14661
rect 797 14597 861 14661
rect 877 14597 941 14661
rect 957 14597 1021 14661
rect 1037 14597 1101 14661
rect 1117 14597 1181 14661
rect 1197 14597 1261 14661
rect 1277 14597 1341 14661
rect 1357 14597 1421 14661
rect 1437 14597 1501 14661
rect 1517 14597 1581 14661
rect 1597 14597 1661 14661
rect 1677 14597 1741 14661
rect 1757 14597 1821 14661
rect 1837 14597 1901 14661
rect 1917 14597 1981 14661
rect 1997 14597 2061 14661
rect 2077 14597 2141 14661
rect 2157 14597 2221 14661
rect 2237 14597 2301 14661
rect 2317 14597 2381 14661
rect 2397 14597 2461 14661
rect 2477 14597 2541 14661
rect 2557 14597 2621 14661
rect 2637 14597 2701 14661
rect 2717 14597 2781 14661
rect 2797 14597 2861 14661
rect 2877 14597 2941 14661
rect 2957 14597 3021 14661
rect 3037 14597 3101 14661
rect 3117 14597 3181 14661
rect 3197 14597 3261 14661
rect 3277 14597 3341 14661
rect 3357 14597 3421 14661
rect 3437 14597 3501 14661
rect 3517 14597 3581 14661
rect 3597 14597 3661 14661
rect 3677 14597 3741 14661
rect 3757 14597 3821 14661
rect 3837 14597 3901 14661
rect 3917 14597 3981 14661
rect 3997 14597 4061 14661
rect 4077 14597 4141 14661
rect 4157 14597 4221 14661
rect 4237 14597 4301 14661
rect 4317 14597 4381 14661
rect 4397 14597 4461 14661
rect 4477 14597 4541 14661
rect 4557 14597 4621 14661
rect 4637 14597 4701 14661
rect 4717 14597 4781 14661
rect 4797 14597 4861 14661
rect 157 14515 221 14579
rect 237 14515 301 14579
rect 317 14515 381 14579
rect 397 14515 461 14579
rect 477 14515 541 14579
rect 557 14515 621 14579
rect 637 14515 701 14579
rect 717 14515 781 14579
rect 797 14515 861 14579
rect 877 14515 941 14579
rect 957 14515 1021 14579
rect 1037 14515 1101 14579
rect 1117 14515 1181 14579
rect 1197 14515 1261 14579
rect 1277 14515 1341 14579
rect 1357 14515 1421 14579
rect 1437 14515 1501 14579
rect 1517 14515 1581 14579
rect 1597 14515 1661 14579
rect 1677 14515 1741 14579
rect 1757 14515 1821 14579
rect 1837 14515 1901 14579
rect 1917 14515 1981 14579
rect 1997 14515 2061 14579
rect 2077 14515 2141 14579
rect 2157 14515 2221 14579
rect 2237 14515 2301 14579
rect 2317 14515 2381 14579
rect 2397 14515 2461 14579
rect 2477 14515 2541 14579
rect 2557 14515 2621 14579
rect 2637 14515 2701 14579
rect 2717 14515 2781 14579
rect 2797 14515 2861 14579
rect 2877 14515 2941 14579
rect 2957 14515 3021 14579
rect 3037 14515 3101 14579
rect 3117 14515 3181 14579
rect 3197 14515 3261 14579
rect 3277 14515 3341 14579
rect 3357 14515 3421 14579
rect 3437 14515 3501 14579
rect 3517 14515 3581 14579
rect 3597 14515 3661 14579
rect 3677 14515 3741 14579
rect 3757 14515 3821 14579
rect 3837 14515 3901 14579
rect 3917 14515 3981 14579
rect 3997 14515 4061 14579
rect 4077 14515 4141 14579
rect 4157 14515 4221 14579
rect 4237 14515 4301 14579
rect 4317 14515 4381 14579
rect 4397 14515 4461 14579
rect 4477 14515 4541 14579
rect 4557 14515 4621 14579
rect 4637 14515 4701 14579
rect 4717 14515 4781 14579
rect 4797 14515 4861 14579
rect 157 14433 221 14497
rect 237 14433 301 14497
rect 317 14433 381 14497
rect 397 14433 461 14497
rect 477 14433 541 14497
rect 557 14433 621 14497
rect 637 14433 701 14497
rect 717 14433 781 14497
rect 797 14433 861 14497
rect 877 14433 941 14497
rect 957 14433 1021 14497
rect 1037 14433 1101 14497
rect 1117 14433 1181 14497
rect 1197 14433 1261 14497
rect 1277 14433 1341 14497
rect 1357 14433 1421 14497
rect 1437 14433 1501 14497
rect 1517 14433 1581 14497
rect 1597 14433 1661 14497
rect 1677 14433 1741 14497
rect 1757 14433 1821 14497
rect 1837 14433 1901 14497
rect 1917 14433 1981 14497
rect 1997 14433 2061 14497
rect 2077 14433 2141 14497
rect 2157 14433 2221 14497
rect 2237 14433 2301 14497
rect 2317 14433 2381 14497
rect 2397 14433 2461 14497
rect 2477 14433 2541 14497
rect 2557 14433 2621 14497
rect 2637 14433 2701 14497
rect 2717 14433 2781 14497
rect 2797 14433 2861 14497
rect 2877 14433 2941 14497
rect 2957 14433 3021 14497
rect 3037 14433 3101 14497
rect 3117 14433 3181 14497
rect 3197 14433 3261 14497
rect 3277 14433 3341 14497
rect 3357 14433 3421 14497
rect 3437 14433 3501 14497
rect 3517 14433 3581 14497
rect 3597 14433 3661 14497
rect 3677 14433 3741 14497
rect 3757 14433 3821 14497
rect 3837 14433 3901 14497
rect 3917 14433 3981 14497
rect 3997 14433 4061 14497
rect 4077 14433 4141 14497
rect 4157 14433 4221 14497
rect 4237 14433 4301 14497
rect 4317 14433 4381 14497
rect 4397 14433 4461 14497
rect 4477 14433 4541 14497
rect 4557 14433 4621 14497
rect 4637 14433 4701 14497
rect 4717 14433 4781 14497
rect 4797 14433 4861 14497
rect 157 14351 221 14415
rect 237 14351 301 14415
rect 317 14351 381 14415
rect 397 14351 461 14415
rect 477 14351 541 14415
rect 557 14351 621 14415
rect 637 14351 701 14415
rect 717 14351 781 14415
rect 797 14351 861 14415
rect 877 14351 941 14415
rect 957 14351 1021 14415
rect 1037 14351 1101 14415
rect 1117 14351 1181 14415
rect 1197 14351 1261 14415
rect 1277 14351 1341 14415
rect 1357 14351 1421 14415
rect 1437 14351 1501 14415
rect 1517 14351 1581 14415
rect 1597 14351 1661 14415
rect 1677 14351 1741 14415
rect 1757 14351 1821 14415
rect 1837 14351 1901 14415
rect 1917 14351 1981 14415
rect 1997 14351 2061 14415
rect 2077 14351 2141 14415
rect 2157 14351 2221 14415
rect 2237 14351 2301 14415
rect 2317 14351 2381 14415
rect 2397 14351 2461 14415
rect 2477 14351 2541 14415
rect 2557 14351 2621 14415
rect 2637 14351 2701 14415
rect 2717 14351 2781 14415
rect 2797 14351 2861 14415
rect 2877 14351 2941 14415
rect 2957 14351 3021 14415
rect 3037 14351 3101 14415
rect 3117 14351 3181 14415
rect 3197 14351 3261 14415
rect 3277 14351 3341 14415
rect 3357 14351 3421 14415
rect 3437 14351 3501 14415
rect 3517 14351 3581 14415
rect 3597 14351 3661 14415
rect 3677 14351 3741 14415
rect 3757 14351 3821 14415
rect 3837 14351 3901 14415
rect 3917 14351 3981 14415
rect 3997 14351 4061 14415
rect 4077 14351 4141 14415
rect 4157 14351 4221 14415
rect 4237 14351 4301 14415
rect 4317 14351 4381 14415
rect 4397 14351 4461 14415
rect 4477 14351 4541 14415
rect 4557 14351 4621 14415
rect 4637 14351 4701 14415
rect 4717 14351 4781 14415
rect 4797 14351 4861 14415
rect 157 14269 221 14333
rect 237 14269 301 14333
rect 317 14269 381 14333
rect 397 14269 461 14333
rect 477 14269 541 14333
rect 557 14269 621 14333
rect 637 14269 701 14333
rect 717 14269 781 14333
rect 797 14269 861 14333
rect 877 14269 941 14333
rect 957 14269 1021 14333
rect 1037 14269 1101 14333
rect 1117 14269 1181 14333
rect 1197 14269 1261 14333
rect 1277 14269 1341 14333
rect 1357 14269 1421 14333
rect 1437 14269 1501 14333
rect 1517 14269 1581 14333
rect 1597 14269 1661 14333
rect 1677 14269 1741 14333
rect 1757 14269 1821 14333
rect 1837 14269 1901 14333
rect 1917 14269 1981 14333
rect 1997 14269 2061 14333
rect 2077 14269 2141 14333
rect 2157 14269 2221 14333
rect 2237 14269 2301 14333
rect 2317 14269 2381 14333
rect 2397 14269 2461 14333
rect 2477 14269 2541 14333
rect 2557 14269 2621 14333
rect 2637 14269 2701 14333
rect 2717 14269 2781 14333
rect 2797 14269 2861 14333
rect 2877 14269 2941 14333
rect 2957 14269 3021 14333
rect 3037 14269 3101 14333
rect 3117 14269 3181 14333
rect 3197 14269 3261 14333
rect 3277 14269 3341 14333
rect 3357 14269 3421 14333
rect 3437 14269 3501 14333
rect 3517 14269 3581 14333
rect 3597 14269 3661 14333
rect 3677 14269 3741 14333
rect 3757 14269 3821 14333
rect 3837 14269 3901 14333
rect 3917 14269 3981 14333
rect 3997 14269 4061 14333
rect 4077 14269 4141 14333
rect 4157 14269 4221 14333
rect 4237 14269 4301 14333
rect 4317 14269 4381 14333
rect 4397 14269 4461 14333
rect 4477 14269 4541 14333
rect 4557 14269 4621 14333
rect 4637 14269 4701 14333
rect 4717 14269 4781 14333
rect 4797 14269 4861 14333
rect 157 14187 221 14251
rect 237 14187 301 14251
rect 317 14187 381 14251
rect 397 14187 461 14251
rect 477 14187 541 14251
rect 557 14187 621 14251
rect 637 14187 701 14251
rect 717 14187 781 14251
rect 797 14187 861 14251
rect 877 14187 941 14251
rect 957 14187 1021 14251
rect 1037 14187 1101 14251
rect 1117 14187 1181 14251
rect 1197 14187 1261 14251
rect 1277 14187 1341 14251
rect 1357 14187 1421 14251
rect 1437 14187 1501 14251
rect 1517 14187 1581 14251
rect 1597 14187 1661 14251
rect 1677 14187 1741 14251
rect 1757 14187 1821 14251
rect 1837 14187 1901 14251
rect 1917 14187 1981 14251
rect 1997 14187 2061 14251
rect 2077 14187 2141 14251
rect 2157 14187 2221 14251
rect 2237 14187 2301 14251
rect 2317 14187 2381 14251
rect 2397 14187 2461 14251
rect 2477 14187 2541 14251
rect 2557 14187 2621 14251
rect 2637 14187 2701 14251
rect 2717 14187 2781 14251
rect 2797 14187 2861 14251
rect 2877 14187 2941 14251
rect 2957 14187 3021 14251
rect 3037 14187 3101 14251
rect 3117 14187 3181 14251
rect 3197 14187 3261 14251
rect 3277 14187 3341 14251
rect 3357 14187 3421 14251
rect 3437 14187 3501 14251
rect 3517 14187 3581 14251
rect 3597 14187 3661 14251
rect 3677 14187 3741 14251
rect 3757 14187 3821 14251
rect 3837 14187 3901 14251
rect 3917 14187 3981 14251
rect 3997 14187 4061 14251
rect 4077 14187 4141 14251
rect 4157 14187 4221 14251
rect 4237 14187 4301 14251
rect 4317 14187 4381 14251
rect 4397 14187 4461 14251
rect 4477 14187 4541 14251
rect 4557 14187 4621 14251
rect 4637 14187 4701 14251
rect 4717 14187 4781 14251
rect 4797 14187 4861 14251
rect 157 14105 221 14169
rect 237 14105 301 14169
rect 317 14105 381 14169
rect 397 14105 461 14169
rect 477 14105 541 14169
rect 557 14105 621 14169
rect 637 14105 701 14169
rect 717 14105 781 14169
rect 797 14105 861 14169
rect 877 14105 941 14169
rect 957 14105 1021 14169
rect 1037 14105 1101 14169
rect 1117 14105 1181 14169
rect 1197 14105 1261 14169
rect 1277 14105 1341 14169
rect 1357 14105 1421 14169
rect 1437 14105 1501 14169
rect 1517 14105 1581 14169
rect 1597 14105 1661 14169
rect 1677 14105 1741 14169
rect 1757 14105 1821 14169
rect 1837 14105 1901 14169
rect 1917 14105 1981 14169
rect 1997 14105 2061 14169
rect 2077 14105 2141 14169
rect 2157 14105 2221 14169
rect 2237 14105 2301 14169
rect 2317 14105 2381 14169
rect 2397 14105 2461 14169
rect 2477 14105 2541 14169
rect 2557 14105 2621 14169
rect 2637 14105 2701 14169
rect 2717 14105 2781 14169
rect 2797 14105 2861 14169
rect 2877 14105 2941 14169
rect 2957 14105 3021 14169
rect 3037 14105 3101 14169
rect 3117 14105 3181 14169
rect 3197 14105 3261 14169
rect 3277 14105 3341 14169
rect 3357 14105 3421 14169
rect 3437 14105 3501 14169
rect 3517 14105 3581 14169
rect 3597 14105 3661 14169
rect 3677 14105 3741 14169
rect 3757 14105 3821 14169
rect 3837 14105 3901 14169
rect 3917 14105 3981 14169
rect 3997 14105 4061 14169
rect 4077 14105 4141 14169
rect 4157 14105 4221 14169
rect 4237 14105 4301 14169
rect 4317 14105 4381 14169
rect 4397 14105 4461 14169
rect 4477 14105 4541 14169
rect 4557 14105 4621 14169
rect 4637 14105 4701 14169
rect 4717 14105 4781 14169
rect 4797 14105 4861 14169
rect 157 14023 221 14087
rect 237 14023 301 14087
rect 317 14023 381 14087
rect 397 14023 461 14087
rect 477 14023 541 14087
rect 557 14023 621 14087
rect 637 14023 701 14087
rect 717 14023 781 14087
rect 797 14023 861 14087
rect 877 14023 941 14087
rect 957 14023 1021 14087
rect 1037 14023 1101 14087
rect 1117 14023 1181 14087
rect 1197 14023 1261 14087
rect 1277 14023 1341 14087
rect 1357 14023 1421 14087
rect 1437 14023 1501 14087
rect 1517 14023 1581 14087
rect 1597 14023 1661 14087
rect 1677 14023 1741 14087
rect 1757 14023 1821 14087
rect 1837 14023 1901 14087
rect 1917 14023 1981 14087
rect 1997 14023 2061 14087
rect 2077 14023 2141 14087
rect 2157 14023 2221 14087
rect 2237 14023 2301 14087
rect 2317 14023 2381 14087
rect 2397 14023 2461 14087
rect 2477 14023 2541 14087
rect 2557 14023 2621 14087
rect 2637 14023 2701 14087
rect 2717 14023 2781 14087
rect 2797 14023 2861 14087
rect 2877 14023 2941 14087
rect 2957 14023 3021 14087
rect 3037 14023 3101 14087
rect 3117 14023 3181 14087
rect 3197 14023 3261 14087
rect 3277 14023 3341 14087
rect 3357 14023 3421 14087
rect 3437 14023 3501 14087
rect 3517 14023 3581 14087
rect 3597 14023 3661 14087
rect 3677 14023 3741 14087
rect 3757 14023 3821 14087
rect 3837 14023 3901 14087
rect 3917 14023 3981 14087
rect 3997 14023 4061 14087
rect 4077 14023 4141 14087
rect 4157 14023 4221 14087
rect 4237 14023 4301 14087
rect 4317 14023 4381 14087
rect 4397 14023 4461 14087
rect 4477 14023 4541 14087
rect 4557 14023 4621 14087
rect 4637 14023 4701 14087
rect 4717 14023 4781 14087
rect 4797 14023 4861 14087
rect 157 13941 221 14005
rect 237 13941 301 14005
rect 317 13941 381 14005
rect 397 13941 461 14005
rect 477 13941 541 14005
rect 557 13941 621 14005
rect 637 13941 701 14005
rect 717 13941 781 14005
rect 797 13941 861 14005
rect 877 13941 941 14005
rect 957 13941 1021 14005
rect 1037 13941 1101 14005
rect 1117 13941 1181 14005
rect 1197 13941 1261 14005
rect 1277 13941 1341 14005
rect 1357 13941 1421 14005
rect 1437 13941 1501 14005
rect 1517 13941 1581 14005
rect 1597 13941 1661 14005
rect 1677 13941 1741 14005
rect 1757 13941 1821 14005
rect 1837 13941 1901 14005
rect 1917 13941 1981 14005
rect 1997 13941 2061 14005
rect 2077 13941 2141 14005
rect 2157 13941 2221 14005
rect 2237 13941 2301 14005
rect 2317 13941 2381 14005
rect 2397 13941 2461 14005
rect 2477 13941 2541 14005
rect 2557 13941 2621 14005
rect 2637 13941 2701 14005
rect 2717 13941 2781 14005
rect 2797 13941 2861 14005
rect 2877 13941 2941 14005
rect 2957 13941 3021 14005
rect 3037 13941 3101 14005
rect 3117 13941 3181 14005
rect 3197 13941 3261 14005
rect 3277 13941 3341 14005
rect 3357 13941 3421 14005
rect 3437 13941 3501 14005
rect 3517 13941 3581 14005
rect 3597 13941 3661 14005
rect 3677 13941 3741 14005
rect 3757 13941 3821 14005
rect 3837 13941 3901 14005
rect 3917 13941 3981 14005
rect 3997 13941 4061 14005
rect 4077 13941 4141 14005
rect 4157 13941 4221 14005
rect 4237 13941 4301 14005
rect 4317 13941 4381 14005
rect 4397 13941 4461 14005
rect 4477 13941 4541 14005
rect 4557 13941 4621 14005
rect 4637 13941 4701 14005
rect 4717 13941 4781 14005
rect 4797 13941 4861 14005
rect 157 13859 221 13923
rect 237 13859 301 13923
rect 317 13859 381 13923
rect 397 13859 461 13923
rect 477 13859 541 13923
rect 557 13859 621 13923
rect 637 13859 701 13923
rect 717 13859 781 13923
rect 797 13859 861 13923
rect 877 13859 941 13923
rect 957 13859 1021 13923
rect 1037 13859 1101 13923
rect 1117 13859 1181 13923
rect 1197 13859 1261 13923
rect 1277 13859 1341 13923
rect 1357 13859 1421 13923
rect 1437 13859 1501 13923
rect 1517 13859 1581 13923
rect 1597 13859 1661 13923
rect 1677 13859 1741 13923
rect 1757 13859 1821 13923
rect 1837 13859 1901 13923
rect 1917 13859 1981 13923
rect 1997 13859 2061 13923
rect 2077 13859 2141 13923
rect 2157 13859 2221 13923
rect 2237 13859 2301 13923
rect 2317 13859 2381 13923
rect 2397 13859 2461 13923
rect 2477 13859 2541 13923
rect 2557 13859 2621 13923
rect 2637 13859 2701 13923
rect 2717 13859 2781 13923
rect 2797 13859 2861 13923
rect 2877 13859 2941 13923
rect 2957 13859 3021 13923
rect 3037 13859 3101 13923
rect 3117 13859 3181 13923
rect 3197 13859 3261 13923
rect 3277 13859 3341 13923
rect 3357 13859 3421 13923
rect 3437 13859 3501 13923
rect 3517 13859 3581 13923
rect 3597 13859 3661 13923
rect 3677 13859 3741 13923
rect 3757 13859 3821 13923
rect 3837 13859 3901 13923
rect 3917 13859 3981 13923
rect 3997 13859 4061 13923
rect 4077 13859 4141 13923
rect 4157 13859 4221 13923
rect 4237 13859 4301 13923
rect 4317 13859 4381 13923
rect 4397 13859 4461 13923
rect 4477 13859 4541 13923
rect 4557 13859 4621 13923
rect 4637 13859 4701 13923
rect 4717 13859 4781 13923
rect 4797 13859 4861 13923
rect 157 13777 221 13841
rect 237 13777 301 13841
rect 317 13777 381 13841
rect 397 13777 461 13841
rect 477 13777 541 13841
rect 557 13777 621 13841
rect 637 13777 701 13841
rect 717 13777 781 13841
rect 797 13777 861 13841
rect 877 13777 941 13841
rect 957 13777 1021 13841
rect 1037 13777 1101 13841
rect 1117 13777 1181 13841
rect 1197 13777 1261 13841
rect 1277 13777 1341 13841
rect 1357 13777 1421 13841
rect 1437 13777 1501 13841
rect 1517 13777 1581 13841
rect 1597 13777 1661 13841
rect 1677 13777 1741 13841
rect 1757 13777 1821 13841
rect 1837 13777 1901 13841
rect 1917 13777 1981 13841
rect 1997 13777 2061 13841
rect 2077 13777 2141 13841
rect 2157 13777 2221 13841
rect 2237 13777 2301 13841
rect 2317 13777 2381 13841
rect 2397 13777 2461 13841
rect 2477 13777 2541 13841
rect 2557 13777 2621 13841
rect 2637 13777 2701 13841
rect 2717 13777 2781 13841
rect 2797 13777 2861 13841
rect 2877 13777 2941 13841
rect 2957 13777 3021 13841
rect 3037 13777 3101 13841
rect 3117 13777 3181 13841
rect 3197 13777 3261 13841
rect 3277 13777 3341 13841
rect 3357 13777 3421 13841
rect 3437 13777 3501 13841
rect 3517 13777 3581 13841
rect 3597 13777 3661 13841
rect 3677 13777 3741 13841
rect 3757 13777 3821 13841
rect 3837 13777 3901 13841
rect 3917 13777 3981 13841
rect 3997 13777 4061 13841
rect 4077 13777 4141 13841
rect 4157 13777 4221 13841
rect 4237 13777 4301 13841
rect 4317 13777 4381 13841
rect 4397 13777 4461 13841
rect 4477 13777 4541 13841
rect 4557 13777 4621 13841
rect 4637 13777 4701 13841
rect 4717 13777 4781 13841
rect 4797 13777 4861 13841
rect 157 13695 221 13759
rect 237 13695 301 13759
rect 317 13695 381 13759
rect 397 13695 461 13759
rect 477 13695 541 13759
rect 557 13695 621 13759
rect 637 13695 701 13759
rect 717 13695 781 13759
rect 797 13695 861 13759
rect 877 13695 941 13759
rect 957 13695 1021 13759
rect 1037 13695 1101 13759
rect 1117 13695 1181 13759
rect 1197 13695 1261 13759
rect 1277 13695 1341 13759
rect 1357 13695 1421 13759
rect 1437 13695 1501 13759
rect 1517 13695 1581 13759
rect 1597 13695 1661 13759
rect 1677 13695 1741 13759
rect 1757 13695 1821 13759
rect 1837 13695 1901 13759
rect 1917 13695 1981 13759
rect 1997 13695 2061 13759
rect 2077 13695 2141 13759
rect 2157 13695 2221 13759
rect 2237 13695 2301 13759
rect 2317 13695 2381 13759
rect 2397 13695 2461 13759
rect 2477 13695 2541 13759
rect 2557 13695 2621 13759
rect 2637 13695 2701 13759
rect 2717 13695 2781 13759
rect 2797 13695 2861 13759
rect 2877 13695 2941 13759
rect 2957 13695 3021 13759
rect 3037 13695 3101 13759
rect 3117 13695 3181 13759
rect 3197 13695 3261 13759
rect 3277 13695 3341 13759
rect 3357 13695 3421 13759
rect 3437 13695 3501 13759
rect 3517 13695 3581 13759
rect 3597 13695 3661 13759
rect 3677 13695 3741 13759
rect 3757 13695 3821 13759
rect 3837 13695 3901 13759
rect 3917 13695 3981 13759
rect 3997 13695 4061 13759
rect 4077 13695 4141 13759
rect 4157 13695 4221 13759
rect 4237 13695 4301 13759
rect 4317 13695 4381 13759
rect 4397 13695 4461 13759
rect 4477 13695 4541 13759
rect 4557 13695 4621 13759
rect 4637 13695 4701 13759
rect 4717 13695 4781 13759
rect 4797 13695 4861 13759
rect 157 13613 221 13677
rect 237 13613 301 13677
rect 317 13613 381 13677
rect 397 13613 461 13677
rect 477 13613 541 13677
rect 557 13613 621 13677
rect 637 13613 701 13677
rect 717 13613 781 13677
rect 797 13613 861 13677
rect 877 13613 941 13677
rect 957 13613 1021 13677
rect 1037 13613 1101 13677
rect 1117 13613 1181 13677
rect 1197 13613 1261 13677
rect 1277 13613 1341 13677
rect 1357 13613 1421 13677
rect 1437 13613 1501 13677
rect 1517 13613 1581 13677
rect 1597 13613 1661 13677
rect 1677 13613 1741 13677
rect 1757 13613 1821 13677
rect 1837 13613 1901 13677
rect 1917 13613 1981 13677
rect 1997 13613 2061 13677
rect 2077 13613 2141 13677
rect 2157 13613 2221 13677
rect 2237 13613 2301 13677
rect 2317 13613 2381 13677
rect 2397 13613 2461 13677
rect 2477 13613 2541 13677
rect 2557 13613 2621 13677
rect 2637 13613 2701 13677
rect 2717 13613 2781 13677
rect 2797 13613 2861 13677
rect 2877 13613 2941 13677
rect 2957 13613 3021 13677
rect 3037 13613 3101 13677
rect 3117 13613 3181 13677
rect 3197 13613 3261 13677
rect 3277 13613 3341 13677
rect 3357 13613 3421 13677
rect 3437 13613 3501 13677
rect 3517 13613 3581 13677
rect 3597 13613 3661 13677
rect 3677 13613 3741 13677
rect 3757 13613 3821 13677
rect 3837 13613 3901 13677
rect 3917 13613 3981 13677
rect 3997 13613 4061 13677
rect 4077 13613 4141 13677
rect 4157 13613 4221 13677
rect 4237 13613 4301 13677
rect 4317 13613 4381 13677
rect 4397 13613 4461 13677
rect 4477 13613 4541 13677
rect 4557 13613 4621 13677
rect 4637 13613 4701 13677
rect 4717 13613 4781 13677
rect 4797 13613 4861 13677
rect 10190 16460 10254 16524
rect 10270 16460 10334 16524
rect 10350 16460 10414 16524
rect 10430 16460 10494 16524
rect 10510 16460 10574 16524
rect 10590 16460 10654 16524
rect 10670 16460 10734 16524
rect 10750 16460 10814 16524
rect 10830 16460 10894 16524
rect 10910 16460 10974 16524
rect 10990 16460 11054 16524
rect 11070 16460 11134 16524
rect 11150 16460 11214 16524
rect 11230 16460 11294 16524
rect 11310 16460 11374 16524
rect 11390 16460 11454 16524
rect 11470 16460 11534 16524
rect 11550 16460 11614 16524
rect 11630 16460 11694 16524
rect 11710 16460 11774 16524
rect 11790 16460 11854 16524
rect 11870 16460 11934 16524
rect 11950 16460 12014 16524
rect 12030 16460 12094 16524
rect 12110 16460 12174 16524
rect 12190 16460 12254 16524
rect 12270 16460 12334 16524
rect 12350 16460 12414 16524
rect 12430 16460 12494 16524
rect 12510 16460 12574 16524
rect 12590 16460 12654 16524
rect 12670 16460 12734 16524
rect 12750 16460 12814 16524
rect 12830 16460 12894 16524
rect 12910 16460 12974 16524
rect 12990 16460 13054 16524
rect 13070 16460 13134 16524
rect 13150 16460 13214 16524
rect 13230 16460 13294 16524
rect 13310 16460 13374 16524
rect 13390 16460 13454 16524
rect 13470 16460 13534 16524
rect 13550 16460 13614 16524
rect 13630 16460 13694 16524
rect 13710 16460 13774 16524
rect 13790 16460 13854 16524
rect 13870 16460 13934 16524
rect 13950 16460 14014 16524
rect 14030 16460 14094 16524
rect 14110 16460 14174 16524
rect 14190 16460 14254 16524
rect 14270 16460 14334 16524
rect 14350 16460 14414 16524
rect 14430 16460 14494 16524
rect 14510 16460 14574 16524
rect 14590 16460 14654 16524
rect 14670 16460 14734 16524
rect 14750 16460 14814 16524
rect 14830 16460 14894 16524
rect 10190 16379 10254 16443
rect 10270 16379 10334 16443
rect 10350 16379 10414 16443
rect 10430 16379 10494 16443
rect 10510 16379 10574 16443
rect 10590 16379 10654 16443
rect 10670 16379 10734 16443
rect 10750 16379 10814 16443
rect 10830 16379 10894 16443
rect 10910 16379 10974 16443
rect 10990 16379 11054 16443
rect 11070 16379 11134 16443
rect 11150 16379 11214 16443
rect 11230 16379 11294 16443
rect 11310 16379 11374 16443
rect 11390 16379 11454 16443
rect 11470 16379 11534 16443
rect 11550 16379 11614 16443
rect 11630 16379 11694 16443
rect 11710 16379 11774 16443
rect 11790 16379 11854 16443
rect 11870 16379 11934 16443
rect 11950 16379 12014 16443
rect 12030 16379 12094 16443
rect 12110 16379 12174 16443
rect 12190 16379 12254 16443
rect 12270 16379 12334 16443
rect 12350 16379 12414 16443
rect 12430 16379 12494 16443
rect 12510 16379 12574 16443
rect 12590 16379 12654 16443
rect 12670 16379 12734 16443
rect 12750 16379 12814 16443
rect 12830 16379 12894 16443
rect 12910 16379 12974 16443
rect 12990 16379 13054 16443
rect 13070 16379 13134 16443
rect 13150 16379 13214 16443
rect 13230 16379 13294 16443
rect 13310 16379 13374 16443
rect 13390 16379 13454 16443
rect 13470 16379 13534 16443
rect 13550 16379 13614 16443
rect 13630 16379 13694 16443
rect 13710 16379 13774 16443
rect 13790 16379 13854 16443
rect 13870 16379 13934 16443
rect 13950 16379 14014 16443
rect 14030 16379 14094 16443
rect 14110 16379 14174 16443
rect 14190 16379 14254 16443
rect 14270 16379 14334 16443
rect 14350 16379 14414 16443
rect 14430 16379 14494 16443
rect 14510 16379 14574 16443
rect 14590 16379 14654 16443
rect 14670 16379 14734 16443
rect 14750 16379 14814 16443
rect 14830 16379 14894 16443
rect 10190 16298 10254 16362
rect 10270 16298 10334 16362
rect 10350 16298 10414 16362
rect 10430 16298 10494 16362
rect 10510 16298 10574 16362
rect 10590 16298 10654 16362
rect 10670 16298 10734 16362
rect 10750 16298 10814 16362
rect 10830 16298 10894 16362
rect 10910 16298 10974 16362
rect 10990 16298 11054 16362
rect 11070 16298 11134 16362
rect 11150 16298 11214 16362
rect 11230 16298 11294 16362
rect 11310 16298 11374 16362
rect 11390 16298 11454 16362
rect 11470 16298 11534 16362
rect 11550 16298 11614 16362
rect 11630 16298 11694 16362
rect 11710 16298 11774 16362
rect 11790 16298 11854 16362
rect 11870 16298 11934 16362
rect 11950 16298 12014 16362
rect 12030 16298 12094 16362
rect 12110 16298 12174 16362
rect 12190 16298 12254 16362
rect 12270 16298 12334 16362
rect 12350 16298 12414 16362
rect 12430 16298 12494 16362
rect 12510 16298 12574 16362
rect 12590 16298 12654 16362
rect 12670 16298 12734 16362
rect 12750 16298 12814 16362
rect 12830 16298 12894 16362
rect 12910 16298 12974 16362
rect 12990 16298 13054 16362
rect 13070 16298 13134 16362
rect 13150 16298 13214 16362
rect 13230 16298 13294 16362
rect 13310 16298 13374 16362
rect 13390 16298 13454 16362
rect 13470 16298 13534 16362
rect 13550 16298 13614 16362
rect 13630 16298 13694 16362
rect 13710 16298 13774 16362
rect 13790 16298 13854 16362
rect 13870 16298 13934 16362
rect 13950 16298 14014 16362
rect 14030 16298 14094 16362
rect 14110 16298 14174 16362
rect 14190 16298 14254 16362
rect 14270 16298 14334 16362
rect 14350 16298 14414 16362
rect 14430 16298 14494 16362
rect 14510 16298 14574 16362
rect 14590 16298 14654 16362
rect 14670 16298 14734 16362
rect 14750 16298 14814 16362
rect 14830 16298 14894 16362
rect 10190 16217 10254 16281
rect 10270 16217 10334 16281
rect 10350 16217 10414 16281
rect 10430 16217 10494 16281
rect 10510 16217 10574 16281
rect 10590 16217 10654 16281
rect 10670 16217 10734 16281
rect 10750 16217 10814 16281
rect 10830 16217 10894 16281
rect 10910 16217 10974 16281
rect 10990 16217 11054 16281
rect 11070 16217 11134 16281
rect 11150 16217 11214 16281
rect 11230 16217 11294 16281
rect 11310 16217 11374 16281
rect 11390 16217 11454 16281
rect 11470 16217 11534 16281
rect 11550 16217 11614 16281
rect 11630 16217 11694 16281
rect 11710 16217 11774 16281
rect 11790 16217 11854 16281
rect 11870 16217 11934 16281
rect 11950 16217 12014 16281
rect 12030 16217 12094 16281
rect 12110 16217 12174 16281
rect 12190 16217 12254 16281
rect 12270 16217 12334 16281
rect 12350 16217 12414 16281
rect 12430 16217 12494 16281
rect 12510 16217 12574 16281
rect 12590 16217 12654 16281
rect 12670 16217 12734 16281
rect 12750 16217 12814 16281
rect 12830 16217 12894 16281
rect 12910 16217 12974 16281
rect 12990 16217 13054 16281
rect 13070 16217 13134 16281
rect 13150 16217 13214 16281
rect 13230 16217 13294 16281
rect 13310 16217 13374 16281
rect 13390 16217 13454 16281
rect 13470 16217 13534 16281
rect 13550 16217 13614 16281
rect 13630 16217 13694 16281
rect 13710 16217 13774 16281
rect 13790 16217 13854 16281
rect 13870 16217 13934 16281
rect 13950 16217 14014 16281
rect 14030 16217 14094 16281
rect 14110 16217 14174 16281
rect 14190 16217 14254 16281
rect 14270 16217 14334 16281
rect 14350 16217 14414 16281
rect 14430 16217 14494 16281
rect 14510 16217 14574 16281
rect 14590 16217 14654 16281
rect 14670 16217 14734 16281
rect 14750 16217 14814 16281
rect 14830 16217 14894 16281
rect 10190 16136 10254 16200
rect 10270 16136 10334 16200
rect 10350 16136 10414 16200
rect 10430 16136 10494 16200
rect 10510 16136 10574 16200
rect 10590 16136 10654 16200
rect 10670 16136 10734 16200
rect 10750 16136 10814 16200
rect 10830 16136 10894 16200
rect 10910 16136 10974 16200
rect 10990 16136 11054 16200
rect 11070 16136 11134 16200
rect 11150 16136 11214 16200
rect 11230 16136 11294 16200
rect 11310 16136 11374 16200
rect 11390 16136 11454 16200
rect 11470 16136 11534 16200
rect 11550 16136 11614 16200
rect 11630 16136 11694 16200
rect 11710 16136 11774 16200
rect 11790 16136 11854 16200
rect 11870 16136 11934 16200
rect 11950 16136 12014 16200
rect 12030 16136 12094 16200
rect 12110 16136 12174 16200
rect 12190 16136 12254 16200
rect 12270 16136 12334 16200
rect 12350 16136 12414 16200
rect 12430 16136 12494 16200
rect 12510 16136 12574 16200
rect 12590 16136 12654 16200
rect 12670 16136 12734 16200
rect 12750 16136 12814 16200
rect 12830 16136 12894 16200
rect 12910 16136 12974 16200
rect 12990 16136 13054 16200
rect 13070 16136 13134 16200
rect 13150 16136 13214 16200
rect 13230 16136 13294 16200
rect 13310 16136 13374 16200
rect 13390 16136 13454 16200
rect 13470 16136 13534 16200
rect 13550 16136 13614 16200
rect 13630 16136 13694 16200
rect 13710 16136 13774 16200
rect 13790 16136 13854 16200
rect 13870 16136 13934 16200
rect 13950 16136 14014 16200
rect 14030 16136 14094 16200
rect 14110 16136 14174 16200
rect 14190 16136 14254 16200
rect 14270 16136 14334 16200
rect 14350 16136 14414 16200
rect 14430 16136 14494 16200
rect 14510 16136 14574 16200
rect 14590 16136 14654 16200
rect 14670 16136 14734 16200
rect 14750 16136 14814 16200
rect 14830 16136 14894 16200
rect 10190 16055 10254 16119
rect 10270 16055 10334 16119
rect 10350 16055 10414 16119
rect 10430 16055 10494 16119
rect 10510 16055 10574 16119
rect 10590 16055 10654 16119
rect 10670 16055 10734 16119
rect 10750 16055 10814 16119
rect 10830 16055 10894 16119
rect 10910 16055 10974 16119
rect 10990 16055 11054 16119
rect 11070 16055 11134 16119
rect 11150 16055 11214 16119
rect 11230 16055 11294 16119
rect 11310 16055 11374 16119
rect 11390 16055 11454 16119
rect 11470 16055 11534 16119
rect 11550 16055 11614 16119
rect 11630 16055 11694 16119
rect 11710 16055 11774 16119
rect 11790 16055 11854 16119
rect 11870 16055 11934 16119
rect 11950 16055 12014 16119
rect 12030 16055 12094 16119
rect 12110 16055 12174 16119
rect 12190 16055 12254 16119
rect 12270 16055 12334 16119
rect 12350 16055 12414 16119
rect 12430 16055 12494 16119
rect 12510 16055 12574 16119
rect 12590 16055 12654 16119
rect 12670 16055 12734 16119
rect 12750 16055 12814 16119
rect 12830 16055 12894 16119
rect 12910 16055 12974 16119
rect 12990 16055 13054 16119
rect 13070 16055 13134 16119
rect 13150 16055 13214 16119
rect 13230 16055 13294 16119
rect 13310 16055 13374 16119
rect 13390 16055 13454 16119
rect 13470 16055 13534 16119
rect 13550 16055 13614 16119
rect 13630 16055 13694 16119
rect 13710 16055 13774 16119
rect 13790 16055 13854 16119
rect 13870 16055 13934 16119
rect 13950 16055 14014 16119
rect 14030 16055 14094 16119
rect 14110 16055 14174 16119
rect 14190 16055 14254 16119
rect 14270 16055 14334 16119
rect 14350 16055 14414 16119
rect 14430 16055 14494 16119
rect 14510 16055 14574 16119
rect 14590 16055 14654 16119
rect 14670 16055 14734 16119
rect 14750 16055 14814 16119
rect 14830 16055 14894 16119
rect 10190 15974 10254 16038
rect 10270 15974 10334 16038
rect 10350 15974 10414 16038
rect 10430 15974 10494 16038
rect 10510 15974 10574 16038
rect 10590 15974 10654 16038
rect 10670 15974 10734 16038
rect 10750 15974 10814 16038
rect 10830 15974 10894 16038
rect 10910 15974 10974 16038
rect 10990 15974 11054 16038
rect 11070 15974 11134 16038
rect 11150 15974 11214 16038
rect 11230 15974 11294 16038
rect 11310 15974 11374 16038
rect 11390 15974 11454 16038
rect 11470 15974 11534 16038
rect 11550 15974 11614 16038
rect 11630 15974 11694 16038
rect 11710 15974 11774 16038
rect 11790 15974 11854 16038
rect 11870 15974 11934 16038
rect 11950 15974 12014 16038
rect 12030 15974 12094 16038
rect 12110 15974 12174 16038
rect 12190 15974 12254 16038
rect 12270 15974 12334 16038
rect 12350 15974 12414 16038
rect 12430 15974 12494 16038
rect 12510 15974 12574 16038
rect 12590 15974 12654 16038
rect 12670 15974 12734 16038
rect 12750 15974 12814 16038
rect 12830 15974 12894 16038
rect 12910 15974 12974 16038
rect 12990 15974 13054 16038
rect 13070 15974 13134 16038
rect 13150 15974 13214 16038
rect 13230 15974 13294 16038
rect 13310 15974 13374 16038
rect 13390 15974 13454 16038
rect 13470 15974 13534 16038
rect 13550 15974 13614 16038
rect 13630 15974 13694 16038
rect 13710 15974 13774 16038
rect 13790 15974 13854 16038
rect 13870 15974 13934 16038
rect 13950 15974 14014 16038
rect 14030 15974 14094 16038
rect 14110 15974 14174 16038
rect 14190 15974 14254 16038
rect 14270 15974 14334 16038
rect 14350 15974 14414 16038
rect 14430 15974 14494 16038
rect 14510 15974 14574 16038
rect 14590 15974 14654 16038
rect 14670 15974 14734 16038
rect 14750 15974 14814 16038
rect 14830 15974 14894 16038
rect 10190 15893 10254 15957
rect 10270 15893 10334 15957
rect 10350 15893 10414 15957
rect 10430 15893 10494 15957
rect 10510 15893 10574 15957
rect 10590 15893 10654 15957
rect 10670 15893 10734 15957
rect 10750 15893 10814 15957
rect 10830 15893 10894 15957
rect 10910 15893 10974 15957
rect 10990 15893 11054 15957
rect 11070 15893 11134 15957
rect 11150 15893 11214 15957
rect 11230 15893 11294 15957
rect 11310 15893 11374 15957
rect 11390 15893 11454 15957
rect 11470 15893 11534 15957
rect 11550 15893 11614 15957
rect 11630 15893 11694 15957
rect 11710 15893 11774 15957
rect 11790 15893 11854 15957
rect 11870 15893 11934 15957
rect 11950 15893 12014 15957
rect 12030 15893 12094 15957
rect 12110 15893 12174 15957
rect 12190 15893 12254 15957
rect 12270 15893 12334 15957
rect 12350 15893 12414 15957
rect 12430 15893 12494 15957
rect 12510 15893 12574 15957
rect 12590 15893 12654 15957
rect 12670 15893 12734 15957
rect 12750 15893 12814 15957
rect 12830 15893 12894 15957
rect 12910 15893 12974 15957
rect 12990 15893 13054 15957
rect 13070 15893 13134 15957
rect 13150 15893 13214 15957
rect 13230 15893 13294 15957
rect 13310 15893 13374 15957
rect 13390 15893 13454 15957
rect 13470 15893 13534 15957
rect 13550 15893 13614 15957
rect 13630 15893 13694 15957
rect 13710 15893 13774 15957
rect 13790 15893 13854 15957
rect 13870 15893 13934 15957
rect 13950 15893 14014 15957
rect 14030 15893 14094 15957
rect 14110 15893 14174 15957
rect 14190 15893 14254 15957
rect 14270 15893 14334 15957
rect 14350 15893 14414 15957
rect 14430 15893 14494 15957
rect 14510 15893 14574 15957
rect 14590 15893 14654 15957
rect 14670 15893 14734 15957
rect 14750 15893 14814 15957
rect 14830 15893 14894 15957
rect 10190 15812 10254 15876
rect 10270 15812 10334 15876
rect 10350 15812 10414 15876
rect 10430 15812 10494 15876
rect 10510 15812 10574 15876
rect 10590 15812 10654 15876
rect 10670 15812 10734 15876
rect 10750 15812 10814 15876
rect 10830 15812 10894 15876
rect 10910 15812 10974 15876
rect 10990 15812 11054 15876
rect 11070 15812 11134 15876
rect 11150 15812 11214 15876
rect 11230 15812 11294 15876
rect 11310 15812 11374 15876
rect 11390 15812 11454 15876
rect 11470 15812 11534 15876
rect 11550 15812 11614 15876
rect 11630 15812 11694 15876
rect 11710 15812 11774 15876
rect 11790 15812 11854 15876
rect 11870 15812 11934 15876
rect 11950 15812 12014 15876
rect 12030 15812 12094 15876
rect 12110 15812 12174 15876
rect 12190 15812 12254 15876
rect 12270 15812 12334 15876
rect 12350 15812 12414 15876
rect 12430 15812 12494 15876
rect 12510 15812 12574 15876
rect 12590 15812 12654 15876
rect 12670 15812 12734 15876
rect 12750 15812 12814 15876
rect 12830 15812 12894 15876
rect 12910 15812 12974 15876
rect 12990 15812 13054 15876
rect 13070 15812 13134 15876
rect 13150 15812 13214 15876
rect 13230 15812 13294 15876
rect 13310 15812 13374 15876
rect 13390 15812 13454 15876
rect 13470 15812 13534 15876
rect 13550 15812 13614 15876
rect 13630 15812 13694 15876
rect 13710 15812 13774 15876
rect 13790 15812 13854 15876
rect 13870 15812 13934 15876
rect 13950 15812 14014 15876
rect 14030 15812 14094 15876
rect 14110 15812 14174 15876
rect 14190 15812 14254 15876
rect 14270 15812 14334 15876
rect 14350 15812 14414 15876
rect 14430 15812 14494 15876
rect 14510 15812 14574 15876
rect 14590 15812 14654 15876
rect 14670 15812 14734 15876
rect 14750 15812 14814 15876
rect 14830 15812 14894 15876
rect 10190 15731 10254 15795
rect 10270 15731 10334 15795
rect 10350 15731 10414 15795
rect 10430 15731 10494 15795
rect 10510 15731 10574 15795
rect 10590 15731 10654 15795
rect 10670 15731 10734 15795
rect 10750 15731 10814 15795
rect 10830 15731 10894 15795
rect 10910 15731 10974 15795
rect 10990 15731 11054 15795
rect 11070 15731 11134 15795
rect 11150 15731 11214 15795
rect 11230 15731 11294 15795
rect 11310 15731 11374 15795
rect 11390 15731 11454 15795
rect 11470 15731 11534 15795
rect 11550 15731 11614 15795
rect 11630 15731 11694 15795
rect 11710 15731 11774 15795
rect 11790 15731 11854 15795
rect 11870 15731 11934 15795
rect 11950 15731 12014 15795
rect 12030 15731 12094 15795
rect 12110 15731 12174 15795
rect 12190 15731 12254 15795
rect 12270 15731 12334 15795
rect 12350 15731 12414 15795
rect 12430 15731 12494 15795
rect 12510 15731 12574 15795
rect 12590 15731 12654 15795
rect 12670 15731 12734 15795
rect 12750 15731 12814 15795
rect 12830 15731 12894 15795
rect 12910 15731 12974 15795
rect 12990 15731 13054 15795
rect 13070 15731 13134 15795
rect 13150 15731 13214 15795
rect 13230 15731 13294 15795
rect 13310 15731 13374 15795
rect 13390 15731 13454 15795
rect 13470 15731 13534 15795
rect 13550 15731 13614 15795
rect 13630 15731 13694 15795
rect 13710 15731 13774 15795
rect 13790 15731 13854 15795
rect 13870 15731 13934 15795
rect 13950 15731 14014 15795
rect 14030 15731 14094 15795
rect 14110 15731 14174 15795
rect 14190 15731 14254 15795
rect 14270 15731 14334 15795
rect 14350 15731 14414 15795
rect 14430 15731 14494 15795
rect 14510 15731 14574 15795
rect 14590 15731 14654 15795
rect 14670 15731 14734 15795
rect 14750 15731 14814 15795
rect 14830 15731 14894 15795
rect 10190 15650 10254 15714
rect 10270 15650 10334 15714
rect 10350 15650 10414 15714
rect 10430 15650 10494 15714
rect 10510 15650 10574 15714
rect 10590 15650 10654 15714
rect 10670 15650 10734 15714
rect 10750 15650 10814 15714
rect 10830 15650 10894 15714
rect 10910 15650 10974 15714
rect 10990 15650 11054 15714
rect 11070 15650 11134 15714
rect 11150 15650 11214 15714
rect 11230 15650 11294 15714
rect 11310 15650 11374 15714
rect 11390 15650 11454 15714
rect 11470 15650 11534 15714
rect 11550 15650 11614 15714
rect 11630 15650 11694 15714
rect 11710 15650 11774 15714
rect 11790 15650 11854 15714
rect 11870 15650 11934 15714
rect 11950 15650 12014 15714
rect 12030 15650 12094 15714
rect 12110 15650 12174 15714
rect 12190 15650 12254 15714
rect 12270 15650 12334 15714
rect 12350 15650 12414 15714
rect 12430 15650 12494 15714
rect 12510 15650 12574 15714
rect 12590 15650 12654 15714
rect 12670 15650 12734 15714
rect 12750 15650 12814 15714
rect 12830 15650 12894 15714
rect 12910 15650 12974 15714
rect 12990 15650 13054 15714
rect 13070 15650 13134 15714
rect 13150 15650 13214 15714
rect 13230 15650 13294 15714
rect 13310 15650 13374 15714
rect 13390 15650 13454 15714
rect 13470 15650 13534 15714
rect 13550 15650 13614 15714
rect 13630 15650 13694 15714
rect 13710 15650 13774 15714
rect 13790 15650 13854 15714
rect 13870 15650 13934 15714
rect 13950 15650 14014 15714
rect 14030 15650 14094 15714
rect 14110 15650 14174 15714
rect 14190 15650 14254 15714
rect 14270 15650 14334 15714
rect 14350 15650 14414 15714
rect 14430 15650 14494 15714
rect 14510 15650 14574 15714
rect 14590 15650 14654 15714
rect 14670 15650 14734 15714
rect 14750 15650 14814 15714
rect 14830 15650 14894 15714
rect 10190 15569 10254 15633
rect 10270 15569 10334 15633
rect 10350 15569 10414 15633
rect 10430 15569 10494 15633
rect 10510 15569 10574 15633
rect 10590 15569 10654 15633
rect 10670 15569 10734 15633
rect 10750 15569 10814 15633
rect 10830 15569 10894 15633
rect 10910 15569 10974 15633
rect 10990 15569 11054 15633
rect 11070 15569 11134 15633
rect 11150 15569 11214 15633
rect 11230 15569 11294 15633
rect 11310 15569 11374 15633
rect 11390 15569 11454 15633
rect 11470 15569 11534 15633
rect 11550 15569 11614 15633
rect 11630 15569 11694 15633
rect 11710 15569 11774 15633
rect 11790 15569 11854 15633
rect 11870 15569 11934 15633
rect 11950 15569 12014 15633
rect 12030 15569 12094 15633
rect 12110 15569 12174 15633
rect 12190 15569 12254 15633
rect 12270 15569 12334 15633
rect 12350 15569 12414 15633
rect 12430 15569 12494 15633
rect 12510 15569 12574 15633
rect 12590 15569 12654 15633
rect 12670 15569 12734 15633
rect 12750 15569 12814 15633
rect 12830 15569 12894 15633
rect 12910 15569 12974 15633
rect 12990 15569 13054 15633
rect 13070 15569 13134 15633
rect 13150 15569 13214 15633
rect 13230 15569 13294 15633
rect 13310 15569 13374 15633
rect 13390 15569 13454 15633
rect 13470 15569 13534 15633
rect 13550 15569 13614 15633
rect 13630 15569 13694 15633
rect 13710 15569 13774 15633
rect 13790 15569 13854 15633
rect 13870 15569 13934 15633
rect 13950 15569 14014 15633
rect 14030 15569 14094 15633
rect 14110 15569 14174 15633
rect 14190 15569 14254 15633
rect 14270 15569 14334 15633
rect 14350 15569 14414 15633
rect 14430 15569 14494 15633
rect 14510 15569 14574 15633
rect 14590 15569 14654 15633
rect 14670 15569 14734 15633
rect 14750 15569 14814 15633
rect 14830 15569 14894 15633
rect 10190 15488 10254 15552
rect 10270 15488 10334 15552
rect 10350 15488 10414 15552
rect 10430 15488 10494 15552
rect 10510 15488 10574 15552
rect 10590 15488 10654 15552
rect 10670 15488 10734 15552
rect 10750 15488 10814 15552
rect 10830 15488 10894 15552
rect 10910 15488 10974 15552
rect 10990 15488 11054 15552
rect 11070 15488 11134 15552
rect 11150 15488 11214 15552
rect 11230 15488 11294 15552
rect 11310 15488 11374 15552
rect 11390 15488 11454 15552
rect 11470 15488 11534 15552
rect 11550 15488 11614 15552
rect 11630 15488 11694 15552
rect 11710 15488 11774 15552
rect 11790 15488 11854 15552
rect 11870 15488 11934 15552
rect 11950 15488 12014 15552
rect 12030 15488 12094 15552
rect 12110 15488 12174 15552
rect 12190 15488 12254 15552
rect 12270 15488 12334 15552
rect 12350 15488 12414 15552
rect 12430 15488 12494 15552
rect 12510 15488 12574 15552
rect 12590 15488 12654 15552
rect 12670 15488 12734 15552
rect 12750 15488 12814 15552
rect 12830 15488 12894 15552
rect 12910 15488 12974 15552
rect 12990 15488 13054 15552
rect 13070 15488 13134 15552
rect 13150 15488 13214 15552
rect 13230 15488 13294 15552
rect 13310 15488 13374 15552
rect 13390 15488 13454 15552
rect 13470 15488 13534 15552
rect 13550 15488 13614 15552
rect 13630 15488 13694 15552
rect 13710 15488 13774 15552
rect 13790 15488 13854 15552
rect 13870 15488 13934 15552
rect 13950 15488 14014 15552
rect 14030 15488 14094 15552
rect 14110 15488 14174 15552
rect 14190 15488 14254 15552
rect 14270 15488 14334 15552
rect 14350 15488 14414 15552
rect 14430 15488 14494 15552
rect 14510 15488 14574 15552
rect 14590 15488 14654 15552
rect 14670 15488 14734 15552
rect 14750 15488 14814 15552
rect 14830 15488 14894 15552
rect 10190 15407 10254 15471
rect 10270 15407 10334 15471
rect 10350 15407 10414 15471
rect 10430 15407 10494 15471
rect 10510 15407 10574 15471
rect 10590 15407 10654 15471
rect 10670 15407 10734 15471
rect 10750 15407 10814 15471
rect 10830 15407 10894 15471
rect 10910 15407 10974 15471
rect 10990 15407 11054 15471
rect 11070 15407 11134 15471
rect 11150 15407 11214 15471
rect 11230 15407 11294 15471
rect 11310 15407 11374 15471
rect 11390 15407 11454 15471
rect 11470 15407 11534 15471
rect 11550 15407 11614 15471
rect 11630 15407 11694 15471
rect 11710 15407 11774 15471
rect 11790 15407 11854 15471
rect 11870 15407 11934 15471
rect 11950 15407 12014 15471
rect 12030 15407 12094 15471
rect 12110 15407 12174 15471
rect 12190 15407 12254 15471
rect 12270 15407 12334 15471
rect 12350 15407 12414 15471
rect 12430 15407 12494 15471
rect 12510 15407 12574 15471
rect 12590 15407 12654 15471
rect 12670 15407 12734 15471
rect 12750 15407 12814 15471
rect 12830 15407 12894 15471
rect 12910 15407 12974 15471
rect 12990 15407 13054 15471
rect 13070 15407 13134 15471
rect 13150 15407 13214 15471
rect 13230 15407 13294 15471
rect 13310 15407 13374 15471
rect 13390 15407 13454 15471
rect 13470 15407 13534 15471
rect 13550 15407 13614 15471
rect 13630 15407 13694 15471
rect 13710 15407 13774 15471
rect 13790 15407 13854 15471
rect 13870 15407 13934 15471
rect 13950 15407 14014 15471
rect 14030 15407 14094 15471
rect 14110 15407 14174 15471
rect 14190 15407 14254 15471
rect 14270 15407 14334 15471
rect 14350 15407 14414 15471
rect 14430 15407 14494 15471
rect 14510 15407 14574 15471
rect 14590 15407 14654 15471
rect 14670 15407 14734 15471
rect 14750 15407 14814 15471
rect 14830 15407 14894 15471
rect 10190 15326 10254 15390
rect 10270 15326 10334 15390
rect 10350 15326 10414 15390
rect 10430 15326 10494 15390
rect 10510 15326 10574 15390
rect 10590 15326 10654 15390
rect 10670 15326 10734 15390
rect 10750 15326 10814 15390
rect 10830 15326 10894 15390
rect 10910 15326 10974 15390
rect 10990 15326 11054 15390
rect 11070 15326 11134 15390
rect 11150 15326 11214 15390
rect 11230 15326 11294 15390
rect 11310 15326 11374 15390
rect 11390 15326 11454 15390
rect 11470 15326 11534 15390
rect 11550 15326 11614 15390
rect 11630 15326 11694 15390
rect 11710 15326 11774 15390
rect 11790 15326 11854 15390
rect 11870 15326 11934 15390
rect 11950 15326 12014 15390
rect 12030 15326 12094 15390
rect 12110 15326 12174 15390
rect 12190 15326 12254 15390
rect 12270 15326 12334 15390
rect 12350 15326 12414 15390
rect 12430 15326 12494 15390
rect 12510 15326 12574 15390
rect 12590 15326 12654 15390
rect 12670 15326 12734 15390
rect 12750 15326 12814 15390
rect 12830 15326 12894 15390
rect 12910 15326 12974 15390
rect 12990 15326 13054 15390
rect 13070 15326 13134 15390
rect 13150 15326 13214 15390
rect 13230 15326 13294 15390
rect 13310 15326 13374 15390
rect 13390 15326 13454 15390
rect 13470 15326 13534 15390
rect 13550 15326 13614 15390
rect 13630 15326 13694 15390
rect 13710 15326 13774 15390
rect 13790 15326 13854 15390
rect 13870 15326 13934 15390
rect 13950 15326 14014 15390
rect 14030 15326 14094 15390
rect 14110 15326 14174 15390
rect 14190 15326 14254 15390
rect 14270 15326 14334 15390
rect 14350 15326 14414 15390
rect 14430 15326 14494 15390
rect 14510 15326 14574 15390
rect 14590 15326 14654 15390
rect 14670 15326 14734 15390
rect 14750 15326 14814 15390
rect 14830 15326 14894 15390
rect 10190 15245 10254 15309
rect 10270 15245 10334 15309
rect 10350 15245 10414 15309
rect 10430 15245 10494 15309
rect 10510 15245 10574 15309
rect 10590 15245 10654 15309
rect 10670 15245 10734 15309
rect 10750 15245 10814 15309
rect 10830 15245 10894 15309
rect 10910 15245 10974 15309
rect 10990 15245 11054 15309
rect 11070 15245 11134 15309
rect 11150 15245 11214 15309
rect 11230 15245 11294 15309
rect 11310 15245 11374 15309
rect 11390 15245 11454 15309
rect 11470 15245 11534 15309
rect 11550 15245 11614 15309
rect 11630 15245 11694 15309
rect 11710 15245 11774 15309
rect 11790 15245 11854 15309
rect 11870 15245 11934 15309
rect 11950 15245 12014 15309
rect 12030 15245 12094 15309
rect 12110 15245 12174 15309
rect 12190 15245 12254 15309
rect 12270 15245 12334 15309
rect 12350 15245 12414 15309
rect 12430 15245 12494 15309
rect 12510 15245 12574 15309
rect 12590 15245 12654 15309
rect 12670 15245 12734 15309
rect 12750 15245 12814 15309
rect 12830 15245 12894 15309
rect 12910 15245 12974 15309
rect 12990 15245 13054 15309
rect 13070 15245 13134 15309
rect 13150 15245 13214 15309
rect 13230 15245 13294 15309
rect 13310 15245 13374 15309
rect 13390 15245 13454 15309
rect 13470 15245 13534 15309
rect 13550 15245 13614 15309
rect 13630 15245 13694 15309
rect 13710 15245 13774 15309
rect 13790 15245 13854 15309
rect 13870 15245 13934 15309
rect 13950 15245 14014 15309
rect 14030 15245 14094 15309
rect 14110 15245 14174 15309
rect 14190 15245 14254 15309
rect 14270 15245 14334 15309
rect 14350 15245 14414 15309
rect 14430 15245 14494 15309
rect 14510 15245 14574 15309
rect 14590 15245 14654 15309
rect 14670 15245 14734 15309
rect 14750 15245 14814 15309
rect 14830 15245 14894 15309
rect 10190 15164 10254 15228
rect 10270 15164 10334 15228
rect 10350 15164 10414 15228
rect 10430 15164 10494 15228
rect 10510 15164 10574 15228
rect 10590 15164 10654 15228
rect 10670 15164 10734 15228
rect 10750 15164 10814 15228
rect 10830 15164 10894 15228
rect 10910 15164 10974 15228
rect 10990 15164 11054 15228
rect 11070 15164 11134 15228
rect 11150 15164 11214 15228
rect 11230 15164 11294 15228
rect 11310 15164 11374 15228
rect 11390 15164 11454 15228
rect 11470 15164 11534 15228
rect 11550 15164 11614 15228
rect 11630 15164 11694 15228
rect 11710 15164 11774 15228
rect 11790 15164 11854 15228
rect 11870 15164 11934 15228
rect 11950 15164 12014 15228
rect 12030 15164 12094 15228
rect 12110 15164 12174 15228
rect 12190 15164 12254 15228
rect 12270 15164 12334 15228
rect 12350 15164 12414 15228
rect 12430 15164 12494 15228
rect 12510 15164 12574 15228
rect 12590 15164 12654 15228
rect 12670 15164 12734 15228
rect 12750 15164 12814 15228
rect 12830 15164 12894 15228
rect 12910 15164 12974 15228
rect 12990 15164 13054 15228
rect 13070 15164 13134 15228
rect 13150 15164 13214 15228
rect 13230 15164 13294 15228
rect 13310 15164 13374 15228
rect 13390 15164 13454 15228
rect 13470 15164 13534 15228
rect 13550 15164 13614 15228
rect 13630 15164 13694 15228
rect 13710 15164 13774 15228
rect 13790 15164 13854 15228
rect 13870 15164 13934 15228
rect 13950 15164 14014 15228
rect 14030 15164 14094 15228
rect 14110 15164 14174 15228
rect 14190 15164 14254 15228
rect 14270 15164 14334 15228
rect 14350 15164 14414 15228
rect 14430 15164 14494 15228
rect 14510 15164 14574 15228
rect 14590 15164 14654 15228
rect 14670 15164 14734 15228
rect 14750 15164 14814 15228
rect 14830 15164 14894 15228
rect 10190 15083 10254 15147
rect 10270 15083 10334 15147
rect 10350 15083 10414 15147
rect 10430 15083 10494 15147
rect 10510 15083 10574 15147
rect 10590 15083 10654 15147
rect 10670 15083 10734 15147
rect 10750 15083 10814 15147
rect 10830 15083 10894 15147
rect 10910 15083 10974 15147
rect 10990 15083 11054 15147
rect 11070 15083 11134 15147
rect 11150 15083 11214 15147
rect 11230 15083 11294 15147
rect 11310 15083 11374 15147
rect 11390 15083 11454 15147
rect 11470 15083 11534 15147
rect 11550 15083 11614 15147
rect 11630 15083 11694 15147
rect 11710 15083 11774 15147
rect 11790 15083 11854 15147
rect 11870 15083 11934 15147
rect 11950 15083 12014 15147
rect 12030 15083 12094 15147
rect 12110 15083 12174 15147
rect 12190 15083 12254 15147
rect 12270 15083 12334 15147
rect 12350 15083 12414 15147
rect 12430 15083 12494 15147
rect 12510 15083 12574 15147
rect 12590 15083 12654 15147
rect 12670 15083 12734 15147
rect 12750 15083 12814 15147
rect 12830 15083 12894 15147
rect 12910 15083 12974 15147
rect 12990 15083 13054 15147
rect 13070 15083 13134 15147
rect 13150 15083 13214 15147
rect 13230 15083 13294 15147
rect 13310 15083 13374 15147
rect 13390 15083 13454 15147
rect 13470 15083 13534 15147
rect 13550 15083 13614 15147
rect 13630 15083 13694 15147
rect 13710 15083 13774 15147
rect 13790 15083 13854 15147
rect 13870 15083 13934 15147
rect 13950 15083 14014 15147
rect 14030 15083 14094 15147
rect 14110 15083 14174 15147
rect 14190 15083 14254 15147
rect 14270 15083 14334 15147
rect 14350 15083 14414 15147
rect 14430 15083 14494 15147
rect 14510 15083 14574 15147
rect 14590 15083 14654 15147
rect 14670 15083 14734 15147
rect 14750 15083 14814 15147
rect 14830 15083 14894 15147
rect 10190 15002 10254 15066
rect 10270 15002 10334 15066
rect 10350 15002 10414 15066
rect 10430 15002 10494 15066
rect 10510 15002 10574 15066
rect 10590 15002 10654 15066
rect 10670 15002 10734 15066
rect 10750 15002 10814 15066
rect 10830 15002 10894 15066
rect 10910 15002 10974 15066
rect 10990 15002 11054 15066
rect 11070 15002 11134 15066
rect 11150 15002 11214 15066
rect 11230 15002 11294 15066
rect 11310 15002 11374 15066
rect 11390 15002 11454 15066
rect 11470 15002 11534 15066
rect 11550 15002 11614 15066
rect 11630 15002 11694 15066
rect 11710 15002 11774 15066
rect 11790 15002 11854 15066
rect 11870 15002 11934 15066
rect 11950 15002 12014 15066
rect 12030 15002 12094 15066
rect 12110 15002 12174 15066
rect 12190 15002 12254 15066
rect 12270 15002 12334 15066
rect 12350 15002 12414 15066
rect 12430 15002 12494 15066
rect 12510 15002 12574 15066
rect 12590 15002 12654 15066
rect 12670 15002 12734 15066
rect 12750 15002 12814 15066
rect 12830 15002 12894 15066
rect 12910 15002 12974 15066
rect 12990 15002 13054 15066
rect 13070 15002 13134 15066
rect 13150 15002 13214 15066
rect 13230 15002 13294 15066
rect 13310 15002 13374 15066
rect 13390 15002 13454 15066
rect 13470 15002 13534 15066
rect 13550 15002 13614 15066
rect 13630 15002 13694 15066
rect 13710 15002 13774 15066
rect 13790 15002 13854 15066
rect 13870 15002 13934 15066
rect 13950 15002 14014 15066
rect 14030 15002 14094 15066
rect 14110 15002 14174 15066
rect 14190 15002 14254 15066
rect 14270 15002 14334 15066
rect 14350 15002 14414 15066
rect 14430 15002 14494 15066
rect 14510 15002 14574 15066
rect 14590 15002 14654 15066
rect 14670 15002 14734 15066
rect 14750 15002 14814 15066
rect 14830 15002 14894 15066
rect 10190 14921 10254 14985
rect 10270 14921 10334 14985
rect 10350 14921 10414 14985
rect 10430 14921 10494 14985
rect 10510 14921 10574 14985
rect 10590 14921 10654 14985
rect 10670 14921 10734 14985
rect 10750 14921 10814 14985
rect 10830 14921 10894 14985
rect 10910 14921 10974 14985
rect 10990 14921 11054 14985
rect 11070 14921 11134 14985
rect 11150 14921 11214 14985
rect 11230 14921 11294 14985
rect 11310 14921 11374 14985
rect 11390 14921 11454 14985
rect 11470 14921 11534 14985
rect 11550 14921 11614 14985
rect 11630 14921 11694 14985
rect 11710 14921 11774 14985
rect 11790 14921 11854 14985
rect 11870 14921 11934 14985
rect 11950 14921 12014 14985
rect 12030 14921 12094 14985
rect 12110 14921 12174 14985
rect 12190 14921 12254 14985
rect 12270 14921 12334 14985
rect 12350 14921 12414 14985
rect 12430 14921 12494 14985
rect 12510 14921 12574 14985
rect 12590 14921 12654 14985
rect 12670 14921 12734 14985
rect 12750 14921 12814 14985
rect 12830 14921 12894 14985
rect 12910 14921 12974 14985
rect 12990 14921 13054 14985
rect 13070 14921 13134 14985
rect 13150 14921 13214 14985
rect 13230 14921 13294 14985
rect 13310 14921 13374 14985
rect 13390 14921 13454 14985
rect 13470 14921 13534 14985
rect 13550 14921 13614 14985
rect 13630 14921 13694 14985
rect 13710 14921 13774 14985
rect 13790 14921 13854 14985
rect 13870 14921 13934 14985
rect 13950 14921 14014 14985
rect 14030 14921 14094 14985
rect 14110 14921 14174 14985
rect 14190 14921 14254 14985
rect 14270 14921 14334 14985
rect 14350 14921 14414 14985
rect 14430 14921 14494 14985
rect 14510 14921 14574 14985
rect 14590 14921 14654 14985
rect 14670 14921 14734 14985
rect 14750 14921 14814 14985
rect 14830 14921 14894 14985
rect 10190 14840 10254 14904
rect 10270 14840 10334 14904
rect 10350 14840 10414 14904
rect 10430 14840 10494 14904
rect 10510 14840 10574 14904
rect 10590 14840 10654 14904
rect 10670 14840 10734 14904
rect 10750 14840 10814 14904
rect 10830 14840 10894 14904
rect 10910 14840 10974 14904
rect 10990 14840 11054 14904
rect 11070 14840 11134 14904
rect 11150 14840 11214 14904
rect 11230 14840 11294 14904
rect 11310 14840 11374 14904
rect 11390 14840 11454 14904
rect 11470 14840 11534 14904
rect 11550 14840 11614 14904
rect 11630 14840 11694 14904
rect 11710 14840 11774 14904
rect 11790 14840 11854 14904
rect 11870 14840 11934 14904
rect 11950 14840 12014 14904
rect 12030 14840 12094 14904
rect 12110 14840 12174 14904
rect 12190 14840 12254 14904
rect 12270 14840 12334 14904
rect 12350 14840 12414 14904
rect 12430 14840 12494 14904
rect 12510 14840 12574 14904
rect 12590 14840 12654 14904
rect 12670 14840 12734 14904
rect 12750 14840 12814 14904
rect 12830 14840 12894 14904
rect 12910 14840 12974 14904
rect 12990 14840 13054 14904
rect 13070 14840 13134 14904
rect 13150 14840 13214 14904
rect 13230 14840 13294 14904
rect 13310 14840 13374 14904
rect 13390 14840 13454 14904
rect 13470 14840 13534 14904
rect 13550 14840 13614 14904
rect 13630 14840 13694 14904
rect 13710 14840 13774 14904
rect 13790 14840 13854 14904
rect 13870 14840 13934 14904
rect 13950 14840 14014 14904
rect 14030 14840 14094 14904
rect 14110 14840 14174 14904
rect 14190 14840 14254 14904
rect 14270 14840 14334 14904
rect 14350 14840 14414 14904
rect 14430 14840 14494 14904
rect 14510 14840 14574 14904
rect 14590 14840 14654 14904
rect 14670 14840 14734 14904
rect 14750 14840 14814 14904
rect 14830 14840 14894 14904
rect 10190 14759 10254 14823
rect 10270 14759 10334 14823
rect 10350 14759 10414 14823
rect 10430 14759 10494 14823
rect 10510 14759 10574 14823
rect 10590 14759 10654 14823
rect 10670 14759 10734 14823
rect 10750 14759 10814 14823
rect 10830 14759 10894 14823
rect 10910 14759 10974 14823
rect 10990 14759 11054 14823
rect 11070 14759 11134 14823
rect 11150 14759 11214 14823
rect 11230 14759 11294 14823
rect 11310 14759 11374 14823
rect 11390 14759 11454 14823
rect 11470 14759 11534 14823
rect 11550 14759 11614 14823
rect 11630 14759 11694 14823
rect 11710 14759 11774 14823
rect 11790 14759 11854 14823
rect 11870 14759 11934 14823
rect 11950 14759 12014 14823
rect 12030 14759 12094 14823
rect 12110 14759 12174 14823
rect 12190 14759 12254 14823
rect 12270 14759 12334 14823
rect 12350 14759 12414 14823
rect 12430 14759 12494 14823
rect 12510 14759 12574 14823
rect 12590 14759 12654 14823
rect 12670 14759 12734 14823
rect 12750 14759 12814 14823
rect 12830 14759 12894 14823
rect 12910 14759 12974 14823
rect 12990 14759 13054 14823
rect 13070 14759 13134 14823
rect 13150 14759 13214 14823
rect 13230 14759 13294 14823
rect 13310 14759 13374 14823
rect 13390 14759 13454 14823
rect 13470 14759 13534 14823
rect 13550 14759 13614 14823
rect 13630 14759 13694 14823
rect 13710 14759 13774 14823
rect 13790 14759 13854 14823
rect 13870 14759 13934 14823
rect 13950 14759 14014 14823
rect 14030 14759 14094 14823
rect 14110 14759 14174 14823
rect 14190 14759 14254 14823
rect 14270 14759 14334 14823
rect 14350 14759 14414 14823
rect 14430 14759 14494 14823
rect 14510 14759 14574 14823
rect 14590 14759 14654 14823
rect 14670 14759 14734 14823
rect 14750 14759 14814 14823
rect 14830 14759 14894 14823
rect 10190 14678 10254 14742
rect 10270 14678 10334 14742
rect 10350 14678 10414 14742
rect 10430 14678 10494 14742
rect 10510 14678 10574 14742
rect 10590 14678 10654 14742
rect 10670 14678 10734 14742
rect 10750 14678 10814 14742
rect 10830 14678 10894 14742
rect 10910 14678 10974 14742
rect 10990 14678 11054 14742
rect 11070 14678 11134 14742
rect 11150 14678 11214 14742
rect 11230 14678 11294 14742
rect 11310 14678 11374 14742
rect 11390 14678 11454 14742
rect 11470 14678 11534 14742
rect 11550 14678 11614 14742
rect 11630 14678 11694 14742
rect 11710 14678 11774 14742
rect 11790 14678 11854 14742
rect 11870 14678 11934 14742
rect 11950 14678 12014 14742
rect 12030 14678 12094 14742
rect 12110 14678 12174 14742
rect 12190 14678 12254 14742
rect 12270 14678 12334 14742
rect 12350 14678 12414 14742
rect 12430 14678 12494 14742
rect 12510 14678 12574 14742
rect 12590 14678 12654 14742
rect 12670 14678 12734 14742
rect 12750 14678 12814 14742
rect 12830 14678 12894 14742
rect 12910 14678 12974 14742
rect 12990 14678 13054 14742
rect 13070 14678 13134 14742
rect 13150 14678 13214 14742
rect 13230 14678 13294 14742
rect 13310 14678 13374 14742
rect 13390 14678 13454 14742
rect 13470 14678 13534 14742
rect 13550 14678 13614 14742
rect 13630 14678 13694 14742
rect 13710 14678 13774 14742
rect 13790 14678 13854 14742
rect 13870 14678 13934 14742
rect 13950 14678 14014 14742
rect 14030 14678 14094 14742
rect 14110 14678 14174 14742
rect 14190 14678 14254 14742
rect 14270 14678 14334 14742
rect 14350 14678 14414 14742
rect 14430 14678 14494 14742
rect 14510 14678 14574 14742
rect 14590 14678 14654 14742
rect 14670 14678 14734 14742
rect 14750 14678 14814 14742
rect 14830 14678 14894 14742
rect 10190 14597 10254 14661
rect 10270 14597 10334 14661
rect 10350 14597 10414 14661
rect 10430 14597 10494 14661
rect 10510 14597 10574 14661
rect 10590 14597 10654 14661
rect 10670 14597 10734 14661
rect 10750 14597 10814 14661
rect 10830 14597 10894 14661
rect 10910 14597 10974 14661
rect 10990 14597 11054 14661
rect 11070 14597 11134 14661
rect 11150 14597 11214 14661
rect 11230 14597 11294 14661
rect 11310 14597 11374 14661
rect 11390 14597 11454 14661
rect 11470 14597 11534 14661
rect 11550 14597 11614 14661
rect 11630 14597 11694 14661
rect 11710 14597 11774 14661
rect 11790 14597 11854 14661
rect 11870 14597 11934 14661
rect 11950 14597 12014 14661
rect 12030 14597 12094 14661
rect 12110 14597 12174 14661
rect 12190 14597 12254 14661
rect 12270 14597 12334 14661
rect 12350 14597 12414 14661
rect 12430 14597 12494 14661
rect 12510 14597 12574 14661
rect 12590 14597 12654 14661
rect 12670 14597 12734 14661
rect 12750 14597 12814 14661
rect 12830 14597 12894 14661
rect 12910 14597 12974 14661
rect 12990 14597 13054 14661
rect 13070 14597 13134 14661
rect 13150 14597 13214 14661
rect 13230 14597 13294 14661
rect 13310 14597 13374 14661
rect 13390 14597 13454 14661
rect 13470 14597 13534 14661
rect 13550 14597 13614 14661
rect 13630 14597 13694 14661
rect 13710 14597 13774 14661
rect 13790 14597 13854 14661
rect 13870 14597 13934 14661
rect 13950 14597 14014 14661
rect 14030 14597 14094 14661
rect 14110 14597 14174 14661
rect 14190 14597 14254 14661
rect 14270 14597 14334 14661
rect 14350 14597 14414 14661
rect 14430 14597 14494 14661
rect 14510 14597 14574 14661
rect 14590 14597 14654 14661
rect 14670 14597 14734 14661
rect 14750 14597 14814 14661
rect 14830 14597 14894 14661
rect 10190 14515 10254 14579
rect 10270 14515 10334 14579
rect 10350 14515 10414 14579
rect 10430 14515 10494 14579
rect 10510 14515 10574 14579
rect 10590 14515 10654 14579
rect 10670 14515 10734 14579
rect 10750 14515 10814 14579
rect 10830 14515 10894 14579
rect 10910 14515 10974 14579
rect 10990 14515 11054 14579
rect 11070 14515 11134 14579
rect 11150 14515 11214 14579
rect 11230 14515 11294 14579
rect 11310 14515 11374 14579
rect 11390 14515 11454 14579
rect 11470 14515 11534 14579
rect 11550 14515 11614 14579
rect 11630 14515 11694 14579
rect 11710 14515 11774 14579
rect 11790 14515 11854 14579
rect 11870 14515 11934 14579
rect 11950 14515 12014 14579
rect 12030 14515 12094 14579
rect 12110 14515 12174 14579
rect 12190 14515 12254 14579
rect 12270 14515 12334 14579
rect 12350 14515 12414 14579
rect 12430 14515 12494 14579
rect 12510 14515 12574 14579
rect 12590 14515 12654 14579
rect 12670 14515 12734 14579
rect 12750 14515 12814 14579
rect 12830 14515 12894 14579
rect 12910 14515 12974 14579
rect 12990 14515 13054 14579
rect 13070 14515 13134 14579
rect 13150 14515 13214 14579
rect 13230 14515 13294 14579
rect 13310 14515 13374 14579
rect 13390 14515 13454 14579
rect 13470 14515 13534 14579
rect 13550 14515 13614 14579
rect 13630 14515 13694 14579
rect 13710 14515 13774 14579
rect 13790 14515 13854 14579
rect 13870 14515 13934 14579
rect 13950 14515 14014 14579
rect 14030 14515 14094 14579
rect 14110 14515 14174 14579
rect 14190 14515 14254 14579
rect 14270 14515 14334 14579
rect 14350 14515 14414 14579
rect 14430 14515 14494 14579
rect 14510 14515 14574 14579
rect 14590 14515 14654 14579
rect 14670 14515 14734 14579
rect 14750 14515 14814 14579
rect 14830 14515 14894 14579
rect 10190 14433 10254 14497
rect 10270 14433 10334 14497
rect 10350 14433 10414 14497
rect 10430 14433 10494 14497
rect 10510 14433 10574 14497
rect 10590 14433 10654 14497
rect 10670 14433 10734 14497
rect 10750 14433 10814 14497
rect 10830 14433 10894 14497
rect 10910 14433 10974 14497
rect 10990 14433 11054 14497
rect 11070 14433 11134 14497
rect 11150 14433 11214 14497
rect 11230 14433 11294 14497
rect 11310 14433 11374 14497
rect 11390 14433 11454 14497
rect 11470 14433 11534 14497
rect 11550 14433 11614 14497
rect 11630 14433 11694 14497
rect 11710 14433 11774 14497
rect 11790 14433 11854 14497
rect 11870 14433 11934 14497
rect 11950 14433 12014 14497
rect 12030 14433 12094 14497
rect 12110 14433 12174 14497
rect 12190 14433 12254 14497
rect 12270 14433 12334 14497
rect 12350 14433 12414 14497
rect 12430 14433 12494 14497
rect 12510 14433 12574 14497
rect 12590 14433 12654 14497
rect 12670 14433 12734 14497
rect 12750 14433 12814 14497
rect 12830 14433 12894 14497
rect 12910 14433 12974 14497
rect 12990 14433 13054 14497
rect 13070 14433 13134 14497
rect 13150 14433 13214 14497
rect 13230 14433 13294 14497
rect 13310 14433 13374 14497
rect 13390 14433 13454 14497
rect 13470 14433 13534 14497
rect 13550 14433 13614 14497
rect 13630 14433 13694 14497
rect 13710 14433 13774 14497
rect 13790 14433 13854 14497
rect 13870 14433 13934 14497
rect 13950 14433 14014 14497
rect 14030 14433 14094 14497
rect 14110 14433 14174 14497
rect 14190 14433 14254 14497
rect 14270 14433 14334 14497
rect 14350 14433 14414 14497
rect 14430 14433 14494 14497
rect 14510 14433 14574 14497
rect 14590 14433 14654 14497
rect 14670 14433 14734 14497
rect 14750 14433 14814 14497
rect 14830 14433 14894 14497
rect 10190 14351 10254 14415
rect 10270 14351 10334 14415
rect 10350 14351 10414 14415
rect 10430 14351 10494 14415
rect 10510 14351 10574 14415
rect 10590 14351 10654 14415
rect 10670 14351 10734 14415
rect 10750 14351 10814 14415
rect 10830 14351 10894 14415
rect 10910 14351 10974 14415
rect 10990 14351 11054 14415
rect 11070 14351 11134 14415
rect 11150 14351 11214 14415
rect 11230 14351 11294 14415
rect 11310 14351 11374 14415
rect 11390 14351 11454 14415
rect 11470 14351 11534 14415
rect 11550 14351 11614 14415
rect 11630 14351 11694 14415
rect 11710 14351 11774 14415
rect 11790 14351 11854 14415
rect 11870 14351 11934 14415
rect 11950 14351 12014 14415
rect 12030 14351 12094 14415
rect 12110 14351 12174 14415
rect 12190 14351 12254 14415
rect 12270 14351 12334 14415
rect 12350 14351 12414 14415
rect 12430 14351 12494 14415
rect 12510 14351 12574 14415
rect 12590 14351 12654 14415
rect 12670 14351 12734 14415
rect 12750 14351 12814 14415
rect 12830 14351 12894 14415
rect 12910 14351 12974 14415
rect 12990 14351 13054 14415
rect 13070 14351 13134 14415
rect 13150 14351 13214 14415
rect 13230 14351 13294 14415
rect 13310 14351 13374 14415
rect 13390 14351 13454 14415
rect 13470 14351 13534 14415
rect 13550 14351 13614 14415
rect 13630 14351 13694 14415
rect 13710 14351 13774 14415
rect 13790 14351 13854 14415
rect 13870 14351 13934 14415
rect 13950 14351 14014 14415
rect 14030 14351 14094 14415
rect 14110 14351 14174 14415
rect 14190 14351 14254 14415
rect 14270 14351 14334 14415
rect 14350 14351 14414 14415
rect 14430 14351 14494 14415
rect 14510 14351 14574 14415
rect 14590 14351 14654 14415
rect 14670 14351 14734 14415
rect 14750 14351 14814 14415
rect 14830 14351 14894 14415
rect 10190 14269 10254 14333
rect 10270 14269 10334 14333
rect 10350 14269 10414 14333
rect 10430 14269 10494 14333
rect 10510 14269 10574 14333
rect 10590 14269 10654 14333
rect 10670 14269 10734 14333
rect 10750 14269 10814 14333
rect 10830 14269 10894 14333
rect 10910 14269 10974 14333
rect 10990 14269 11054 14333
rect 11070 14269 11134 14333
rect 11150 14269 11214 14333
rect 11230 14269 11294 14333
rect 11310 14269 11374 14333
rect 11390 14269 11454 14333
rect 11470 14269 11534 14333
rect 11550 14269 11614 14333
rect 11630 14269 11694 14333
rect 11710 14269 11774 14333
rect 11790 14269 11854 14333
rect 11870 14269 11934 14333
rect 11950 14269 12014 14333
rect 12030 14269 12094 14333
rect 12110 14269 12174 14333
rect 12190 14269 12254 14333
rect 12270 14269 12334 14333
rect 12350 14269 12414 14333
rect 12430 14269 12494 14333
rect 12510 14269 12574 14333
rect 12590 14269 12654 14333
rect 12670 14269 12734 14333
rect 12750 14269 12814 14333
rect 12830 14269 12894 14333
rect 12910 14269 12974 14333
rect 12990 14269 13054 14333
rect 13070 14269 13134 14333
rect 13150 14269 13214 14333
rect 13230 14269 13294 14333
rect 13310 14269 13374 14333
rect 13390 14269 13454 14333
rect 13470 14269 13534 14333
rect 13550 14269 13614 14333
rect 13630 14269 13694 14333
rect 13710 14269 13774 14333
rect 13790 14269 13854 14333
rect 13870 14269 13934 14333
rect 13950 14269 14014 14333
rect 14030 14269 14094 14333
rect 14110 14269 14174 14333
rect 14190 14269 14254 14333
rect 14270 14269 14334 14333
rect 14350 14269 14414 14333
rect 14430 14269 14494 14333
rect 14510 14269 14574 14333
rect 14590 14269 14654 14333
rect 14670 14269 14734 14333
rect 14750 14269 14814 14333
rect 14830 14269 14894 14333
rect 10190 14187 10254 14251
rect 10270 14187 10334 14251
rect 10350 14187 10414 14251
rect 10430 14187 10494 14251
rect 10510 14187 10574 14251
rect 10590 14187 10654 14251
rect 10670 14187 10734 14251
rect 10750 14187 10814 14251
rect 10830 14187 10894 14251
rect 10910 14187 10974 14251
rect 10990 14187 11054 14251
rect 11070 14187 11134 14251
rect 11150 14187 11214 14251
rect 11230 14187 11294 14251
rect 11310 14187 11374 14251
rect 11390 14187 11454 14251
rect 11470 14187 11534 14251
rect 11550 14187 11614 14251
rect 11630 14187 11694 14251
rect 11710 14187 11774 14251
rect 11790 14187 11854 14251
rect 11870 14187 11934 14251
rect 11950 14187 12014 14251
rect 12030 14187 12094 14251
rect 12110 14187 12174 14251
rect 12190 14187 12254 14251
rect 12270 14187 12334 14251
rect 12350 14187 12414 14251
rect 12430 14187 12494 14251
rect 12510 14187 12574 14251
rect 12590 14187 12654 14251
rect 12670 14187 12734 14251
rect 12750 14187 12814 14251
rect 12830 14187 12894 14251
rect 12910 14187 12974 14251
rect 12990 14187 13054 14251
rect 13070 14187 13134 14251
rect 13150 14187 13214 14251
rect 13230 14187 13294 14251
rect 13310 14187 13374 14251
rect 13390 14187 13454 14251
rect 13470 14187 13534 14251
rect 13550 14187 13614 14251
rect 13630 14187 13694 14251
rect 13710 14187 13774 14251
rect 13790 14187 13854 14251
rect 13870 14187 13934 14251
rect 13950 14187 14014 14251
rect 14030 14187 14094 14251
rect 14110 14187 14174 14251
rect 14190 14187 14254 14251
rect 14270 14187 14334 14251
rect 14350 14187 14414 14251
rect 14430 14187 14494 14251
rect 14510 14187 14574 14251
rect 14590 14187 14654 14251
rect 14670 14187 14734 14251
rect 14750 14187 14814 14251
rect 14830 14187 14894 14251
rect 10190 14105 10254 14169
rect 10270 14105 10334 14169
rect 10350 14105 10414 14169
rect 10430 14105 10494 14169
rect 10510 14105 10574 14169
rect 10590 14105 10654 14169
rect 10670 14105 10734 14169
rect 10750 14105 10814 14169
rect 10830 14105 10894 14169
rect 10910 14105 10974 14169
rect 10990 14105 11054 14169
rect 11070 14105 11134 14169
rect 11150 14105 11214 14169
rect 11230 14105 11294 14169
rect 11310 14105 11374 14169
rect 11390 14105 11454 14169
rect 11470 14105 11534 14169
rect 11550 14105 11614 14169
rect 11630 14105 11694 14169
rect 11710 14105 11774 14169
rect 11790 14105 11854 14169
rect 11870 14105 11934 14169
rect 11950 14105 12014 14169
rect 12030 14105 12094 14169
rect 12110 14105 12174 14169
rect 12190 14105 12254 14169
rect 12270 14105 12334 14169
rect 12350 14105 12414 14169
rect 12430 14105 12494 14169
rect 12510 14105 12574 14169
rect 12590 14105 12654 14169
rect 12670 14105 12734 14169
rect 12750 14105 12814 14169
rect 12830 14105 12894 14169
rect 12910 14105 12974 14169
rect 12990 14105 13054 14169
rect 13070 14105 13134 14169
rect 13150 14105 13214 14169
rect 13230 14105 13294 14169
rect 13310 14105 13374 14169
rect 13390 14105 13454 14169
rect 13470 14105 13534 14169
rect 13550 14105 13614 14169
rect 13630 14105 13694 14169
rect 13710 14105 13774 14169
rect 13790 14105 13854 14169
rect 13870 14105 13934 14169
rect 13950 14105 14014 14169
rect 14030 14105 14094 14169
rect 14110 14105 14174 14169
rect 14190 14105 14254 14169
rect 14270 14105 14334 14169
rect 14350 14105 14414 14169
rect 14430 14105 14494 14169
rect 14510 14105 14574 14169
rect 14590 14105 14654 14169
rect 14670 14105 14734 14169
rect 14750 14105 14814 14169
rect 14830 14105 14894 14169
rect 10190 14023 10254 14087
rect 10270 14023 10334 14087
rect 10350 14023 10414 14087
rect 10430 14023 10494 14087
rect 10510 14023 10574 14087
rect 10590 14023 10654 14087
rect 10670 14023 10734 14087
rect 10750 14023 10814 14087
rect 10830 14023 10894 14087
rect 10910 14023 10974 14087
rect 10990 14023 11054 14087
rect 11070 14023 11134 14087
rect 11150 14023 11214 14087
rect 11230 14023 11294 14087
rect 11310 14023 11374 14087
rect 11390 14023 11454 14087
rect 11470 14023 11534 14087
rect 11550 14023 11614 14087
rect 11630 14023 11694 14087
rect 11710 14023 11774 14087
rect 11790 14023 11854 14087
rect 11870 14023 11934 14087
rect 11950 14023 12014 14087
rect 12030 14023 12094 14087
rect 12110 14023 12174 14087
rect 12190 14023 12254 14087
rect 12270 14023 12334 14087
rect 12350 14023 12414 14087
rect 12430 14023 12494 14087
rect 12510 14023 12574 14087
rect 12590 14023 12654 14087
rect 12670 14023 12734 14087
rect 12750 14023 12814 14087
rect 12830 14023 12894 14087
rect 12910 14023 12974 14087
rect 12990 14023 13054 14087
rect 13070 14023 13134 14087
rect 13150 14023 13214 14087
rect 13230 14023 13294 14087
rect 13310 14023 13374 14087
rect 13390 14023 13454 14087
rect 13470 14023 13534 14087
rect 13550 14023 13614 14087
rect 13630 14023 13694 14087
rect 13710 14023 13774 14087
rect 13790 14023 13854 14087
rect 13870 14023 13934 14087
rect 13950 14023 14014 14087
rect 14030 14023 14094 14087
rect 14110 14023 14174 14087
rect 14190 14023 14254 14087
rect 14270 14023 14334 14087
rect 14350 14023 14414 14087
rect 14430 14023 14494 14087
rect 14510 14023 14574 14087
rect 14590 14023 14654 14087
rect 14670 14023 14734 14087
rect 14750 14023 14814 14087
rect 14830 14023 14894 14087
rect 10190 13941 10254 14005
rect 10270 13941 10334 14005
rect 10350 13941 10414 14005
rect 10430 13941 10494 14005
rect 10510 13941 10574 14005
rect 10590 13941 10654 14005
rect 10670 13941 10734 14005
rect 10750 13941 10814 14005
rect 10830 13941 10894 14005
rect 10910 13941 10974 14005
rect 10990 13941 11054 14005
rect 11070 13941 11134 14005
rect 11150 13941 11214 14005
rect 11230 13941 11294 14005
rect 11310 13941 11374 14005
rect 11390 13941 11454 14005
rect 11470 13941 11534 14005
rect 11550 13941 11614 14005
rect 11630 13941 11694 14005
rect 11710 13941 11774 14005
rect 11790 13941 11854 14005
rect 11870 13941 11934 14005
rect 11950 13941 12014 14005
rect 12030 13941 12094 14005
rect 12110 13941 12174 14005
rect 12190 13941 12254 14005
rect 12270 13941 12334 14005
rect 12350 13941 12414 14005
rect 12430 13941 12494 14005
rect 12510 13941 12574 14005
rect 12590 13941 12654 14005
rect 12670 13941 12734 14005
rect 12750 13941 12814 14005
rect 12830 13941 12894 14005
rect 12910 13941 12974 14005
rect 12990 13941 13054 14005
rect 13070 13941 13134 14005
rect 13150 13941 13214 14005
rect 13230 13941 13294 14005
rect 13310 13941 13374 14005
rect 13390 13941 13454 14005
rect 13470 13941 13534 14005
rect 13550 13941 13614 14005
rect 13630 13941 13694 14005
rect 13710 13941 13774 14005
rect 13790 13941 13854 14005
rect 13870 13941 13934 14005
rect 13950 13941 14014 14005
rect 14030 13941 14094 14005
rect 14110 13941 14174 14005
rect 14190 13941 14254 14005
rect 14270 13941 14334 14005
rect 14350 13941 14414 14005
rect 14430 13941 14494 14005
rect 14510 13941 14574 14005
rect 14590 13941 14654 14005
rect 14670 13941 14734 14005
rect 14750 13941 14814 14005
rect 14830 13941 14894 14005
rect 10190 13859 10254 13923
rect 10270 13859 10334 13923
rect 10350 13859 10414 13923
rect 10430 13859 10494 13923
rect 10510 13859 10574 13923
rect 10590 13859 10654 13923
rect 10670 13859 10734 13923
rect 10750 13859 10814 13923
rect 10830 13859 10894 13923
rect 10910 13859 10974 13923
rect 10990 13859 11054 13923
rect 11070 13859 11134 13923
rect 11150 13859 11214 13923
rect 11230 13859 11294 13923
rect 11310 13859 11374 13923
rect 11390 13859 11454 13923
rect 11470 13859 11534 13923
rect 11550 13859 11614 13923
rect 11630 13859 11694 13923
rect 11710 13859 11774 13923
rect 11790 13859 11854 13923
rect 11870 13859 11934 13923
rect 11950 13859 12014 13923
rect 12030 13859 12094 13923
rect 12110 13859 12174 13923
rect 12190 13859 12254 13923
rect 12270 13859 12334 13923
rect 12350 13859 12414 13923
rect 12430 13859 12494 13923
rect 12510 13859 12574 13923
rect 12590 13859 12654 13923
rect 12670 13859 12734 13923
rect 12750 13859 12814 13923
rect 12830 13859 12894 13923
rect 12910 13859 12974 13923
rect 12990 13859 13054 13923
rect 13070 13859 13134 13923
rect 13150 13859 13214 13923
rect 13230 13859 13294 13923
rect 13310 13859 13374 13923
rect 13390 13859 13454 13923
rect 13470 13859 13534 13923
rect 13550 13859 13614 13923
rect 13630 13859 13694 13923
rect 13710 13859 13774 13923
rect 13790 13859 13854 13923
rect 13870 13859 13934 13923
rect 13950 13859 14014 13923
rect 14030 13859 14094 13923
rect 14110 13859 14174 13923
rect 14190 13859 14254 13923
rect 14270 13859 14334 13923
rect 14350 13859 14414 13923
rect 14430 13859 14494 13923
rect 14510 13859 14574 13923
rect 14590 13859 14654 13923
rect 14670 13859 14734 13923
rect 14750 13859 14814 13923
rect 14830 13859 14894 13923
rect 10190 13777 10254 13841
rect 10270 13777 10334 13841
rect 10350 13777 10414 13841
rect 10430 13777 10494 13841
rect 10510 13777 10574 13841
rect 10590 13777 10654 13841
rect 10670 13777 10734 13841
rect 10750 13777 10814 13841
rect 10830 13777 10894 13841
rect 10910 13777 10974 13841
rect 10990 13777 11054 13841
rect 11070 13777 11134 13841
rect 11150 13777 11214 13841
rect 11230 13777 11294 13841
rect 11310 13777 11374 13841
rect 11390 13777 11454 13841
rect 11470 13777 11534 13841
rect 11550 13777 11614 13841
rect 11630 13777 11694 13841
rect 11710 13777 11774 13841
rect 11790 13777 11854 13841
rect 11870 13777 11934 13841
rect 11950 13777 12014 13841
rect 12030 13777 12094 13841
rect 12110 13777 12174 13841
rect 12190 13777 12254 13841
rect 12270 13777 12334 13841
rect 12350 13777 12414 13841
rect 12430 13777 12494 13841
rect 12510 13777 12574 13841
rect 12590 13777 12654 13841
rect 12670 13777 12734 13841
rect 12750 13777 12814 13841
rect 12830 13777 12894 13841
rect 12910 13777 12974 13841
rect 12990 13777 13054 13841
rect 13070 13777 13134 13841
rect 13150 13777 13214 13841
rect 13230 13777 13294 13841
rect 13310 13777 13374 13841
rect 13390 13777 13454 13841
rect 13470 13777 13534 13841
rect 13550 13777 13614 13841
rect 13630 13777 13694 13841
rect 13710 13777 13774 13841
rect 13790 13777 13854 13841
rect 13870 13777 13934 13841
rect 13950 13777 14014 13841
rect 14030 13777 14094 13841
rect 14110 13777 14174 13841
rect 14190 13777 14254 13841
rect 14270 13777 14334 13841
rect 14350 13777 14414 13841
rect 14430 13777 14494 13841
rect 14510 13777 14574 13841
rect 14590 13777 14654 13841
rect 14670 13777 14734 13841
rect 14750 13777 14814 13841
rect 14830 13777 14894 13841
rect 10190 13695 10254 13759
rect 10270 13695 10334 13759
rect 10350 13695 10414 13759
rect 10430 13695 10494 13759
rect 10510 13695 10574 13759
rect 10590 13695 10654 13759
rect 10670 13695 10734 13759
rect 10750 13695 10814 13759
rect 10830 13695 10894 13759
rect 10910 13695 10974 13759
rect 10990 13695 11054 13759
rect 11070 13695 11134 13759
rect 11150 13695 11214 13759
rect 11230 13695 11294 13759
rect 11310 13695 11374 13759
rect 11390 13695 11454 13759
rect 11470 13695 11534 13759
rect 11550 13695 11614 13759
rect 11630 13695 11694 13759
rect 11710 13695 11774 13759
rect 11790 13695 11854 13759
rect 11870 13695 11934 13759
rect 11950 13695 12014 13759
rect 12030 13695 12094 13759
rect 12110 13695 12174 13759
rect 12190 13695 12254 13759
rect 12270 13695 12334 13759
rect 12350 13695 12414 13759
rect 12430 13695 12494 13759
rect 12510 13695 12574 13759
rect 12590 13695 12654 13759
rect 12670 13695 12734 13759
rect 12750 13695 12814 13759
rect 12830 13695 12894 13759
rect 12910 13695 12974 13759
rect 12990 13695 13054 13759
rect 13070 13695 13134 13759
rect 13150 13695 13214 13759
rect 13230 13695 13294 13759
rect 13310 13695 13374 13759
rect 13390 13695 13454 13759
rect 13470 13695 13534 13759
rect 13550 13695 13614 13759
rect 13630 13695 13694 13759
rect 13710 13695 13774 13759
rect 13790 13695 13854 13759
rect 13870 13695 13934 13759
rect 13950 13695 14014 13759
rect 14030 13695 14094 13759
rect 14110 13695 14174 13759
rect 14190 13695 14254 13759
rect 14270 13695 14334 13759
rect 14350 13695 14414 13759
rect 14430 13695 14494 13759
rect 14510 13695 14574 13759
rect 14590 13695 14654 13759
rect 14670 13695 14734 13759
rect 14750 13695 14814 13759
rect 14830 13695 14894 13759
rect 10190 13613 10254 13677
rect 10270 13613 10334 13677
rect 10350 13613 10414 13677
rect 10430 13613 10494 13677
rect 10510 13613 10574 13677
rect 10590 13613 10654 13677
rect 10670 13613 10734 13677
rect 10750 13613 10814 13677
rect 10830 13613 10894 13677
rect 10910 13613 10974 13677
rect 10990 13613 11054 13677
rect 11070 13613 11134 13677
rect 11150 13613 11214 13677
rect 11230 13613 11294 13677
rect 11310 13613 11374 13677
rect 11390 13613 11454 13677
rect 11470 13613 11534 13677
rect 11550 13613 11614 13677
rect 11630 13613 11694 13677
rect 11710 13613 11774 13677
rect 11790 13613 11854 13677
rect 11870 13613 11934 13677
rect 11950 13613 12014 13677
rect 12030 13613 12094 13677
rect 12110 13613 12174 13677
rect 12190 13613 12254 13677
rect 12270 13613 12334 13677
rect 12350 13613 12414 13677
rect 12430 13613 12494 13677
rect 12510 13613 12574 13677
rect 12590 13613 12654 13677
rect 12670 13613 12734 13677
rect 12750 13613 12814 13677
rect 12830 13613 12894 13677
rect 12910 13613 12974 13677
rect 12990 13613 13054 13677
rect 13070 13613 13134 13677
rect 13150 13613 13214 13677
rect 13230 13613 13294 13677
rect 13310 13613 13374 13677
rect 13390 13613 13454 13677
rect 13470 13613 13534 13677
rect 13550 13613 13614 13677
rect 13630 13613 13694 13677
rect 13710 13613 13774 13677
rect 13790 13613 13854 13677
rect 13870 13613 13934 13677
rect 13950 13613 14014 13677
rect 14030 13613 14094 13677
rect 14110 13613 14174 13677
rect 14190 13613 14254 13677
rect 14270 13613 14334 13677
rect 14350 13613 14414 13677
rect 14430 13613 14494 13677
rect 14510 13613 14574 13677
rect 14590 13613 14654 13677
rect 14670 13613 14734 13677
rect 14750 13613 14814 13677
rect 14830 13613 14894 13677
rect 126 13240 190 13304
rect 207 13240 271 13304
rect 288 13240 352 13304
rect 369 13240 433 13304
rect 450 13240 514 13304
rect 531 13240 595 13304
rect 612 13240 676 13304
rect 693 13240 757 13304
rect 774 13240 838 13304
rect 855 13240 919 13304
rect 936 13240 1000 13304
rect 1017 13240 1081 13304
rect 1098 13240 1162 13304
rect 1179 13240 1243 13304
rect 1260 13240 1324 13304
rect 1341 13240 1405 13304
rect 1422 13240 1486 13304
rect 1503 13240 1567 13304
rect 1584 13240 1648 13304
rect 1665 13240 1729 13304
rect 1746 13240 1810 13304
rect 1827 13240 1891 13304
rect 1908 13240 1972 13304
rect 1989 13240 2053 13304
rect 2070 13240 2134 13304
rect 2151 13240 2215 13304
rect 2232 13240 2296 13304
rect 2313 13240 2377 13304
rect 2394 13240 2458 13304
rect 2475 13240 2539 13304
rect 2556 13240 2620 13304
rect 2637 13240 2701 13304
rect 2718 13240 2782 13304
rect 2799 13240 2863 13304
rect 2880 13240 2944 13304
rect 2961 13240 3025 13304
rect 3042 13240 3106 13304
rect 3123 13240 3187 13304
rect 3204 13240 3268 13304
rect 3285 13240 3349 13304
rect 3366 13240 3430 13304
rect 3447 13240 3511 13304
rect 3528 13240 3592 13304
rect 3609 13240 3673 13304
rect 3690 13240 3754 13304
rect 3771 13240 3835 13304
rect 3852 13240 3916 13304
rect 3933 13240 3997 13304
rect 4014 13240 4078 13304
rect 4095 13240 4159 13304
rect 4176 13240 4240 13304
rect 4257 13240 4321 13304
rect 4338 13240 4402 13304
rect 4420 13240 4484 13304
rect 4502 13240 4566 13304
rect 4584 13240 4648 13304
rect 4666 13240 4730 13304
rect 4748 13240 4812 13304
rect 4830 13240 4894 13304
rect 126 13158 190 13222
rect 207 13158 271 13222
rect 288 13158 352 13222
rect 369 13158 433 13222
rect 450 13158 514 13222
rect 531 13158 595 13222
rect 612 13158 676 13222
rect 693 13158 757 13222
rect 774 13158 838 13222
rect 855 13158 919 13222
rect 936 13158 1000 13222
rect 1017 13158 1081 13222
rect 1098 13158 1162 13222
rect 1179 13158 1243 13222
rect 1260 13158 1324 13222
rect 1341 13158 1405 13222
rect 1422 13158 1486 13222
rect 1503 13158 1567 13222
rect 1584 13158 1648 13222
rect 1665 13158 1729 13222
rect 1746 13158 1810 13222
rect 1827 13158 1891 13222
rect 1908 13158 1972 13222
rect 1989 13158 2053 13222
rect 2070 13158 2134 13222
rect 2151 13158 2215 13222
rect 2232 13158 2296 13222
rect 2313 13158 2377 13222
rect 2394 13158 2458 13222
rect 2475 13158 2539 13222
rect 2556 13158 2620 13222
rect 2637 13158 2701 13222
rect 2718 13158 2782 13222
rect 2799 13158 2863 13222
rect 2880 13158 2944 13222
rect 2961 13158 3025 13222
rect 3042 13158 3106 13222
rect 3123 13158 3187 13222
rect 3204 13158 3268 13222
rect 3285 13158 3349 13222
rect 3366 13158 3430 13222
rect 3447 13158 3511 13222
rect 3528 13158 3592 13222
rect 3609 13158 3673 13222
rect 3690 13158 3754 13222
rect 3771 13158 3835 13222
rect 3852 13158 3916 13222
rect 3933 13158 3997 13222
rect 4014 13158 4078 13222
rect 4095 13158 4159 13222
rect 4176 13158 4240 13222
rect 4257 13158 4321 13222
rect 4338 13158 4402 13222
rect 4420 13158 4484 13222
rect 4502 13158 4566 13222
rect 4584 13158 4648 13222
rect 4666 13158 4730 13222
rect 4748 13158 4812 13222
rect 4830 13158 4894 13222
rect 126 13076 190 13140
rect 207 13076 271 13140
rect 288 13076 352 13140
rect 369 13076 433 13140
rect 450 13076 514 13140
rect 531 13076 595 13140
rect 612 13076 676 13140
rect 693 13076 757 13140
rect 774 13076 838 13140
rect 855 13076 919 13140
rect 936 13076 1000 13140
rect 1017 13076 1081 13140
rect 1098 13076 1162 13140
rect 1179 13076 1243 13140
rect 1260 13076 1324 13140
rect 1341 13076 1405 13140
rect 1422 13076 1486 13140
rect 1503 13076 1567 13140
rect 1584 13076 1648 13140
rect 1665 13076 1729 13140
rect 1746 13076 1810 13140
rect 1827 13076 1891 13140
rect 1908 13076 1972 13140
rect 1989 13076 2053 13140
rect 2070 13076 2134 13140
rect 2151 13076 2215 13140
rect 2232 13076 2296 13140
rect 2313 13076 2377 13140
rect 2394 13076 2458 13140
rect 2475 13076 2539 13140
rect 2556 13076 2620 13140
rect 2637 13076 2701 13140
rect 2718 13076 2782 13140
rect 2799 13076 2863 13140
rect 2880 13076 2944 13140
rect 2961 13076 3025 13140
rect 3042 13076 3106 13140
rect 3123 13076 3187 13140
rect 3204 13076 3268 13140
rect 3285 13076 3349 13140
rect 3366 13076 3430 13140
rect 3447 13076 3511 13140
rect 3528 13076 3592 13140
rect 3609 13076 3673 13140
rect 3690 13076 3754 13140
rect 3771 13076 3835 13140
rect 3852 13076 3916 13140
rect 3933 13076 3997 13140
rect 4014 13076 4078 13140
rect 4095 13076 4159 13140
rect 4176 13076 4240 13140
rect 4257 13076 4321 13140
rect 4338 13076 4402 13140
rect 4420 13076 4484 13140
rect 4502 13076 4566 13140
rect 4584 13076 4648 13140
rect 4666 13076 4730 13140
rect 4748 13076 4812 13140
rect 4830 13076 4894 13140
rect 126 12994 190 13058
rect 207 12994 271 13058
rect 288 12994 352 13058
rect 369 12994 433 13058
rect 450 12994 514 13058
rect 531 12994 595 13058
rect 612 12994 676 13058
rect 693 12994 757 13058
rect 774 12994 838 13058
rect 855 12994 919 13058
rect 936 12994 1000 13058
rect 1017 12994 1081 13058
rect 1098 12994 1162 13058
rect 1179 12994 1243 13058
rect 1260 12994 1324 13058
rect 1341 12994 1405 13058
rect 1422 12994 1486 13058
rect 1503 12994 1567 13058
rect 1584 12994 1648 13058
rect 1665 12994 1729 13058
rect 1746 12994 1810 13058
rect 1827 12994 1891 13058
rect 1908 12994 1972 13058
rect 1989 12994 2053 13058
rect 2070 12994 2134 13058
rect 2151 12994 2215 13058
rect 2232 12994 2296 13058
rect 2313 12994 2377 13058
rect 2394 12994 2458 13058
rect 2475 12994 2539 13058
rect 2556 12994 2620 13058
rect 2637 12994 2701 13058
rect 2718 12994 2782 13058
rect 2799 12994 2863 13058
rect 2880 12994 2944 13058
rect 2961 12994 3025 13058
rect 3042 12994 3106 13058
rect 3123 12994 3187 13058
rect 3204 12994 3268 13058
rect 3285 12994 3349 13058
rect 3366 12994 3430 13058
rect 3447 12994 3511 13058
rect 3528 12994 3592 13058
rect 3609 12994 3673 13058
rect 3690 12994 3754 13058
rect 3771 12994 3835 13058
rect 3852 12994 3916 13058
rect 3933 12994 3997 13058
rect 4014 12994 4078 13058
rect 4095 12994 4159 13058
rect 4176 12994 4240 13058
rect 4257 12994 4321 13058
rect 4338 12994 4402 13058
rect 4420 12994 4484 13058
rect 4502 12994 4566 13058
rect 4584 12994 4648 13058
rect 4666 12994 4730 13058
rect 4748 12994 4812 13058
rect 4830 12994 4894 13058
rect 126 12912 190 12976
rect 207 12912 271 12976
rect 288 12912 352 12976
rect 369 12912 433 12976
rect 450 12912 514 12976
rect 531 12912 595 12976
rect 612 12912 676 12976
rect 693 12912 757 12976
rect 774 12912 838 12976
rect 855 12912 919 12976
rect 936 12912 1000 12976
rect 1017 12912 1081 12976
rect 1098 12912 1162 12976
rect 1179 12912 1243 12976
rect 1260 12912 1324 12976
rect 1341 12912 1405 12976
rect 1422 12912 1486 12976
rect 1503 12912 1567 12976
rect 1584 12912 1648 12976
rect 1665 12912 1729 12976
rect 1746 12912 1810 12976
rect 1827 12912 1891 12976
rect 1908 12912 1972 12976
rect 1989 12912 2053 12976
rect 2070 12912 2134 12976
rect 2151 12912 2215 12976
rect 2232 12912 2296 12976
rect 2313 12912 2377 12976
rect 2394 12912 2458 12976
rect 2475 12912 2539 12976
rect 2556 12912 2620 12976
rect 2637 12912 2701 12976
rect 2718 12912 2782 12976
rect 2799 12912 2863 12976
rect 2880 12912 2944 12976
rect 2961 12912 3025 12976
rect 3042 12912 3106 12976
rect 3123 12912 3187 12976
rect 3204 12912 3268 12976
rect 3285 12912 3349 12976
rect 3366 12912 3430 12976
rect 3447 12912 3511 12976
rect 3528 12912 3592 12976
rect 3609 12912 3673 12976
rect 3690 12912 3754 12976
rect 3771 12912 3835 12976
rect 3852 12912 3916 12976
rect 3933 12912 3997 12976
rect 4014 12912 4078 12976
rect 4095 12912 4159 12976
rect 4176 12912 4240 12976
rect 4257 12912 4321 12976
rect 4338 12912 4402 12976
rect 4420 12912 4484 12976
rect 4502 12912 4566 12976
rect 4584 12912 4648 12976
rect 4666 12912 4730 12976
rect 4748 12912 4812 12976
rect 4830 12912 4894 12976
rect 126 12830 190 12894
rect 207 12830 271 12894
rect 288 12830 352 12894
rect 369 12830 433 12894
rect 450 12830 514 12894
rect 531 12830 595 12894
rect 612 12830 676 12894
rect 693 12830 757 12894
rect 774 12830 838 12894
rect 855 12830 919 12894
rect 936 12830 1000 12894
rect 1017 12830 1081 12894
rect 1098 12830 1162 12894
rect 1179 12830 1243 12894
rect 1260 12830 1324 12894
rect 1341 12830 1405 12894
rect 1422 12830 1486 12894
rect 1503 12830 1567 12894
rect 1584 12830 1648 12894
rect 1665 12830 1729 12894
rect 1746 12830 1810 12894
rect 1827 12830 1891 12894
rect 1908 12830 1972 12894
rect 1989 12830 2053 12894
rect 2070 12830 2134 12894
rect 2151 12830 2215 12894
rect 2232 12830 2296 12894
rect 2313 12830 2377 12894
rect 2394 12830 2458 12894
rect 2475 12830 2539 12894
rect 2556 12830 2620 12894
rect 2637 12830 2701 12894
rect 2718 12830 2782 12894
rect 2799 12830 2863 12894
rect 2880 12830 2944 12894
rect 2961 12830 3025 12894
rect 3042 12830 3106 12894
rect 3123 12830 3187 12894
rect 3204 12830 3268 12894
rect 3285 12830 3349 12894
rect 3366 12830 3430 12894
rect 3447 12830 3511 12894
rect 3528 12830 3592 12894
rect 3609 12830 3673 12894
rect 3690 12830 3754 12894
rect 3771 12830 3835 12894
rect 3852 12830 3916 12894
rect 3933 12830 3997 12894
rect 4014 12830 4078 12894
rect 4095 12830 4159 12894
rect 4176 12830 4240 12894
rect 4257 12830 4321 12894
rect 4338 12830 4402 12894
rect 4420 12830 4484 12894
rect 4502 12830 4566 12894
rect 4584 12830 4648 12894
rect 4666 12830 4730 12894
rect 4748 12830 4812 12894
rect 4830 12830 4894 12894
rect 126 12748 190 12812
rect 207 12748 271 12812
rect 288 12748 352 12812
rect 369 12748 433 12812
rect 450 12748 514 12812
rect 531 12748 595 12812
rect 612 12748 676 12812
rect 693 12748 757 12812
rect 774 12748 838 12812
rect 855 12748 919 12812
rect 936 12748 1000 12812
rect 1017 12748 1081 12812
rect 1098 12748 1162 12812
rect 1179 12748 1243 12812
rect 1260 12748 1324 12812
rect 1341 12748 1405 12812
rect 1422 12748 1486 12812
rect 1503 12748 1567 12812
rect 1584 12748 1648 12812
rect 1665 12748 1729 12812
rect 1746 12748 1810 12812
rect 1827 12748 1891 12812
rect 1908 12748 1972 12812
rect 1989 12748 2053 12812
rect 2070 12748 2134 12812
rect 2151 12748 2215 12812
rect 2232 12748 2296 12812
rect 2313 12748 2377 12812
rect 2394 12748 2458 12812
rect 2475 12748 2539 12812
rect 2556 12748 2620 12812
rect 2637 12748 2701 12812
rect 2718 12748 2782 12812
rect 2799 12748 2863 12812
rect 2880 12748 2944 12812
rect 2961 12748 3025 12812
rect 3042 12748 3106 12812
rect 3123 12748 3187 12812
rect 3204 12748 3268 12812
rect 3285 12748 3349 12812
rect 3366 12748 3430 12812
rect 3447 12748 3511 12812
rect 3528 12748 3592 12812
rect 3609 12748 3673 12812
rect 3690 12748 3754 12812
rect 3771 12748 3835 12812
rect 3852 12748 3916 12812
rect 3933 12748 3997 12812
rect 4014 12748 4078 12812
rect 4095 12748 4159 12812
rect 4176 12748 4240 12812
rect 4257 12748 4321 12812
rect 4338 12748 4402 12812
rect 4420 12748 4484 12812
rect 4502 12748 4566 12812
rect 4584 12748 4648 12812
rect 4666 12748 4730 12812
rect 4748 12748 4812 12812
rect 4830 12748 4894 12812
rect 126 12666 190 12730
rect 207 12666 271 12730
rect 288 12666 352 12730
rect 369 12666 433 12730
rect 450 12666 514 12730
rect 531 12666 595 12730
rect 612 12666 676 12730
rect 693 12666 757 12730
rect 774 12666 838 12730
rect 855 12666 919 12730
rect 936 12666 1000 12730
rect 1017 12666 1081 12730
rect 1098 12666 1162 12730
rect 1179 12666 1243 12730
rect 1260 12666 1324 12730
rect 1341 12666 1405 12730
rect 1422 12666 1486 12730
rect 1503 12666 1567 12730
rect 1584 12666 1648 12730
rect 1665 12666 1729 12730
rect 1746 12666 1810 12730
rect 1827 12666 1891 12730
rect 1908 12666 1972 12730
rect 1989 12666 2053 12730
rect 2070 12666 2134 12730
rect 2151 12666 2215 12730
rect 2232 12666 2296 12730
rect 2313 12666 2377 12730
rect 2394 12666 2458 12730
rect 2475 12666 2539 12730
rect 2556 12666 2620 12730
rect 2637 12666 2701 12730
rect 2718 12666 2782 12730
rect 2799 12666 2863 12730
rect 2880 12666 2944 12730
rect 2961 12666 3025 12730
rect 3042 12666 3106 12730
rect 3123 12666 3187 12730
rect 3204 12666 3268 12730
rect 3285 12666 3349 12730
rect 3366 12666 3430 12730
rect 3447 12666 3511 12730
rect 3528 12666 3592 12730
rect 3609 12666 3673 12730
rect 3690 12666 3754 12730
rect 3771 12666 3835 12730
rect 3852 12666 3916 12730
rect 3933 12666 3997 12730
rect 4014 12666 4078 12730
rect 4095 12666 4159 12730
rect 4176 12666 4240 12730
rect 4257 12666 4321 12730
rect 4338 12666 4402 12730
rect 4420 12666 4484 12730
rect 4502 12666 4566 12730
rect 4584 12666 4648 12730
rect 4666 12666 4730 12730
rect 4748 12666 4812 12730
rect 4830 12666 4894 12730
rect 126 12584 190 12648
rect 207 12584 271 12648
rect 288 12584 352 12648
rect 369 12584 433 12648
rect 450 12584 514 12648
rect 531 12584 595 12648
rect 612 12584 676 12648
rect 693 12584 757 12648
rect 774 12584 838 12648
rect 855 12584 919 12648
rect 936 12584 1000 12648
rect 1017 12584 1081 12648
rect 1098 12584 1162 12648
rect 1179 12584 1243 12648
rect 1260 12584 1324 12648
rect 1341 12584 1405 12648
rect 1422 12584 1486 12648
rect 1503 12584 1567 12648
rect 1584 12584 1648 12648
rect 1665 12584 1729 12648
rect 1746 12584 1810 12648
rect 1827 12584 1891 12648
rect 1908 12584 1972 12648
rect 1989 12584 2053 12648
rect 2070 12584 2134 12648
rect 2151 12584 2215 12648
rect 2232 12584 2296 12648
rect 2313 12584 2377 12648
rect 2394 12584 2458 12648
rect 2475 12584 2539 12648
rect 2556 12584 2620 12648
rect 2637 12584 2701 12648
rect 2718 12584 2782 12648
rect 2799 12584 2863 12648
rect 2880 12584 2944 12648
rect 2961 12584 3025 12648
rect 3042 12584 3106 12648
rect 3123 12584 3187 12648
rect 3204 12584 3268 12648
rect 3285 12584 3349 12648
rect 3366 12584 3430 12648
rect 3447 12584 3511 12648
rect 3528 12584 3592 12648
rect 3609 12584 3673 12648
rect 3690 12584 3754 12648
rect 3771 12584 3835 12648
rect 3852 12584 3916 12648
rect 3933 12584 3997 12648
rect 4014 12584 4078 12648
rect 4095 12584 4159 12648
rect 4176 12584 4240 12648
rect 4257 12584 4321 12648
rect 4338 12584 4402 12648
rect 4420 12584 4484 12648
rect 4502 12584 4566 12648
rect 4584 12584 4648 12648
rect 4666 12584 4730 12648
rect 4748 12584 4812 12648
rect 4830 12584 4894 12648
rect 126 12502 190 12566
rect 207 12502 271 12566
rect 288 12502 352 12566
rect 369 12502 433 12566
rect 450 12502 514 12566
rect 531 12502 595 12566
rect 612 12502 676 12566
rect 693 12502 757 12566
rect 774 12502 838 12566
rect 855 12502 919 12566
rect 936 12502 1000 12566
rect 1017 12502 1081 12566
rect 1098 12502 1162 12566
rect 1179 12502 1243 12566
rect 1260 12502 1324 12566
rect 1341 12502 1405 12566
rect 1422 12502 1486 12566
rect 1503 12502 1567 12566
rect 1584 12502 1648 12566
rect 1665 12502 1729 12566
rect 1746 12502 1810 12566
rect 1827 12502 1891 12566
rect 1908 12502 1972 12566
rect 1989 12502 2053 12566
rect 2070 12502 2134 12566
rect 2151 12502 2215 12566
rect 2232 12502 2296 12566
rect 2313 12502 2377 12566
rect 2394 12502 2458 12566
rect 2475 12502 2539 12566
rect 2556 12502 2620 12566
rect 2637 12502 2701 12566
rect 2718 12502 2782 12566
rect 2799 12502 2863 12566
rect 2880 12502 2944 12566
rect 2961 12502 3025 12566
rect 3042 12502 3106 12566
rect 3123 12502 3187 12566
rect 3204 12502 3268 12566
rect 3285 12502 3349 12566
rect 3366 12502 3430 12566
rect 3447 12502 3511 12566
rect 3528 12502 3592 12566
rect 3609 12502 3673 12566
rect 3690 12502 3754 12566
rect 3771 12502 3835 12566
rect 3852 12502 3916 12566
rect 3933 12502 3997 12566
rect 4014 12502 4078 12566
rect 4095 12502 4159 12566
rect 4176 12502 4240 12566
rect 4257 12502 4321 12566
rect 4338 12502 4402 12566
rect 4420 12502 4484 12566
rect 4502 12502 4566 12566
rect 4584 12502 4648 12566
rect 4666 12502 4730 12566
rect 4748 12502 4812 12566
rect 4830 12502 4894 12566
rect 126 12420 190 12484
rect 207 12420 271 12484
rect 288 12420 352 12484
rect 369 12420 433 12484
rect 450 12420 514 12484
rect 531 12420 595 12484
rect 612 12420 676 12484
rect 693 12420 757 12484
rect 774 12420 838 12484
rect 855 12420 919 12484
rect 936 12420 1000 12484
rect 1017 12420 1081 12484
rect 1098 12420 1162 12484
rect 1179 12420 1243 12484
rect 1260 12420 1324 12484
rect 1341 12420 1405 12484
rect 1422 12420 1486 12484
rect 1503 12420 1567 12484
rect 1584 12420 1648 12484
rect 1665 12420 1729 12484
rect 1746 12420 1810 12484
rect 1827 12420 1891 12484
rect 1908 12420 1972 12484
rect 1989 12420 2053 12484
rect 2070 12420 2134 12484
rect 2151 12420 2215 12484
rect 2232 12420 2296 12484
rect 2313 12420 2377 12484
rect 2394 12420 2458 12484
rect 2475 12420 2539 12484
rect 2556 12420 2620 12484
rect 2637 12420 2701 12484
rect 2718 12420 2782 12484
rect 2799 12420 2863 12484
rect 2880 12420 2944 12484
rect 2961 12420 3025 12484
rect 3042 12420 3106 12484
rect 3123 12420 3187 12484
rect 3204 12420 3268 12484
rect 3285 12420 3349 12484
rect 3366 12420 3430 12484
rect 3447 12420 3511 12484
rect 3528 12420 3592 12484
rect 3609 12420 3673 12484
rect 3690 12420 3754 12484
rect 3771 12420 3835 12484
rect 3852 12420 3916 12484
rect 3933 12420 3997 12484
rect 4014 12420 4078 12484
rect 4095 12420 4159 12484
rect 4176 12420 4240 12484
rect 4257 12420 4321 12484
rect 4338 12420 4402 12484
rect 4420 12420 4484 12484
rect 4502 12420 4566 12484
rect 4584 12420 4648 12484
rect 4666 12420 4730 12484
rect 4748 12420 4812 12484
rect 4830 12420 4894 12484
rect 10157 13240 10221 13304
rect 10238 13240 10302 13304
rect 10319 13240 10383 13304
rect 10400 13240 10464 13304
rect 10481 13240 10545 13304
rect 10562 13240 10626 13304
rect 10643 13240 10707 13304
rect 10724 13240 10788 13304
rect 10805 13240 10869 13304
rect 10886 13240 10950 13304
rect 10967 13240 11031 13304
rect 11048 13240 11112 13304
rect 11129 13240 11193 13304
rect 11210 13240 11274 13304
rect 11291 13240 11355 13304
rect 11372 13240 11436 13304
rect 11453 13240 11517 13304
rect 11534 13240 11598 13304
rect 11615 13240 11679 13304
rect 11696 13240 11760 13304
rect 11777 13240 11841 13304
rect 11858 13240 11922 13304
rect 11939 13240 12003 13304
rect 12020 13240 12084 13304
rect 12101 13240 12165 13304
rect 12182 13240 12246 13304
rect 12263 13240 12327 13304
rect 12344 13240 12408 13304
rect 12425 13240 12489 13304
rect 12506 13240 12570 13304
rect 12587 13240 12651 13304
rect 12668 13240 12732 13304
rect 12749 13240 12813 13304
rect 12830 13240 12894 13304
rect 12911 13240 12975 13304
rect 12992 13240 13056 13304
rect 13073 13240 13137 13304
rect 13154 13240 13218 13304
rect 13235 13240 13299 13304
rect 13316 13240 13380 13304
rect 13397 13240 13461 13304
rect 13478 13240 13542 13304
rect 13559 13240 13623 13304
rect 13640 13240 13704 13304
rect 13721 13240 13785 13304
rect 13802 13240 13866 13304
rect 13883 13240 13947 13304
rect 13964 13240 14028 13304
rect 14045 13240 14109 13304
rect 14126 13240 14190 13304
rect 14207 13240 14271 13304
rect 14288 13240 14352 13304
rect 14369 13240 14433 13304
rect 14451 13240 14515 13304
rect 14533 13240 14597 13304
rect 14615 13240 14679 13304
rect 14697 13240 14761 13304
rect 14779 13240 14843 13304
rect 14861 13240 14925 13304
rect 10157 13158 10221 13222
rect 10238 13158 10302 13222
rect 10319 13158 10383 13222
rect 10400 13158 10464 13222
rect 10481 13158 10545 13222
rect 10562 13158 10626 13222
rect 10643 13158 10707 13222
rect 10724 13158 10788 13222
rect 10805 13158 10869 13222
rect 10886 13158 10950 13222
rect 10967 13158 11031 13222
rect 11048 13158 11112 13222
rect 11129 13158 11193 13222
rect 11210 13158 11274 13222
rect 11291 13158 11355 13222
rect 11372 13158 11436 13222
rect 11453 13158 11517 13222
rect 11534 13158 11598 13222
rect 11615 13158 11679 13222
rect 11696 13158 11760 13222
rect 11777 13158 11841 13222
rect 11858 13158 11922 13222
rect 11939 13158 12003 13222
rect 12020 13158 12084 13222
rect 12101 13158 12165 13222
rect 12182 13158 12246 13222
rect 12263 13158 12327 13222
rect 12344 13158 12408 13222
rect 12425 13158 12489 13222
rect 12506 13158 12570 13222
rect 12587 13158 12651 13222
rect 12668 13158 12732 13222
rect 12749 13158 12813 13222
rect 12830 13158 12894 13222
rect 12911 13158 12975 13222
rect 12992 13158 13056 13222
rect 13073 13158 13137 13222
rect 13154 13158 13218 13222
rect 13235 13158 13299 13222
rect 13316 13158 13380 13222
rect 13397 13158 13461 13222
rect 13478 13158 13542 13222
rect 13559 13158 13623 13222
rect 13640 13158 13704 13222
rect 13721 13158 13785 13222
rect 13802 13158 13866 13222
rect 13883 13158 13947 13222
rect 13964 13158 14028 13222
rect 14045 13158 14109 13222
rect 14126 13158 14190 13222
rect 14207 13158 14271 13222
rect 14288 13158 14352 13222
rect 14369 13158 14433 13222
rect 14451 13158 14515 13222
rect 14533 13158 14597 13222
rect 14615 13158 14679 13222
rect 14697 13158 14761 13222
rect 14779 13158 14843 13222
rect 14861 13158 14925 13222
rect 10157 13076 10221 13140
rect 10238 13076 10302 13140
rect 10319 13076 10383 13140
rect 10400 13076 10464 13140
rect 10481 13076 10545 13140
rect 10562 13076 10626 13140
rect 10643 13076 10707 13140
rect 10724 13076 10788 13140
rect 10805 13076 10869 13140
rect 10886 13076 10950 13140
rect 10967 13076 11031 13140
rect 11048 13076 11112 13140
rect 11129 13076 11193 13140
rect 11210 13076 11274 13140
rect 11291 13076 11355 13140
rect 11372 13076 11436 13140
rect 11453 13076 11517 13140
rect 11534 13076 11598 13140
rect 11615 13076 11679 13140
rect 11696 13076 11760 13140
rect 11777 13076 11841 13140
rect 11858 13076 11922 13140
rect 11939 13076 12003 13140
rect 12020 13076 12084 13140
rect 12101 13076 12165 13140
rect 12182 13076 12246 13140
rect 12263 13076 12327 13140
rect 12344 13076 12408 13140
rect 12425 13076 12489 13140
rect 12506 13076 12570 13140
rect 12587 13076 12651 13140
rect 12668 13076 12732 13140
rect 12749 13076 12813 13140
rect 12830 13076 12894 13140
rect 12911 13076 12975 13140
rect 12992 13076 13056 13140
rect 13073 13076 13137 13140
rect 13154 13076 13218 13140
rect 13235 13076 13299 13140
rect 13316 13076 13380 13140
rect 13397 13076 13461 13140
rect 13478 13076 13542 13140
rect 13559 13076 13623 13140
rect 13640 13076 13704 13140
rect 13721 13076 13785 13140
rect 13802 13076 13866 13140
rect 13883 13076 13947 13140
rect 13964 13076 14028 13140
rect 14045 13076 14109 13140
rect 14126 13076 14190 13140
rect 14207 13076 14271 13140
rect 14288 13076 14352 13140
rect 14369 13076 14433 13140
rect 14451 13076 14515 13140
rect 14533 13076 14597 13140
rect 14615 13076 14679 13140
rect 14697 13076 14761 13140
rect 14779 13076 14843 13140
rect 14861 13076 14925 13140
rect 10157 12994 10221 13058
rect 10238 12994 10302 13058
rect 10319 12994 10383 13058
rect 10400 12994 10464 13058
rect 10481 12994 10545 13058
rect 10562 12994 10626 13058
rect 10643 12994 10707 13058
rect 10724 12994 10788 13058
rect 10805 12994 10869 13058
rect 10886 12994 10950 13058
rect 10967 12994 11031 13058
rect 11048 12994 11112 13058
rect 11129 12994 11193 13058
rect 11210 12994 11274 13058
rect 11291 12994 11355 13058
rect 11372 12994 11436 13058
rect 11453 12994 11517 13058
rect 11534 12994 11598 13058
rect 11615 12994 11679 13058
rect 11696 12994 11760 13058
rect 11777 12994 11841 13058
rect 11858 12994 11922 13058
rect 11939 12994 12003 13058
rect 12020 12994 12084 13058
rect 12101 12994 12165 13058
rect 12182 12994 12246 13058
rect 12263 12994 12327 13058
rect 12344 12994 12408 13058
rect 12425 12994 12489 13058
rect 12506 12994 12570 13058
rect 12587 12994 12651 13058
rect 12668 12994 12732 13058
rect 12749 12994 12813 13058
rect 12830 12994 12894 13058
rect 12911 12994 12975 13058
rect 12992 12994 13056 13058
rect 13073 12994 13137 13058
rect 13154 12994 13218 13058
rect 13235 12994 13299 13058
rect 13316 12994 13380 13058
rect 13397 12994 13461 13058
rect 13478 12994 13542 13058
rect 13559 12994 13623 13058
rect 13640 12994 13704 13058
rect 13721 12994 13785 13058
rect 13802 12994 13866 13058
rect 13883 12994 13947 13058
rect 13964 12994 14028 13058
rect 14045 12994 14109 13058
rect 14126 12994 14190 13058
rect 14207 12994 14271 13058
rect 14288 12994 14352 13058
rect 14369 12994 14433 13058
rect 14451 12994 14515 13058
rect 14533 12994 14597 13058
rect 14615 12994 14679 13058
rect 14697 12994 14761 13058
rect 14779 12994 14843 13058
rect 14861 12994 14925 13058
rect 10157 12912 10221 12976
rect 10238 12912 10302 12976
rect 10319 12912 10383 12976
rect 10400 12912 10464 12976
rect 10481 12912 10545 12976
rect 10562 12912 10626 12976
rect 10643 12912 10707 12976
rect 10724 12912 10788 12976
rect 10805 12912 10869 12976
rect 10886 12912 10950 12976
rect 10967 12912 11031 12976
rect 11048 12912 11112 12976
rect 11129 12912 11193 12976
rect 11210 12912 11274 12976
rect 11291 12912 11355 12976
rect 11372 12912 11436 12976
rect 11453 12912 11517 12976
rect 11534 12912 11598 12976
rect 11615 12912 11679 12976
rect 11696 12912 11760 12976
rect 11777 12912 11841 12976
rect 11858 12912 11922 12976
rect 11939 12912 12003 12976
rect 12020 12912 12084 12976
rect 12101 12912 12165 12976
rect 12182 12912 12246 12976
rect 12263 12912 12327 12976
rect 12344 12912 12408 12976
rect 12425 12912 12489 12976
rect 12506 12912 12570 12976
rect 12587 12912 12651 12976
rect 12668 12912 12732 12976
rect 12749 12912 12813 12976
rect 12830 12912 12894 12976
rect 12911 12912 12975 12976
rect 12992 12912 13056 12976
rect 13073 12912 13137 12976
rect 13154 12912 13218 12976
rect 13235 12912 13299 12976
rect 13316 12912 13380 12976
rect 13397 12912 13461 12976
rect 13478 12912 13542 12976
rect 13559 12912 13623 12976
rect 13640 12912 13704 12976
rect 13721 12912 13785 12976
rect 13802 12912 13866 12976
rect 13883 12912 13947 12976
rect 13964 12912 14028 12976
rect 14045 12912 14109 12976
rect 14126 12912 14190 12976
rect 14207 12912 14271 12976
rect 14288 12912 14352 12976
rect 14369 12912 14433 12976
rect 14451 12912 14515 12976
rect 14533 12912 14597 12976
rect 14615 12912 14679 12976
rect 14697 12912 14761 12976
rect 14779 12912 14843 12976
rect 14861 12912 14925 12976
rect 10157 12830 10221 12894
rect 10238 12830 10302 12894
rect 10319 12830 10383 12894
rect 10400 12830 10464 12894
rect 10481 12830 10545 12894
rect 10562 12830 10626 12894
rect 10643 12830 10707 12894
rect 10724 12830 10788 12894
rect 10805 12830 10869 12894
rect 10886 12830 10950 12894
rect 10967 12830 11031 12894
rect 11048 12830 11112 12894
rect 11129 12830 11193 12894
rect 11210 12830 11274 12894
rect 11291 12830 11355 12894
rect 11372 12830 11436 12894
rect 11453 12830 11517 12894
rect 11534 12830 11598 12894
rect 11615 12830 11679 12894
rect 11696 12830 11760 12894
rect 11777 12830 11841 12894
rect 11858 12830 11922 12894
rect 11939 12830 12003 12894
rect 12020 12830 12084 12894
rect 12101 12830 12165 12894
rect 12182 12830 12246 12894
rect 12263 12830 12327 12894
rect 12344 12830 12408 12894
rect 12425 12830 12489 12894
rect 12506 12830 12570 12894
rect 12587 12830 12651 12894
rect 12668 12830 12732 12894
rect 12749 12830 12813 12894
rect 12830 12830 12894 12894
rect 12911 12830 12975 12894
rect 12992 12830 13056 12894
rect 13073 12830 13137 12894
rect 13154 12830 13218 12894
rect 13235 12830 13299 12894
rect 13316 12830 13380 12894
rect 13397 12830 13461 12894
rect 13478 12830 13542 12894
rect 13559 12830 13623 12894
rect 13640 12830 13704 12894
rect 13721 12830 13785 12894
rect 13802 12830 13866 12894
rect 13883 12830 13947 12894
rect 13964 12830 14028 12894
rect 14045 12830 14109 12894
rect 14126 12830 14190 12894
rect 14207 12830 14271 12894
rect 14288 12830 14352 12894
rect 14369 12830 14433 12894
rect 14451 12830 14515 12894
rect 14533 12830 14597 12894
rect 14615 12830 14679 12894
rect 14697 12830 14761 12894
rect 14779 12830 14843 12894
rect 14861 12830 14925 12894
rect 10157 12748 10221 12812
rect 10238 12748 10302 12812
rect 10319 12748 10383 12812
rect 10400 12748 10464 12812
rect 10481 12748 10545 12812
rect 10562 12748 10626 12812
rect 10643 12748 10707 12812
rect 10724 12748 10788 12812
rect 10805 12748 10869 12812
rect 10886 12748 10950 12812
rect 10967 12748 11031 12812
rect 11048 12748 11112 12812
rect 11129 12748 11193 12812
rect 11210 12748 11274 12812
rect 11291 12748 11355 12812
rect 11372 12748 11436 12812
rect 11453 12748 11517 12812
rect 11534 12748 11598 12812
rect 11615 12748 11679 12812
rect 11696 12748 11760 12812
rect 11777 12748 11841 12812
rect 11858 12748 11922 12812
rect 11939 12748 12003 12812
rect 12020 12748 12084 12812
rect 12101 12748 12165 12812
rect 12182 12748 12246 12812
rect 12263 12748 12327 12812
rect 12344 12748 12408 12812
rect 12425 12748 12489 12812
rect 12506 12748 12570 12812
rect 12587 12748 12651 12812
rect 12668 12748 12732 12812
rect 12749 12748 12813 12812
rect 12830 12748 12894 12812
rect 12911 12748 12975 12812
rect 12992 12748 13056 12812
rect 13073 12748 13137 12812
rect 13154 12748 13218 12812
rect 13235 12748 13299 12812
rect 13316 12748 13380 12812
rect 13397 12748 13461 12812
rect 13478 12748 13542 12812
rect 13559 12748 13623 12812
rect 13640 12748 13704 12812
rect 13721 12748 13785 12812
rect 13802 12748 13866 12812
rect 13883 12748 13947 12812
rect 13964 12748 14028 12812
rect 14045 12748 14109 12812
rect 14126 12748 14190 12812
rect 14207 12748 14271 12812
rect 14288 12748 14352 12812
rect 14369 12748 14433 12812
rect 14451 12748 14515 12812
rect 14533 12748 14597 12812
rect 14615 12748 14679 12812
rect 14697 12748 14761 12812
rect 14779 12748 14843 12812
rect 14861 12748 14925 12812
rect 10157 12666 10221 12730
rect 10238 12666 10302 12730
rect 10319 12666 10383 12730
rect 10400 12666 10464 12730
rect 10481 12666 10545 12730
rect 10562 12666 10626 12730
rect 10643 12666 10707 12730
rect 10724 12666 10788 12730
rect 10805 12666 10869 12730
rect 10886 12666 10950 12730
rect 10967 12666 11031 12730
rect 11048 12666 11112 12730
rect 11129 12666 11193 12730
rect 11210 12666 11274 12730
rect 11291 12666 11355 12730
rect 11372 12666 11436 12730
rect 11453 12666 11517 12730
rect 11534 12666 11598 12730
rect 11615 12666 11679 12730
rect 11696 12666 11760 12730
rect 11777 12666 11841 12730
rect 11858 12666 11922 12730
rect 11939 12666 12003 12730
rect 12020 12666 12084 12730
rect 12101 12666 12165 12730
rect 12182 12666 12246 12730
rect 12263 12666 12327 12730
rect 12344 12666 12408 12730
rect 12425 12666 12489 12730
rect 12506 12666 12570 12730
rect 12587 12666 12651 12730
rect 12668 12666 12732 12730
rect 12749 12666 12813 12730
rect 12830 12666 12894 12730
rect 12911 12666 12975 12730
rect 12992 12666 13056 12730
rect 13073 12666 13137 12730
rect 13154 12666 13218 12730
rect 13235 12666 13299 12730
rect 13316 12666 13380 12730
rect 13397 12666 13461 12730
rect 13478 12666 13542 12730
rect 13559 12666 13623 12730
rect 13640 12666 13704 12730
rect 13721 12666 13785 12730
rect 13802 12666 13866 12730
rect 13883 12666 13947 12730
rect 13964 12666 14028 12730
rect 14045 12666 14109 12730
rect 14126 12666 14190 12730
rect 14207 12666 14271 12730
rect 14288 12666 14352 12730
rect 14369 12666 14433 12730
rect 14451 12666 14515 12730
rect 14533 12666 14597 12730
rect 14615 12666 14679 12730
rect 14697 12666 14761 12730
rect 14779 12666 14843 12730
rect 14861 12666 14925 12730
rect 10157 12584 10221 12648
rect 10238 12584 10302 12648
rect 10319 12584 10383 12648
rect 10400 12584 10464 12648
rect 10481 12584 10545 12648
rect 10562 12584 10626 12648
rect 10643 12584 10707 12648
rect 10724 12584 10788 12648
rect 10805 12584 10869 12648
rect 10886 12584 10950 12648
rect 10967 12584 11031 12648
rect 11048 12584 11112 12648
rect 11129 12584 11193 12648
rect 11210 12584 11274 12648
rect 11291 12584 11355 12648
rect 11372 12584 11436 12648
rect 11453 12584 11517 12648
rect 11534 12584 11598 12648
rect 11615 12584 11679 12648
rect 11696 12584 11760 12648
rect 11777 12584 11841 12648
rect 11858 12584 11922 12648
rect 11939 12584 12003 12648
rect 12020 12584 12084 12648
rect 12101 12584 12165 12648
rect 12182 12584 12246 12648
rect 12263 12584 12327 12648
rect 12344 12584 12408 12648
rect 12425 12584 12489 12648
rect 12506 12584 12570 12648
rect 12587 12584 12651 12648
rect 12668 12584 12732 12648
rect 12749 12584 12813 12648
rect 12830 12584 12894 12648
rect 12911 12584 12975 12648
rect 12992 12584 13056 12648
rect 13073 12584 13137 12648
rect 13154 12584 13218 12648
rect 13235 12584 13299 12648
rect 13316 12584 13380 12648
rect 13397 12584 13461 12648
rect 13478 12584 13542 12648
rect 13559 12584 13623 12648
rect 13640 12584 13704 12648
rect 13721 12584 13785 12648
rect 13802 12584 13866 12648
rect 13883 12584 13947 12648
rect 13964 12584 14028 12648
rect 14045 12584 14109 12648
rect 14126 12584 14190 12648
rect 14207 12584 14271 12648
rect 14288 12584 14352 12648
rect 14369 12584 14433 12648
rect 14451 12584 14515 12648
rect 14533 12584 14597 12648
rect 14615 12584 14679 12648
rect 14697 12584 14761 12648
rect 14779 12584 14843 12648
rect 14861 12584 14925 12648
rect 10157 12502 10221 12566
rect 10238 12502 10302 12566
rect 10319 12502 10383 12566
rect 10400 12502 10464 12566
rect 10481 12502 10545 12566
rect 10562 12502 10626 12566
rect 10643 12502 10707 12566
rect 10724 12502 10788 12566
rect 10805 12502 10869 12566
rect 10886 12502 10950 12566
rect 10967 12502 11031 12566
rect 11048 12502 11112 12566
rect 11129 12502 11193 12566
rect 11210 12502 11274 12566
rect 11291 12502 11355 12566
rect 11372 12502 11436 12566
rect 11453 12502 11517 12566
rect 11534 12502 11598 12566
rect 11615 12502 11679 12566
rect 11696 12502 11760 12566
rect 11777 12502 11841 12566
rect 11858 12502 11922 12566
rect 11939 12502 12003 12566
rect 12020 12502 12084 12566
rect 12101 12502 12165 12566
rect 12182 12502 12246 12566
rect 12263 12502 12327 12566
rect 12344 12502 12408 12566
rect 12425 12502 12489 12566
rect 12506 12502 12570 12566
rect 12587 12502 12651 12566
rect 12668 12502 12732 12566
rect 12749 12502 12813 12566
rect 12830 12502 12894 12566
rect 12911 12502 12975 12566
rect 12992 12502 13056 12566
rect 13073 12502 13137 12566
rect 13154 12502 13218 12566
rect 13235 12502 13299 12566
rect 13316 12502 13380 12566
rect 13397 12502 13461 12566
rect 13478 12502 13542 12566
rect 13559 12502 13623 12566
rect 13640 12502 13704 12566
rect 13721 12502 13785 12566
rect 13802 12502 13866 12566
rect 13883 12502 13947 12566
rect 13964 12502 14028 12566
rect 14045 12502 14109 12566
rect 14126 12502 14190 12566
rect 14207 12502 14271 12566
rect 14288 12502 14352 12566
rect 14369 12502 14433 12566
rect 14451 12502 14515 12566
rect 14533 12502 14597 12566
rect 14615 12502 14679 12566
rect 14697 12502 14761 12566
rect 14779 12502 14843 12566
rect 14861 12502 14925 12566
rect 10157 12420 10221 12484
rect 10238 12420 10302 12484
rect 10319 12420 10383 12484
rect 10400 12420 10464 12484
rect 10481 12420 10545 12484
rect 10562 12420 10626 12484
rect 10643 12420 10707 12484
rect 10724 12420 10788 12484
rect 10805 12420 10869 12484
rect 10886 12420 10950 12484
rect 10967 12420 11031 12484
rect 11048 12420 11112 12484
rect 11129 12420 11193 12484
rect 11210 12420 11274 12484
rect 11291 12420 11355 12484
rect 11372 12420 11436 12484
rect 11453 12420 11517 12484
rect 11534 12420 11598 12484
rect 11615 12420 11679 12484
rect 11696 12420 11760 12484
rect 11777 12420 11841 12484
rect 11858 12420 11922 12484
rect 11939 12420 12003 12484
rect 12020 12420 12084 12484
rect 12101 12420 12165 12484
rect 12182 12420 12246 12484
rect 12263 12420 12327 12484
rect 12344 12420 12408 12484
rect 12425 12420 12489 12484
rect 12506 12420 12570 12484
rect 12587 12420 12651 12484
rect 12668 12420 12732 12484
rect 12749 12420 12813 12484
rect 12830 12420 12894 12484
rect 12911 12420 12975 12484
rect 12992 12420 13056 12484
rect 13073 12420 13137 12484
rect 13154 12420 13218 12484
rect 13235 12420 13299 12484
rect 13316 12420 13380 12484
rect 13397 12420 13461 12484
rect 13478 12420 13542 12484
rect 13559 12420 13623 12484
rect 13640 12420 13704 12484
rect 13721 12420 13785 12484
rect 13802 12420 13866 12484
rect 13883 12420 13947 12484
rect 13964 12420 14028 12484
rect 14045 12420 14109 12484
rect 14126 12420 14190 12484
rect 14207 12420 14271 12484
rect 14288 12420 14352 12484
rect 14369 12420 14433 12484
rect 14451 12420 14515 12484
rect 14533 12420 14597 12484
rect 14615 12420 14679 12484
rect 14697 12420 14761 12484
rect 14779 12420 14843 12484
rect 14861 12420 14925 12484
rect 126 4420 190 4484
rect 207 4420 271 4484
rect 288 4420 352 4484
rect 369 4420 433 4484
rect 450 4420 514 4484
rect 531 4420 595 4484
rect 612 4420 676 4484
rect 693 4420 757 4484
rect 774 4420 838 4484
rect 855 4420 919 4484
rect 936 4420 1000 4484
rect 1017 4420 1081 4484
rect 1098 4420 1162 4484
rect 1179 4420 1243 4484
rect 1260 4420 1324 4484
rect 1341 4420 1405 4484
rect 1422 4420 1486 4484
rect 1503 4420 1567 4484
rect 1584 4420 1648 4484
rect 1665 4420 1729 4484
rect 1746 4420 1810 4484
rect 1827 4420 1891 4484
rect 1908 4420 1972 4484
rect 1989 4420 2053 4484
rect 2070 4420 2134 4484
rect 2151 4420 2215 4484
rect 2232 4420 2296 4484
rect 2313 4420 2377 4484
rect 2394 4420 2458 4484
rect 2475 4420 2539 4484
rect 2556 4420 2620 4484
rect 2637 4420 2701 4484
rect 2718 4420 2782 4484
rect 2799 4420 2863 4484
rect 2880 4420 2944 4484
rect 2961 4420 3025 4484
rect 3042 4420 3106 4484
rect 3123 4420 3187 4484
rect 3204 4420 3268 4484
rect 3285 4420 3349 4484
rect 3366 4420 3430 4484
rect 3447 4420 3511 4484
rect 3528 4420 3592 4484
rect 3609 4420 3673 4484
rect 3690 4420 3754 4484
rect 3771 4420 3835 4484
rect 3852 4420 3916 4484
rect 3933 4420 3997 4484
rect 4014 4420 4078 4484
rect 4095 4420 4159 4484
rect 4176 4420 4240 4484
rect 4257 4420 4321 4484
rect 4338 4420 4402 4484
rect 4420 4420 4484 4484
rect 4502 4420 4566 4484
rect 4584 4420 4648 4484
rect 4666 4420 4730 4484
rect 4748 4420 4812 4484
rect 4830 4420 4894 4484
rect 126 4334 190 4398
rect 207 4334 271 4398
rect 288 4334 352 4398
rect 369 4334 433 4398
rect 450 4334 514 4398
rect 531 4334 595 4398
rect 612 4334 676 4398
rect 693 4334 757 4398
rect 774 4334 838 4398
rect 855 4334 919 4398
rect 936 4334 1000 4398
rect 1017 4334 1081 4398
rect 1098 4334 1162 4398
rect 1179 4334 1243 4398
rect 1260 4334 1324 4398
rect 1341 4334 1405 4398
rect 1422 4334 1486 4398
rect 1503 4334 1567 4398
rect 1584 4334 1648 4398
rect 1665 4334 1729 4398
rect 1746 4334 1810 4398
rect 1827 4334 1891 4398
rect 1908 4334 1972 4398
rect 1989 4334 2053 4398
rect 2070 4334 2134 4398
rect 2151 4334 2215 4398
rect 2232 4334 2296 4398
rect 2313 4334 2377 4398
rect 2394 4334 2458 4398
rect 2475 4334 2539 4398
rect 2556 4334 2620 4398
rect 2637 4334 2701 4398
rect 2718 4334 2782 4398
rect 2799 4334 2863 4398
rect 2880 4334 2944 4398
rect 2961 4334 3025 4398
rect 3042 4334 3106 4398
rect 3123 4334 3187 4398
rect 3204 4334 3268 4398
rect 3285 4334 3349 4398
rect 3366 4334 3430 4398
rect 3447 4334 3511 4398
rect 3528 4334 3592 4398
rect 3609 4334 3673 4398
rect 3690 4334 3754 4398
rect 3771 4334 3835 4398
rect 3852 4334 3916 4398
rect 3933 4334 3997 4398
rect 4014 4334 4078 4398
rect 4095 4334 4159 4398
rect 4176 4334 4240 4398
rect 4257 4334 4321 4398
rect 4338 4334 4402 4398
rect 4420 4334 4484 4398
rect 4502 4334 4566 4398
rect 4584 4334 4648 4398
rect 4666 4334 4730 4398
rect 4748 4334 4812 4398
rect 4830 4334 4894 4398
rect 126 4248 190 4312
rect 207 4248 271 4312
rect 288 4248 352 4312
rect 369 4248 433 4312
rect 450 4248 514 4312
rect 531 4248 595 4312
rect 612 4248 676 4312
rect 693 4248 757 4312
rect 774 4248 838 4312
rect 855 4248 919 4312
rect 936 4248 1000 4312
rect 1017 4248 1081 4312
rect 1098 4248 1162 4312
rect 1179 4248 1243 4312
rect 1260 4248 1324 4312
rect 1341 4248 1405 4312
rect 1422 4248 1486 4312
rect 1503 4248 1567 4312
rect 1584 4248 1648 4312
rect 1665 4248 1729 4312
rect 1746 4248 1810 4312
rect 1827 4248 1891 4312
rect 1908 4248 1972 4312
rect 1989 4248 2053 4312
rect 2070 4248 2134 4312
rect 2151 4248 2215 4312
rect 2232 4248 2296 4312
rect 2313 4248 2377 4312
rect 2394 4248 2458 4312
rect 2475 4248 2539 4312
rect 2556 4248 2620 4312
rect 2637 4248 2701 4312
rect 2718 4248 2782 4312
rect 2799 4248 2863 4312
rect 2880 4248 2944 4312
rect 2961 4248 3025 4312
rect 3042 4248 3106 4312
rect 3123 4248 3187 4312
rect 3204 4248 3268 4312
rect 3285 4248 3349 4312
rect 3366 4248 3430 4312
rect 3447 4248 3511 4312
rect 3528 4248 3592 4312
rect 3609 4248 3673 4312
rect 3690 4248 3754 4312
rect 3771 4248 3835 4312
rect 3852 4248 3916 4312
rect 3933 4248 3997 4312
rect 4014 4248 4078 4312
rect 4095 4248 4159 4312
rect 4176 4248 4240 4312
rect 4257 4248 4321 4312
rect 4338 4248 4402 4312
rect 4420 4248 4484 4312
rect 4502 4248 4566 4312
rect 4584 4248 4648 4312
rect 4666 4248 4730 4312
rect 4748 4248 4812 4312
rect 4830 4248 4894 4312
rect 126 4162 190 4226
rect 207 4162 271 4226
rect 288 4162 352 4226
rect 369 4162 433 4226
rect 450 4162 514 4226
rect 531 4162 595 4226
rect 612 4162 676 4226
rect 693 4162 757 4226
rect 774 4162 838 4226
rect 855 4162 919 4226
rect 936 4162 1000 4226
rect 1017 4162 1081 4226
rect 1098 4162 1162 4226
rect 1179 4162 1243 4226
rect 1260 4162 1324 4226
rect 1341 4162 1405 4226
rect 1422 4162 1486 4226
rect 1503 4162 1567 4226
rect 1584 4162 1648 4226
rect 1665 4162 1729 4226
rect 1746 4162 1810 4226
rect 1827 4162 1891 4226
rect 1908 4162 1972 4226
rect 1989 4162 2053 4226
rect 2070 4162 2134 4226
rect 2151 4162 2215 4226
rect 2232 4162 2296 4226
rect 2313 4162 2377 4226
rect 2394 4162 2458 4226
rect 2475 4162 2539 4226
rect 2556 4162 2620 4226
rect 2637 4162 2701 4226
rect 2718 4162 2782 4226
rect 2799 4162 2863 4226
rect 2880 4162 2944 4226
rect 2961 4162 3025 4226
rect 3042 4162 3106 4226
rect 3123 4162 3187 4226
rect 3204 4162 3268 4226
rect 3285 4162 3349 4226
rect 3366 4162 3430 4226
rect 3447 4162 3511 4226
rect 3528 4162 3592 4226
rect 3609 4162 3673 4226
rect 3690 4162 3754 4226
rect 3771 4162 3835 4226
rect 3852 4162 3916 4226
rect 3933 4162 3997 4226
rect 4014 4162 4078 4226
rect 4095 4162 4159 4226
rect 4176 4162 4240 4226
rect 4257 4162 4321 4226
rect 4338 4162 4402 4226
rect 4420 4162 4484 4226
rect 4502 4162 4566 4226
rect 4584 4162 4648 4226
rect 4666 4162 4730 4226
rect 4748 4162 4812 4226
rect 4830 4162 4894 4226
rect 126 4076 190 4140
rect 207 4076 271 4140
rect 288 4076 352 4140
rect 369 4076 433 4140
rect 450 4076 514 4140
rect 531 4076 595 4140
rect 612 4076 676 4140
rect 693 4076 757 4140
rect 774 4076 838 4140
rect 855 4076 919 4140
rect 936 4076 1000 4140
rect 1017 4076 1081 4140
rect 1098 4076 1162 4140
rect 1179 4076 1243 4140
rect 1260 4076 1324 4140
rect 1341 4076 1405 4140
rect 1422 4076 1486 4140
rect 1503 4076 1567 4140
rect 1584 4076 1648 4140
rect 1665 4076 1729 4140
rect 1746 4076 1810 4140
rect 1827 4076 1891 4140
rect 1908 4076 1972 4140
rect 1989 4076 2053 4140
rect 2070 4076 2134 4140
rect 2151 4076 2215 4140
rect 2232 4076 2296 4140
rect 2313 4076 2377 4140
rect 2394 4076 2458 4140
rect 2475 4076 2539 4140
rect 2556 4076 2620 4140
rect 2637 4076 2701 4140
rect 2718 4076 2782 4140
rect 2799 4076 2863 4140
rect 2880 4076 2944 4140
rect 2961 4076 3025 4140
rect 3042 4076 3106 4140
rect 3123 4076 3187 4140
rect 3204 4076 3268 4140
rect 3285 4076 3349 4140
rect 3366 4076 3430 4140
rect 3447 4076 3511 4140
rect 3528 4076 3592 4140
rect 3609 4076 3673 4140
rect 3690 4076 3754 4140
rect 3771 4076 3835 4140
rect 3852 4076 3916 4140
rect 3933 4076 3997 4140
rect 4014 4076 4078 4140
rect 4095 4076 4159 4140
rect 4176 4076 4240 4140
rect 4257 4076 4321 4140
rect 4338 4076 4402 4140
rect 4420 4076 4484 4140
rect 4502 4076 4566 4140
rect 4584 4076 4648 4140
rect 4666 4076 4730 4140
rect 4748 4076 4812 4140
rect 4830 4076 4894 4140
rect 126 3990 190 4054
rect 207 3990 271 4054
rect 288 3990 352 4054
rect 369 3990 433 4054
rect 450 3990 514 4054
rect 531 3990 595 4054
rect 612 3990 676 4054
rect 693 3990 757 4054
rect 774 3990 838 4054
rect 855 3990 919 4054
rect 936 3990 1000 4054
rect 1017 3990 1081 4054
rect 1098 3990 1162 4054
rect 1179 3990 1243 4054
rect 1260 3990 1324 4054
rect 1341 3990 1405 4054
rect 1422 3990 1486 4054
rect 1503 3990 1567 4054
rect 1584 3990 1648 4054
rect 1665 3990 1729 4054
rect 1746 3990 1810 4054
rect 1827 3990 1891 4054
rect 1908 3990 1972 4054
rect 1989 3990 2053 4054
rect 2070 3990 2134 4054
rect 2151 3990 2215 4054
rect 2232 3990 2296 4054
rect 2313 3990 2377 4054
rect 2394 3990 2458 4054
rect 2475 3990 2539 4054
rect 2556 3990 2620 4054
rect 2637 3990 2701 4054
rect 2718 3990 2782 4054
rect 2799 3990 2863 4054
rect 2880 3990 2944 4054
rect 2961 3990 3025 4054
rect 3042 3990 3106 4054
rect 3123 3990 3187 4054
rect 3204 3990 3268 4054
rect 3285 3990 3349 4054
rect 3366 3990 3430 4054
rect 3447 3990 3511 4054
rect 3528 3990 3592 4054
rect 3609 3990 3673 4054
rect 3690 3990 3754 4054
rect 3771 3990 3835 4054
rect 3852 3990 3916 4054
rect 3933 3990 3997 4054
rect 4014 3990 4078 4054
rect 4095 3990 4159 4054
rect 4176 3990 4240 4054
rect 4257 3990 4321 4054
rect 4338 3990 4402 4054
rect 4420 3990 4484 4054
rect 4502 3990 4566 4054
rect 4584 3990 4648 4054
rect 4666 3990 4730 4054
rect 4748 3990 4812 4054
rect 4830 3990 4894 4054
rect 126 3904 190 3968
rect 207 3904 271 3968
rect 288 3904 352 3968
rect 369 3904 433 3968
rect 450 3904 514 3968
rect 531 3904 595 3968
rect 612 3904 676 3968
rect 693 3904 757 3968
rect 774 3904 838 3968
rect 855 3904 919 3968
rect 936 3904 1000 3968
rect 1017 3904 1081 3968
rect 1098 3904 1162 3968
rect 1179 3904 1243 3968
rect 1260 3904 1324 3968
rect 1341 3904 1405 3968
rect 1422 3904 1486 3968
rect 1503 3904 1567 3968
rect 1584 3904 1648 3968
rect 1665 3904 1729 3968
rect 1746 3904 1810 3968
rect 1827 3904 1891 3968
rect 1908 3904 1972 3968
rect 1989 3904 2053 3968
rect 2070 3904 2134 3968
rect 2151 3904 2215 3968
rect 2232 3904 2296 3968
rect 2313 3904 2377 3968
rect 2394 3904 2458 3968
rect 2475 3904 2539 3968
rect 2556 3904 2620 3968
rect 2637 3904 2701 3968
rect 2718 3904 2782 3968
rect 2799 3904 2863 3968
rect 2880 3904 2944 3968
rect 2961 3904 3025 3968
rect 3042 3904 3106 3968
rect 3123 3904 3187 3968
rect 3204 3904 3268 3968
rect 3285 3904 3349 3968
rect 3366 3904 3430 3968
rect 3447 3904 3511 3968
rect 3528 3904 3592 3968
rect 3609 3904 3673 3968
rect 3690 3904 3754 3968
rect 3771 3904 3835 3968
rect 3852 3904 3916 3968
rect 3933 3904 3997 3968
rect 4014 3904 4078 3968
rect 4095 3904 4159 3968
rect 4176 3904 4240 3968
rect 4257 3904 4321 3968
rect 4338 3904 4402 3968
rect 4420 3904 4484 3968
rect 4502 3904 4566 3968
rect 4584 3904 4648 3968
rect 4666 3904 4730 3968
rect 4748 3904 4812 3968
rect 4830 3904 4894 3968
rect 126 3818 190 3882
rect 207 3818 271 3882
rect 288 3818 352 3882
rect 369 3818 433 3882
rect 450 3818 514 3882
rect 531 3818 595 3882
rect 612 3818 676 3882
rect 693 3818 757 3882
rect 774 3818 838 3882
rect 855 3818 919 3882
rect 936 3818 1000 3882
rect 1017 3818 1081 3882
rect 1098 3818 1162 3882
rect 1179 3818 1243 3882
rect 1260 3818 1324 3882
rect 1341 3818 1405 3882
rect 1422 3818 1486 3882
rect 1503 3818 1567 3882
rect 1584 3818 1648 3882
rect 1665 3818 1729 3882
rect 1746 3818 1810 3882
rect 1827 3818 1891 3882
rect 1908 3818 1972 3882
rect 1989 3818 2053 3882
rect 2070 3818 2134 3882
rect 2151 3818 2215 3882
rect 2232 3818 2296 3882
rect 2313 3818 2377 3882
rect 2394 3818 2458 3882
rect 2475 3818 2539 3882
rect 2556 3818 2620 3882
rect 2637 3818 2701 3882
rect 2718 3818 2782 3882
rect 2799 3818 2863 3882
rect 2880 3818 2944 3882
rect 2961 3818 3025 3882
rect 3042 3818 3106 3882
rect 3123 3818 3187 3882
rect 3204 3818 3268 3882
rect 3285 3818 3349 3882
rect 3366 3818 3430 3882
rect 3447 3818 3511 3882
rect 3528 3818 3592 3882
rect 3609 3818 3673 3882
rect 3690 3818 3754 3882
rect 3771 3818 3835 3882
rect 3852 3818 3916 3882
rect 3933 3818 3997 3882
rect 4014 3818 4078 3882
rect 4095 3818 4159 3882
rect 4176 3818 4240 3882
rect 4257 3818 4321 3882
rect 4338 3818 4402 3882
rect 4420 3818 4484 3882
rect 4502 3818 4566 3882
rect 4584 3818 4648 3882
rect 4666 3818 4730 3882
rect 4748 3818 4812 3882
rect 4830 3818 4894 3882
rect 126 3732 190 3796
rect 207 3732 271 3796
rect 288 3732 352 3796
rect 369 3732 433 3796
rect 450 3732 514 3796
rect 531 3732 595 3796
rect 612 3732 676 3796
rect 693 3732 757 3796
rect 774 3732 838 3796
rect 855 3732 919 3796
rect 936 3732 1000 3796
rect 1017 3732 1081 3796
rect 1098 3732 1162 3796
rect 1179 3732 1243 3796
rect 1260 3732 1324 3796
rect 1341 3732 1405 3796
rect 1422 3732 1486 3796
rect 1503 3732 1567 3796
rect 1584 3732 1648 3796
rect 1665 3732 1729 3796
rect 1746 3732 1810 3796
rect 1827 3732 1891 3796
rect 1908 3732 1972 3796
rect 1989 3732 2053 3796
rect 2070 3732 2134 3796
rect 2151 3732 2215 3796
rect 2232 3732 2296 3796
rect 2313 3732 2377 3796
rect 2394 3732 2458 3796
rect 2475 3732 2539 3796
rect 2556 3732 2620 3796
rect 2637 3732 2701 3796
rect 2718 3732 2782 3796
rect 2799 3732 2863 3796
rect 2880 3732 2944 3796
rect 2961 3732 3025 3796
rect 3042 3732 3106 3796
rect 3123 3732 3187 3796
rect 3204 3732 3268 3796
rect 3285 3732 3349 3796
rect 3366 3732 3430 3796
rect 3447 3732 3511 3796
rect 3528 3732 3592 3796
rect 3609 3732 3673 3796
rect 3690 3732 3754 3796
rect 3771 3732 3835 3796
rect 3852 3732 3916 3796
rect 3933 3732 3997 3796
rect 4014 3732 4078 3796
rect 4095 3732 4159 3796
rect 4176 3732 4240 3796
rect 4257 3732 4321 3796
rect 4338 3732 4402 3796
rect 4420 3732 4484 3796
rect 4502 3732 4566 3796
rect 4584 3732 4648 3796
rect 4666 3732 4730 3796
rect 4748 3732 4812 3796
rect 4830 3732 4894 3796
rect 126 3646 190 3710
rect 207 3646 271 3710
rect 288 3646 352 3710
rect 369 3646 433 3710
rect 450 3646 514 3710
rect 531 3646 595 3710
rect 612 3646 676 3710
rect 693 3646 757 3710
rect 774 3646 838 3710
rect 855 3646 919 3710
rect 936 3646 1000 3710
rect 1017 3646 1081 3710
rect 1098 3646 1162 3710
rect 1179 3646 1243 3710
rect 1260 3646 1324 3710
rect 1341 3646 1405 3710
rect 1422 3646 1486 3710
rect 1503 3646 1567 3710
rect 1584 3646 1648 3710
rect 1665 3646 1729 3710
rect 1746 3646 1810 3710
rect 1827 3646 1891 3710
rect 1908 3646 1972 3710
rect 1989 3646 2053 3710
rect 2070 3646 2134 3710
rect 2151 3646 2215 3710
rect 2232 3646 2296 3710
rect 2313 3646 2377 3710
rect 2394 3646 2458 3710
rect 2475 3646 2539 3710
rect 2556 3646 2620 3710
rect 2637 3646 2701 3710
rect 2718 3646 2782 3710
rect 2799 3646 2863 3710
rect 2880 3646 2944 3710
rect 2961 3646 3025 3710
rect 3042 3646 3106 3710
rect 3123 3646 3187 3710
rect 3204 3646 3268 3710
rect 3285 3646 3349 3710
rect 3366 3646 3430 3710
rect 3447 3646 3511 3710
rect 3528 3646 3592 3710
rect 3609 3646 3673 3710
rect 3690 3646 3754 3710
rect 3771 3646 3835 3710
rect 3852 3646 3916 3710
rect 3933 3646 3997 3710
rect 4014 3646 4078 3710
rect 4095 3646 4159 3710
rect 4176 3646 4240 3710
rect 4257 3646 4321 3710
rect 4338 3646 4402 3710
rect 4420 3646 4484 3710
rect 4502 3646 4566 3710
rect 4584 3646 4648 3710
rect 4666 3646 4730 3710
rect 4748 3646 4812 3710
rect 4830 3646 4894 3710
rect 126 3560 190 3624
rect 207 3560 271 3624
rect 288 3560 352 3624
rect 369 3560 433 3624
rect 450 3560 514 3624
rect 531 3560 595 3624
rect 612 3560 676 3624
rect 693 3560 757 3624
rect 774 3560 838 3624
rect 855 3560 919 3624
rect 936 3560 1000 3624
rect 1017 3560 1081 3624
rect 1098 3560 1162 3624
rect 1179 3560 1243 3624
rect 1260 3560 1324 3624
rect 1341 3560 1405 3624
rect 1422 3560 1486 3624
rect 1503 3560 1567 3624
rect 1584 3560 1648 3624
rect 1665 3560 1729 3624
rect 1746 3560 1810 3624
rect 1827 3560 1891 3624
rect 1908 3560 1972 3624
rect 1989 3560 2053 3624
rect 2070 3560 2134 3624
rect 2151 3560 2215 3624
rect 2232 3560 2296 3624
rect 2313 3560 2377 3624
rect 2394 3560 2458 3624
rect 2475 3560 2539 3624
rect 2556 3560 2620 3624
rect 2637 3560 2701 3624
rect 2718 3560 2782 3624
rect 2799 3560 2863 3624
rect 2880 3560 2944 3624
rect 2961 3560 3025 3624
rect 3042 3560 3106 3624
rect 3123 3560 3187 3624
rect 3204 3560 3268 3624
rect 3285 3560 3349 3624
rect 3366 3560 3430 3624
rect 3447 3560 3511 3624
rect 3528 3560 3592 3624
rect 3609 3560 3673 3624
rect 3690 3560 3754 3624
rect 3771 3560 3835 3624
rect 3852 3560 3916 3624
rect 3933 3560 3997 3624
rect 4014 3560 4078 3624
rect 4095 3560 4159 3624
rect 4176 3560 4240 3624
rect 4257 3560 4321 3624
rect 4338 3560 4402 3624
rect 4420 3560 4484 3624
rect 4502 3560 4566 3624
rect 4584 3560 4648 3624
rect 4666 3560 4730 3624
rect 4748 3560 4812 3624
rect 4830 3560 4894 3624
rect 10157 4420 10221 4484
rect 10238 4420 10302 4484
rect 10319 4420 10383 4484
rect 10400 4420 10464 4484
rect 10481 4420 10545 4484
rect 10562 4420 10626 4484
rect 10643 4420 10707 4484
rect 10724 4420 10788 4484
rect 10805 4420 10869 4484
rect 10886 4420 10950 4484
rect 10967 4420 11031 4484
rect 11048 4420 11112 4484
rect 11129 4420 11193 4484
rect 11210 4420 11274 4484
rect 11291 4420 11355 4484
rect 11372 4420 11436 4484
rect 11453 4420 11517 4484
rect 11534 4420 11598 4484
rect 11615 4420 11679 4484
rect 11696 4420 11760 4484
rect 11777 4420 11841 4484
rect 11858 4420 11922 4484
rect 11939 4420 12003 4484
rect 12020 4420 12084 4484
rect 12101 4420 12165 4484
rect 12182 4420 12246 4484
rect 12263 4420 12327 4484
rect 12344 4420 12408 4484
rect 12425 4420 12489 4484
rect 12506 4420 12570 4484
rect 12587 4420 12651 4484
rect 12668 4420 12732 4484
rect 12749 4420 12813 4484
rect 12830 4420 12894 4484
rect 12911 4420 12975 4484
rect 12992 4420 13056 4484
rect 13073 4420 13137 4484
rect 13154 4420 13218 4484
rect 13235 4420 13299 4484
rect 13316 4420 13380 4484
rect 13397 4420 13461 4484
rect 13478 4420 13542 4484
rect 13559 4420 13623 4484
rect 13640 4420 13704 4484
rect 13721 4420 13785 4484
rect 13802 4420 13866 4484
rect 13883 4420 13947 4484
rect 13964 4420 14028 4484
rect 14045 4420 14109 4484
rect 14126 4420 14190 4484
rect 14207 4420 14271 4484
rect 14288 4420 14352 4484
rect 14369 4420 14433 4484
rect 14451 4420 14515 4484
rect 14533 4420 14597 4484
rect 14615 4420 14679 4484
rect 14697 4420 14761 4484
rect 14779 4420 14843 4484
rect 14861 4420 14925 4484
rect 10157 4334 10221 4398
rect 10238 4334 10302 4398
rect 10319 4334 10383 4398
rect 10400 4334 10464 4398
rect 10481 4334 10545 4398
rect 10562 4334 10626 4398
rect 10643 4334 10707 4398
rect 10724 4334 10788 4398
rect 10805 4334 10869 4398
rect 10886 4334 10950 4398
rect 10967 4334 11031 4398
rect 11048 4334 11112 4398
rect 11129 4334 11193 4398
rect 11210 4334 11274 4398
rect 11291 4334 11355 4398
rect 11372 4334 11436 4398
rect 11453 4334 11517 4398
rect 11534 4334 11598 4398
rect 11615 4334 11679 4398
rect 11696 4334 11760 4398
rect 11777 4334 11841 4398
rect 11858 4334 11922 4398
rect 11939 4334 12003 4398
rect 12020 4334 12084 4398
rect 12101 4334 12165 4398
rect 12182 4334 12246 4398
rect 12263 4334 12327 4398
rect 12344 4334 12408 4398
rect 12425 4334 12489 4398
rect 12506 4334 12570 4398
rect 12587 4334 12651 4398
rect 12668 4334 12732 4398
rect 12749 4334 12813 4398
rect 12830 4334 12894 4398
rect 12911 4334 12975 4398
rect 12992 4334 13056 4398
rect 13073 4334 13137 4398
rect 13154 4334 13218 4398
rect 13235 4334 13299 4398
rect 13316 4334 13380 4398
rect 13397 4334 13461 4398
rect 13478 4334 13542 4398
rect 13559 4334 13623 4398
rect 13640 4334 13704 4398
rect 13721 4334 13785 4398
rect 13802 4334 13866 4398
rect 13883 4334 13947 4398
rect 13964 4334 14028 4398
rect 14045 4334 14109 4398
rect 14126 4334 14190 4398
rect 14207 4334 14271 4398
rect 14288 4334 14352 4398
rect 14369 4334 14433 4398
rect 14451 4334 14515 4398
rect 14533 4334 14597 4398
rect 14615 4334 14679 4398
rect 14697 4334 14761 4398
rect 14779 4334 14843 4398
rect 14861 4334 14925 4398
rect 10157 4248 10221 4312
rect 10238 4248 10302 4312
rect 10319 4248 10383 4312
rect 10400 4248 10464 4312
rect 10481 4248 10545 4312
rect 10562 4248 10626 4312
rect 10643 4248 10707 4312
rect 10724 4248 10788 4312
rect 10805 4248 10869 4312
rect 10886 4248 10950 4312
rect 10967 4248 11031 4312
rect 11048 4248 11112 4312
rect 11129 4248 11193 4312
rect 11210 4248 11274 4312
rect 11291 4248 11355 4312
rect 11372 4248 11436 4312
rect 11453 4248 11517 4312
rect 11534 4248 11598 4312
rect 11615 4248 11679 4312
rect 11696 4248 11760 4312
rect 11777 4248 11841 4312
rect 11858 4248 11922 4312
rect 11939 4248 12003 4312
rect 12020 4248 12084 4312
rect 12101 4248 12165 4312
rect 12182 4248 12246 4312
rect 12263 4248 12327 4312
rect 12344 4248 12408 4312
rect 12425 4248 12489 4312
rect 12506 4248 12570 4312
rect 12587 4248 12651 4312
rect 12668 4248 12732 4312
rect 12749 4248 12813 4312
rect 12830 4248 12894 4312
rect 12911 4248 12975 4312
rect 12992 4248 13056 4312
rect 13073 4248 13137 4312
rect 13154 4248 13218 4312
rect 13235 4248 13299 4312
rect 13316 4248 13380 4312
rect 13397 4248 13461 4312
rect 13478 4248 13542 4312
rect 13559 4248 13623 4312
rect 13640 4248 13704 4312
rect 13721 4248 13785 4312
rect 13802 4248 13866 4312
rect 13883 4248 13947 4312
rect 13964 4248 14028 4312
rect 14045 4248 14109 4312
rect 14126 4248 14190 4312
rect 14207 4248 14271 4312
rect 14288 4248 14352 4312
rect 14369 4248 14433 4312
rect 14451 4248 14515 4312
rect 14533 4248 14597 4312
rect 14615 4248 14679 4312
rect 14697 4248 14761 4312
rect 14779 4248 14843 4312
rect 14861 4248 14925 4312
rect 10157 4162 10221 4226
rect 10238 4162 10302 4226
rect 10319 4162 10383 4226
rect 10400 4162 10464 4226
rect 10481 4162 10545 4226
rect 10562 4162 10626 4226
rect 10643 4162 10707 4226
rect 10724 4162 10788 4226
rect 10805 4162 10869 4226
rect 10886 4162 10950 4226
rect 10967 4162 11031 4226
rect 11048 4162 11112 4226
rect 11129 4162 11193 4226
rect 11210 4162 11274 4226
rect 11291 4162 11355 4226
rect 11372 4162 11436 4226
rect 11453 4162 11517 4226
rect 11534 4162 11598 4226
rect 11615 4162 11679 4226
rect 11696 4162 11760 4226
rect 11777 4162 11841 4226
rect 11858 4162 11922 4226
rect 11939 4162 12003 4226
rect 12020 4162 12084 4226
rect 12101 4162 12165 4226
rect 12182 4162 12246 4226
rect 12263 4162 12327 4226
rect 12344 4162 12408 4226
rect 12425 4162 12489 4226
rect 12506 4162 12570 4226
rect 12587 4162 12651 4226
rect 12668 4162 12732 4226
rect 12749 4162 12813 4226
rect 12830 4162 12894 4226
rect 12911 4162 12975 4226
rect 12992 4162 13056 4226
rect 13073 4162 13137 4226
rect 13154 4162 13218 4226
rect 13235 4162 13299 4226
rect 13316 4162 13380 4226
rect 13397 4162 13461 4226
rect 13478 4162 13542 4226
rect 13559 4162 13623 4226
rect 13640 4162 13704 4226
rect 13721 4162 13785 4226
rect 13802 4162 13866 4226
rect 13883 4162 13947 4226
rect 13964 4162 14028 4226
rect 14045 4162 14109 4226
rect 14126 4162 14190 4226
rect 14207 4162 14271 4226
rect 14288 4162 14352 4226
rect 14369 4162 14433 4226
rect 14451 4162 14515 4226
rect 14533 4162 14597 4226
rect 14615 4162 14679 4226
rect 14697 4162 14761 4226
rect 14779 4162 14843 4226
rect 14861 4162 14925 4226
rect 10157 4076 10221 4140
rect 10238 4076 10302 4140
rect 10319 4076 10383 4140
rect 10400 4076 10464 4140
rect 10481 4076 10545 4140
rect 10562 4076 10626 4140
rect 10643 4076 10707 4140
rect 10724 4076 10788 4140
rect 10805 4076 10869 4140
rect 10886 4076 10950 4140
rect 10967 4076 11031 4140
rect 11048 4076 11112 4140
rect 11129 4076 11193 4140
rect 11210 4076 11274 4140
rect 11291 4076 11355 4140
rect 11372 4076 11436 4140
rect 11453 4076 11517 4140
rect 11534 4076 11598 4140
rect 11615 4076 11679 4140
rect 11696 4076 11760 4140
rect 11777 4076 11841 4140
rect 11858 4076 11922 4140
rect 11939 4076 12003 4140
rect 12020 4076 12084 4140
rect 12101 4076 12165 4140
rect 12182 4076 12246 4140
rect 12263 4076 12327 4140
rect 12344 4076 12408 4140
rect 12425 4076 12489 4140
rect 12506 4076 12570 4140
rect 12587 4076 12651 4140
rect 12668 4076 12732 4140
rect 12749 4076 12813 4140
rect 12830 4076 12894 4140
rect 12911 4076 12975 4140
rect 12992 4076 13056 4140
rect 13073 4076 13137 4140
rect 13154 4076 13218 4140
rect 13235 4076 13299 4140
rect 13316 4076 13380 4140
rect 13397 4076 13461 4140
rect 13478 4076 13542 4140
rect 13559 4076 13623 4140
rect 13640 4076 13704 4140
rect 13721 4076 13785 4140
rect 13802 4076 13866 4140
rect 13883 4076 13947 4140
rect 13964 4076 14028 4140
rect 14045 4076 14109 4140
rect 14126 4076 14190 4140
rect 14207 4076 14271 4140
rect 14288 4076 14352 4140
rect 14369 4076 14433 4140
rect 14451 4076 14515 4140
rect 14533 4076 14597 4140
rect 14615 4076 14679 4140
rect 14697 4076 14761 4140
rect 14779 4076 14843 4140
rect 14861 4076 14925 4140
rect 10157 3990 10221 4054
rect 10238 3990 10302 4054
rect 10319 3990 10383 4054
rect 10400 3990 10464 4054
rect 10481 3990 10545 4054
rect 10562 3990 10626 4054
rect 10643 3990 10707 4054
rect 10724 3990 10788 4054
rect 10805 3990 10869 4054
rect 10886 3990 10950 4054
rect 10967 3990 11031 4054
rect 11048 3990 11112 4054
rect 11129 3990 11193 4054
rect 11210 3990 11274 4054
rect 11291 3990 11355 4054
rect 11372 3990 11436 4054
rect 11453 3990 11517 4054
rect 11534 3990 11598 4054
rect 11615 3990 11679 4054
rect 11696 3990 11760 4054
rect 11777 3990 11841 4054
rect 11858 3990 11922 4054
rect 11939 3990 12003 4054
rect 12020 3990 12084 4054
rect 12101 3990 12165 4054
rect 12182 3990 12246 4054
rect 12263 3990 12327 4054
rect 12344 3990 12408 4054
rect 12425 3990 12489 4054
rect 12506 3990 12570 4054
rect 12587 3990 12651 4054
rect 12668 3990 12732 4054
rect 12749 3990 12813 4054
rect 12830 3990 12894 4054
rect 12911 3990 12975 4054
rect 12992 3990 13056 4054
rect 13073 3990 13137 4054
rect 13154 3990 13218 4054
rect 13235 3990 13299 4054
rect 13316 3990 13380 4054
rect 13397 3990 13461 4054
rect 13478 3990 13542 4054
rect 13559 3990 13623 4054
rect 13640 3990 13704 4054
rect 13721 3990 13785 4054
rect 13802 3990 13866 4054
rect 13883 3990 13947 4054
rect 13964 3990 14028 4054
rect 14045 3990 14109 4054
rect 14126 3990 14190 4054
rect 14207 3990 14271 4054
rect 14288 3990 14352 4054
rect 14369 3990 14433 4054
rect 14451 3990 14515 4054
rect 14533 3990 14597 4054
rect 14615 3990 14679 4054
rect 14697 3990 14761 4054
rect 14779 3990 14843 4054
rect 14861 3990 14925 4054
rect 10157 3904 10221 3968
rect 10238 3904 10302 3968
rect 10319 3904 10383 3968
rect 10400 3904 10464 3968
rect 10481 3904 10545 3968
rect 10562 3904 10626 3968
rect 10643 3904 10707 3968
rect 10724 3904 10788 3968
rect 10805 3904 10869 3968
rect 10886 3904 10950 3968
rect 10967 3904 11031 3968
rect 11048 3904 11112 3968
rect 11129 3904 11193 3968
rect 11210 3904 11274 3968
rect 11291 3904 11355 3968
rect 11372 3904 11436 3968
rect 11453 3904 11517 3968
rect 11534 3904 11598 3968
rect 11615 3904 11679 3968
rect 11696 3904 11760 3968
rect 11777 3904 11841 3968
rect 11858 3904 11922 3968
rect 11939 3904 12003 3968
rect 12020 3904 12084 3968
rect 12101 3904 12165 3968
rect 12182 3904 12246 3968
rect 12263 3904 12327 3968
rect 12344 3904 12408 3968
rect 12425 3904 12489 3968
rect 12506 3904 12570 3968
rect 12587 3904 12651 3968
rect 12668 3904 12732 3968
rect 12749 3904 12813 3968
rect 12830 3904 12894 3968
rect 12911 3904 12975 3968
rect 12992 3904 13056 3968
rect 13073 3904 13137 3968
rect 13154 3904 13218 3968
rect 13235 3904 13299 3968
rect 13316 3904 13380 3968
rect 13397 3904 13461 3968
rect 13478 3904 13542 3968
rect 13559 3904 13623 3968
rect 13640 3904 13704 3968
rect 13721 3904 13785 3968
rect 13802 3904 13866 3968
rect 13883 3904 13947 3968
rect 13964 3904 14028 3968
rect 14045 3904 14109 3968
rect 14126 3904 14190 3968
rect 14207 3904 14271 3968
rect 14288 3904 14352 3968
rect 14369 3904 14433 3968
rect 14451 3904 14515 3968
rect 14533 3904 14597 3968
rect 14615 3904 14679 3968
rect 14697 3904 14761 3968
rect 14779 3904 14843 3968
rect 14861 3904 14925 3968
rect 10157 3818 10221 3882
rect 10238 3818 10302 3882
rect 10319 3818 10383 3882
rect 10400 3818 10464 3882
rect 10481 3818 10545 3882
rect 10562 3818 10626 3882
rect 10643 3818 10707 3882
rect 10724 3818 10788 3882
rect 10805 3818 10869 3882
rect 10886 3818 10950 3882
rect 10967 3818 11031 3882
rect 11048 3818 11112 3882
rect 11129 3818 11193 3882
rect 11210 3818 11274 3882
rect 11291 3818 11355 3882
rect 11372 3818 11436 3882
rect 11453 3818 11517 3882
rect 11534 3818 11598 3882
rect 11615 3818 11679 3882
rect 11696 3818 11760 3882
rect 11777 3818 11841 3882
rect 11858 3818 11922 3882
rect 11939 3818 12003 3882
rect 12020 3818 12084 3882
rect 12101 3818 12165 3882
rect 12182 3818 12246 3882
rect 12263 3818 12327 3882
rect 12344 3818 12408 3882
rect 12425 3818 12489 3882
rect 12506 3818 12570 3882
rect 12587 3818 12651 3882
rect 12668 3818 12732 3882
rect 12749 3818 12813 3882
rect 12830 3818 12894 3882
rect 12911 3818 12975 3882
rect 12992 3818 13056 3882
rect 13073 3818 13137 3882
rect 13154 3818 13218 3882
rect 13235 3818 13299 3882
rect 13316 3818 13380 3882
rect 13397 3818 13461 3882
rect 13478 3818 13542 3882
rect 13559 3818 13623 3882
rect 13640 3818 13704 3882
rect 13721 3818 13785 3882
rect 13802 3818 13866 3882
rect 13883 3818 13947 3882
rect 13964 3818 14028 3882
rect 14045 3818 14109 3882
rect 14126 3818 14190 3882
rect 14207 3818 14271 3882
rect 14288 3818 14352 3882
rect 14369 3818 14433 3882
rect 14451 3818 14515 3882
rect 14533 3818 14597 3882
rect 14615 3818 14679 3882
rect 14697 3818 14761 3882
rect 14779 3818 14843 3882
rect 14861 3818 14925 3882
rect 10157 3732 10221 3796
rect 10238 3732 10302 3796
rect 10319 3732 10383 3796
rect 10400 3732 10464 3796
rect 10481 3732 10545 3796
rect 10562 3732 10626 3796
rect 10643 3732 10707 3796
rect 10724 3732 10788 3796
rect 10805 3732 10869 3796
rect 10886 3732 10950 3796
rect 10967 3732 11031 3796
rect 11048 3732 11112 3796
rect 11129 3732 11193 3796
rect 11210 3732 11274 3796
rect 11291 3732 11355 3796
rect 11372 3732 11436 3796
rect 11453 3732 11517 3796
rect 11534 3732 11598 3796
rect 11615 3732 11679 3796
rect 11696 3732 11760 3796
rect 11777 3732 11841 3796
rect 11858 3732 11922 3796
rect 11939 3732 12003 3796
rect 12020 3732 12084 3796
rect 12101 3732 12165 3796
rect 12182 3732 12246 3796
rect 12263 3732 12327 3796
rect 12344 3732 12408 3796
rect 12425 3732 12489 3796
rect 12506 3732 12570 3796
rect 12587 3732 12651 3796
rect 12668 3732 12732 3796
rect 12749 3732 12813 3796
rect 12830 3732 12894 3796
rect 12911 3732 12975 3796
rect 12992 3732 13056 3796
rect 13073 3732 13137 3796
rect 13154 3732 13218 3796
rect 13235 3732 13299 3796
rect 13316 3732 13380 3796
rect 13397 3732 13461 3796
rect 13478 3732 13542 3796
rect 13559 3732 13623 3796
rect 13640 3732 13704 3796
rect 13721 3732 13785 3796
rect 13802 3732 13866 3796
rect 13883 3732 13947 3796
rect 13964 3732 14028 3796
rect 14045 3732 14109 3796
rect 14126 3732 14190 3796
rect 14207 3732 14271 3796
rect 14288 3732 14352 3796
rect 14369 3732 14433 3796
rect 14451 3732 14515 3796
rect 14533 3732 14597 3796
rect 14615 3732 14679 3796
rect 14697 3732 14761 3796
rect 14779 3732 14843 3796
rect 14861 3732 14925 3796
rect 10157 3646 10221 3710
rect 10238 3646 10302 3710
rect 10319 3646 10383 3710
rect 10400 3646 10464 3710
rect 10481 3646 10545 3710
rect 10562 3646 10626 3710
rect 10643 3646 10707 3710
rect 10724 3646 10788 3710
rect 10805 3646 10869 3710
rect 10886 3646 10950 3710
rect 10967 3646 11031 3710
rect 11048 3646 11112 3710
rect 11129 3646 11193 3710
rect 11210 3646 11274 3710
rect 11291 3646 11355 3710
rect 11372 3646 11436 3710
rect 11453 3646 11517 3710
rect 11534 3646 11598 3710
rect 11615 3646 11679 3710
rect 11696 3646 11760 3710
rect 11777 3646 11841 3710
rect 11858 3646 11922 3710
rect 11939 3646 12003 3710
rect 12020 3646 12084 3710
rect 12101 3646 12165 3710
rect 12182 3646 12246 3710
rect 12263 3646 12327 3710
rect 12344 3646 12408 3710
rect 12425 3646 12489 3710
rect 12506 3646 12570 3710
rect 12587 3646 12651 3710
rect 12668 3646 12732 3710
rect 12749 3646 12813 3710
rect 12830 3646 12894 3710
rect 12911 3646 12975 3710
rect 12992 3646 13056 3710
rect 13073 3646 13137 3710
rect 13154 3646 13218 3710
rect 13235 3646 13299 3710
rect 13316 3646 13380 3710
rect 13397 3646 13461 3710
rect 13478 3646 13542 3710
rect 13559 3646 13623 3710
rect 13640 3646 13704 3710
rect 13721 3646 13785 3710
rect 13802 3646 13866 3710
rect 13883 3646 13947 3710
rect 13964 3646 14028 3710
rect 14045 3646 14109 3710
rect 14126 3646 14190 3710
rect 14207 3646 14271 3710
rect 14288 3646 14352 3710
rect 14369 3646 14433 3710
rect 14451 3646 14515 3710
rect 14533 3646 14597 3710
rect 14615 3646 14679 3710
rect 14697 3646 14761 3710
rect 14779 3646 14843 3710
rect 14861 3646 14925 3710
rect 10157 3560 10221 3624
rect 10238 3560 10302 3624
rect 10319 3560 10383 3624
rect 10400 3560 10464 3624
rect 10481 3560 10545 3624
rect 10562 3560 10626 3624
rect 10643 3560 10707 3624
rect 10724 3560 10788 3624
rect 10805 3560 10869 3624
rect 10886 3560 10950 3624
rect 10967 3560 11031 3624
rect 11048 3560 11112 3624
rect 11129 3560 11193 3624
rect 11210 3560 11274 3624
rect 11291 3560 11355 3624
rect 11372 3560 11436 3624
rect 11453 3560 11517 3624
rect 11534 3560 11598 3624
rect 11615 3560 11679 3624
rect 11696 3560 11760 3624
rect 11777 3560 11841 3624
rect 11858 3560 11922 3624
rect 11939 3560 12003 3624
rect 12020 3560 12084 3624
rect 12101 3560 12165 3624
rect 12182 3560 12246 3624
rect 12263 3560 12327 3624
rect 12344 3560 12408 3624
rect 12425 3560 12489 3624
rect 12506 3560 12570 3624
rect 12587 3560 12651 3624
rect 12668 3560 12732 3624
rect 12749 3560 12813 3624
rect 12830 3560 12894 3624
rect 12911 3560 12975 3624
rect 12992 3560 13056 3624
rect 13073 3560 13137 3624
rect 13154 3560 13218 3624
rect 13235 3560 13299 3624
rect 13316 3560 13380 3624
rect 13397 3560 13461 3624
rect 13478 3560 13542 3624
rect 13559 3560 13623 3624
rect 13640 3560 13704 3624
rect 13721 3560 13785 3624
rect 13802 3560 13866 3624
rect 13883 3560 13947 3624
rect 13964 3560 14028 3624
rect 14045 3560 14109 3624
rect 14126 3560 14190 3624
rect 14207 3560 14271 3624
rect 14288 3560 14352 3624
rect 14369 3560 14433 3624
rect 14451 3560 14515 3624
rect 14533 3560 14597 3624
rect 14615 3560 14679 3624
rect 14697 3560 14761 3624
rect 14779 3560 14843 3624
rect 14861 3560 14925 3624
<< metal4 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 18592 254 18600
rect 14746 18593 15000 18600
rect 0 18591 2821 18592
rect 0 18527 135 18591
rect 199 18527 217 18591
rect 281 18527 299 18591
rect 363 18527 381 18591
rect 445 18527 463 18591
rect 527 18527 545 18591
rect 609 18527 627 18591
rect 691 18527 709 18591
rect 773 18527 791 18591
rect 855 18527 873 18591
rect 937 18527 955 18591
rect 1019 18527 1037 18591
rect 1101 18527 1119 18591
rect 1183 18527 1201 18591
rect 1265 18527 1283 18591
rect 1347 18527 1365 18591
rect 1429 18527 1447 18591
rect 1511 18527 1529 18591
rect 1593 18527 1611 18591
rect 1675 18527 1693 18591
rect 1757 18527 1775 18591
rect 1839 18527 1857 18591
rect 1921 18527 1939 18591
rect 2003 18527 2021 18591
rect 2085 18527 2103 18591
rect 2167 18527 2185 18591
rect 2249 18527 2267 18591
rect 2331 18527 2349 18591
rect 2413 18527 2431 18591
rect 2495 18527 2513 18591
rect 2577 18527 2594 18591
rect 2658 18527 2675 18591
rect 2739 18527 2756 18591
rect 2820 18527 2821 18591
rect 0 18509 2821 18527
rect 0 18445 135 18509
rect 199 18445 217 18509
rect 281 18445 299 18509
rect 363 18445 381 18509
rect 445 18445 463 18509
rect 527 18445 545 18509
rect 609 18445 627 18509
rect 691 18445 709 18509
rect 773 18445 791 18509
rect 855 18445 873 18509
rect 937 18445 955 18509
rect 1019 18445 1037 18509
rect 1101 18445 1119 18509
rect 1183 18445 1201 18509
rect 1265 18445 1283 18509
rect 1347 18445 1365 18509
rect 1429 18445 1447 18509
rect 1511 18445 1529 18509
rect 1593 18445 1611 18509
rect 1675 18445 1693 18509
rect 1757 18445 1775 18509
rect 1839 18445 1857 18509
rect 1921 18445 1939 18509
rect 2003 18445 2021 18509
rect 2085 18445 2103 18509
rect 2167 18445 2185 18509
rect 2249 18445 2267 18509
rect 2331 18445 2349 18509
rect 2413 18445 2431 18509
rect 2495 18445 2513 18509
rect 2577 18445 2594 18509
rect 2658 18445 2675 18509
rect 2739 18445 2756 18509
rect 2820 18445 2821 18509
rect 0 18427 2821 18445
rect 0 18363 135 18427
rect 199 18363 217 18427
rect 281 18363 299 18427
rect 363 18363 381 18427
rect 445 18363 463 18427
rect 527 18363 545 18427
rect 609 18363 627 18427
rect 691 18363 709 18427
rect 773 18363 791 18427
rect 855 18363 873 18427
rect 937 18363 955 18427
rect 1019 18363 1037 18427
rect 1101 18363 1119 18427
rect 1183 18363 1201 18427
rect 1265 18363 1283 18427
rect 1347 18363 1365 18427
rect 1429 18363 1447 18427
rect 1511 18363 1529 18427
rect 1593 18363 1611 18427
rect 1675 18363 1693 18427
rect 1757 18363 1775 18427
rect 1839 18363 1857 18427
rect 1921 18363 1939 18427
rect 2003 18363 2021 18427
rect 2085 18363 2103 18427
rect 2167 18363 2185 18427
rect 2249 18363 2267 18427
rect 2331 18363 2349 18427
rect 2413 18363 2431 18427
rect 2495 18363 2513 18427
rect 2577 18363 2594 18427
rect 2658 18363 2675 18427
rect 2739 18363 2756 18427
rect 2820 18363 2821 18427
rect 0 18345 2821 18363
rect 0 18281 135 18345
rect 199 18281 217 18345
rect 281 18281 299 18345
rect 363 18281 381 18345
rect 445 18281 463 18345
rect 527 18281 545 18345
rect 609 18281 627 18345
rect 691 18281 709 18345
rect 773 18281 791 18345
rect 855 18281 873 18345
rect 937 18281 955 18345
rect 1019 18281 1037 18345
rect 1101 18281 1119 18345
rect 1183 18281 1201 18345
rect 1265 18281 1283 18345
rect 1347 18281 1365 18345
rect 1429 18281 1447 18345
rect 1511 18281 1529 18345
rect 1593 18281 1611 18345
rect 1675 18281 1693 18345
rect 1757 18281 1775 18345
rect 1839 18281 1857 18345
rect 1921 18281 1939 18345
rect 2003 18281 2021 18345
rect 2085 18281 2103 18345
rect 2167 18281 2185 18345
rect 2249 18281 2267 18345
rect 2331 18281 2349 18345
rect 2413 18281 2431 18345
rect 2495 18281 2513 18345
rect 2577 18281 2594 18345
rect 2658 18281 2675 18345
rect 2739 18281 2756 18345
rect 2820 18281 2821 18345
rect 12230 18591 15000 18593
rect 12230 18527 12231 18591
rect 12295 18527 12312 18591
rect 12376 18527 12393 18591
rect 12457 18527 12474 18591
rect 12538 18527 12556 18591
rect 12620 18527 12638 18591
rect 12702 18527 12720 18591
rect 12784 18527 12802 18591
rect 12866 18527 12884 18591
rect 12948 18527 12966 18591
rect 13030 18527 13048 18591
rect 13112 18527 13130 18591
rect 13194 18527 13212 18591
rect 13276 18527 13294 18591
rect 13358 18527 13376 18591
rect 13440 18527 13458 18591
rect 13522 18527 13540 18591
rect 13604 18527 13622 18591
rect 13686 18527 13704 18591
rect 13768 18527 13786 18591
rect 13850 18527 13868 18591
rect 13932 18527 13950 18591
rect 14014 18527 14032 18591
rect 14096 18527 14114 18591
rect 14178 18527 14196 18591
rect 14260 18527 14278 18591
rect 14342 18527 14360 18591
rect 14424 18527 14442 18591
rect 14506 18527 14524 18591
rect 14588 18527 14606 18591
rect 14670 18527 14688 18591
rect 14752 18527 14770 18591
rect 14834 18527 14852 18591
rect 14916 18527 15000 18591
rect 12230 18509 15000 18527
rect 12230 18445 12231 18509
rect 12295 18445 12312 18509
rect 12376 18445 12393 18509
rect 12457 18445 12474 18509
rect 12538 18445 12556 18509
rect 12620 18445 12638 18509
rect 12702 18445 12720 18509
rect 12784 18445 12802 18509
rect 12866 18445 12884 18509
rect 12948 18445 12966 18509
rect 13030 18445 13048 18509
rect 13112 18445 13130 18509
rect 13194 18445 13212 18509
rect 13276 18445 13294 18509
rect 13358 18445 13376 18509
rect 13440 18445 13458 18509
rect 13522 18445 13540 18509
rect 13604 18445 13622 18509
rect 13686 18445 13704 18509
rect 13768 18445 13786 18509
rect 13850 18445 13868 18509
rect 13932 18445 13950 18509
rect 14014 18445 14032 18509
rect 14096 18445 14114 18509
rect 14178 18445 14196 18509
rect 14260 18445 14278 18509
rect 14342 18445 14360 18509
rect 14424 18445 14442 18509
rect 14506 18445 14524 18509
rect 14588 18445 14606 18509
rect 14670 18445 14688 18509
rect 14752 18445 14770 18509
rect 14834 18445 14852 18509
rect 14916 18445 15000 18509
rect 12230 18427 15000 18445
rect 12230 18363 12231 18427
rect 12295 18363 12312 18427
rect 12376 18363 12393 18427
rect 12457 18363 12474 18427
rect 12538 18363 12556 18427
rect 12620 18363 12638 18427
rect 12702 18363 12720 18427
rect 12784 18363 12802 18427
rect 12866 18363 12884 18427
rect 12948 18363 12966 18427
rect 13030 18363 13048 18427
rect 13112 18363 13130 18427
rect 13194 18363 13212 18427
rect 13276 18363 13294 18427
rect 13358 18363 13376 18427
rect 13440 18363 13458 18427
rect 13522 18363 13540 18427
rect 13604 18363 13622 18427
rect 13686 18363 13704 18427
rect 13768 18363 13786 18427
rect 13850 18363 13868 18427
rect 13932 18363 13950 18427
rect 14014 18363 14032 18427
rect 14096 18363 14114 18427
rect 14178 18363 14196 18427
rect 14260 18363 14278 18427
rect 14342 18363 14360 18427
rect 14424 18363 14442 18427
rect 14506 18363 14524 18427
rect 14588 18363 14606 18427
rect 14670 18363 14688 18427
rect 14752 18363 14770 18427
rect 14834 18363 14852 18427
rect 14916 18363 15000 18427
rect 12230 18345 15000 18363
rect 0 18263 2821 18281
rect 0 18199 135 18263
rect 199 18199 217 18263
rect 281 18199 299 18263
rect 363 18199 381 18263
rect 445 18199 463 18263
rect 527 18199 545 18263
rect 609 18199 627 18263
rect 691 18199 709 18263
rect 773 18199 791 18263
rect 855 18199 873 18263
rect 937 18199 955 18263
rect 1019 18199 1037 18263
rect 1101 18199 1119 18263
rect 1183 18199 1201 18263
rect 1265 18199 1283 18263
rect 1347 18199 1365 18263
rect 1429 18199 1447 18263
rect 1511 18199 1529 18263
rect 1593 18199 1611 18263
rect 1675 18199 1693 18263
rect 1757 18199 1775 18263
rect 1839 18199 1857 18263
rect 1921 18199 1939 18263
rect 2003 18199 2021 18263
rect 2085 18199 2103 18263
rect 2167 18199 2185 18263
rect 2249 18199 2267 18263
rect 2331 18199 2349 18263
rect 2413 18199 2431 18263
rect 2495 18199 2513 18263
rect 2577 18199 2594 18263
rect 2658 18199 2675 18263
rect 2739 18199 2756 18263
rect 2820 18199 2821 18263
rect 0 18181 2821 18199
rect 2851 18341 3073 18342
rect 2851 18277 2852 18341
rect 2916 18277 3008 18341
rect 3072 18277 3073 18341
rect 2851 18255 3073 18277
rect 2851 18191 2852 18255
rect 2916 18191 3008 18255
rect 3072 18191 3073 18255
rect 2851 18190 3073 18191
rect 11978 18341 12200 18342
rect 11978 18277 11979 18341
rect 12043 18277 12135 18341
rect 12199 18277 12200 18341
rect 11978 18255 12200 18277
rect 11978 18191 11979 18255
rect 12043 18191 12135 18255
rect 12199 18191 12200 18255
rect 11978 18190 12200 18191
rect 12230 18281 12231 18345
rect 12295 18281 12312 18345
rect 12376 18281 12393 18345
rect 12457 18281 12474 18345
rect 12538 18281 12556 18345
rect 12620 18281 12638 18345
rect 12702 18281 12720 18345
rect 12784 18281 12802 18345
rect 12866 18281 12884 18345
rect 12948 18281 12966 18345
rect 13030 18281 13048 18345
rect 13112 18281 13130 18345
rect 13194 18281 13212 18345
rect 13276 18281 13294 18345
rect 13358 18281 13376 18345
rect 13440 18281 13458 18345
rect 13522 18281 13540 18345
rect 13604 18281 13622 18345
rect 13686 18281 13704 18345
rect 13768 18281 13786 18345
rect 13850 18281 13868 18345
rect 13932 18281 13950 18345
rect 14014 18281 14032 18345
rect 14096 18281 14114 18345
rect 14178 18281 14196 18345
rect 14260 18281 14278 18345
rect 14342 18281 14360 18345
rect 14424 18281 14442 18345
rect 14506 18281 14524 18345
rect 14588 18281 14606 18345
rect 14670 18281 14688 18345
rect 14752 18281 14770 18345
rect 14834 18281 14852 18345
rect 14916 18281 15000 18345
rect 12230 18263 15000 18281
rect 12230 18199 12231 18263
rect 12295 18199 12312 18263
rect 12376 18199 12393 18263
rect 12457 18199 12474 18263
rect 12538 18199 12556 18263
rect 12620 18199 12638 18263
rect 12702 18199 12720 18263
rect 12784 18199 12802 18263
rect 12866 18199 12884 18263
rect 12948 18199 12966 18263
rect 13030 18199 13048 18263
rect 13112 18199 13130 18263
rect 13194 18199 13212 18263
rect 13276 18199 13294 18263
rect 13358 18199 13376 18263
rect 13440 18199 13458 18263
rect 13522 18199 13540 18263
rect 13604 18199 13622 18263
rect 13686 18199 13704 18263
rect 13768 18199 13786 18263
rect 13850 18199 13868 18263
rect 13932 18199 13950 18263
rect 14014 18199 14032 18263
rect 14096 18199 14114 18263
rect 14178 18199 14196 18263
rect 14260 18199 14278 18263
rect 14342 18199 14360 18263
rect 14424 18199 14442 18263
rect 14506 18199 14524 18263
rect 14588 18199 14606 18263
rect 14670 18199 14688 18263
rect 14752 18199 14770 18263
rect 14834 18199 14852 18263
rect 14916 18199 15000 18263
rect 0 18117 135 18181
rect 199 18117 217 18181
rect 281 18117 299 18181
rect 363 18117 381 18181
rect 445 18117 463 18181
rect 527 18117 545 18181
rect 609 18117 627 18181
rect 691 18117 709 18181
rect 773 18117 791 18181
rect 855 18117 873 18181
rect 937 18117 955 18181
rect 1019 18117 1037 18181
rect 1101 18117 1119 18181
rect 1183 18117 1201 18181
rect 1265 18117 1283 18181
rect 1347 18117 1365 18181
rect 1429 18117 1447 18181
rect 1511 18117 1529 18181
rect 1593 18117 1611 18181
rect 1675 18117 1693 18181
rect 1757 18117 1775 18181
rect 1839 18117 1857 18181
rect 1921 18117 1939 18181
rect 2003 18117 2021 18181
rect 2085 18117 2103 18181
rect 2167 18117 2185 18181
rect 2249 18117 2267 18181
rect 2331 18117 2349 18181
rect 2413 18117 2431 18181
rect 2495 18117 2513 18181
rect 2577 18117 2594 18181
rect 2658 18117 2675 18181
rect 2739 18117 2756 18181
rect 2820 18117 2821 18181
rect 12230 18181 15000 18199
rect 0 18099 2821 18117
rect 0 18035 135 18099
rect 199 18035 217 18099
rect 281 18035 299 18099
rect 363 18035 381 18099
rect 445 18035 463 18099
rect 527 18035 545 18099
rect 609 18035 627 18099
rect 691 18035 709 18099
rect 773 18035 791 18099
rect 855 18035 873 18099
rect 937 18035 955 18099
rect 1019 18035 1037 18099
rect 1101 18035 1119 18099
rect 1183 18035 1201 18099
rect 1265 18035 1283 18099
rect 1347 18035 1365 18099
rect 1429 18035 1447 18099
rect 1511 18035 1529 18099
rect 1593 18035 1611 18099
rect 1675 18035 1693 18099
rect 1757 18035 1775 18099
rect 1839 18035 1857 18099
rect 1921 18035 1939 18099
rect 2003 18035 2021 18099
rect 2085 18035 2103 18099
rect 2167 18035 2185 18099
rect 2249 18035 2267 18099
rect 2331 18035 2349 18099
rect 2413 18035 2431 18099
rect 2495 18035 2513 18099
rect 2577 18035 2594 18099
rect 2658 18035 2675 18099
rect 2739 18035 2756 18099
rect 2820 18035 2821 18099
rect 0 18017 2821 18035
rect 0 17953 135 18017
rect 199 17953 217 18017
rect 281 17953 299 18017
rect 363 17953 381 18017
rect 445 17953 463 18017
rect 527 17953 545 18017
rect 609 17953 627 18017
rect 691 17953 709 18017
rect 773 17953 791 18017
rect 855 17953 873 18017
rect 937 17953 955 18017
rect 1019 17953 1037 18017
rect 1101 17953 1119 18017
rect 1183 17953 1201 18017
rect 1265 17953 1283 18017
rect 1347 17953 1365 18017
rect 1429 17953 1447 18017
rect 1511 17953 1529 18017
rect 1593 17953 1611 18017
rect 1675 17953 1693 18017
rect 1757 17953 1775 18017
rect 1839 17953 1857 18017
rect 1921 17953 1939 18017
rect 2003 17953 2021 18017
rect 2085 17953 2103 18017
rect 2167 17953 2185 18017
rect 2249 17953 2267 18017
rect 2331 17953 2349 18017
rect 2413 17953 2431 18017
rect 2495 17953 2513 18017
rect 2577 17953 2594 18017
rect 2658 17953 2675 18017
rect 2739 17953 2756 18017
rect 2820 17953 2821 18017
rect 0 17935 2821 17953
rect 0 17871 135 17935
rect 199 17871 217 17935
rect 281 17871 299 17935
rect 363 17871 381 17935
rect 445 17871 463 17935
rect 527 17871 545 17935
rect 609 17871 627 17935
rect 691 17871 709 17935
rect 773 17871 791 17935
rect 855 17871 873 17935
rect 937 17871 955 17935
rect 1019 17871 1037 17935
rect 1101 17871 1119 17935
rect 1183 17871 1201 17935
rect 1265 17871 1283 17935
rect 1347 17871 1365 17935
rect 1429 17871 1447 17935
rect 1511 17871 1529 17935
rect 1593 17871 1611 17935
rect 1675 17871 1693 17935
rect 1757 17871 1775 17935
rect 1839 17871 1857 17935
rect 1921 17871 1939 17935
rect 2003 17871 2021 17935
rect 2085 17871 2103 17935
rect 2167 17871 2185 17935
rect 2249 17871 2267 17935
rect 2331 17871 2349 17935
rect 2413 17871 2431 17935
rect 2495 17871 2513 17935
rect 2577 17871 2594 17935
rect 2658 17871 2675 17935
rect 2739 17871 2756 17935
rect 2820 17871 2821 17935
rect 0 17853 2821 17871
rect 0 17789 135 17853
rect 199 17789 217 17853
rect 281 17789 299 17853
rect 363 17789 381 17853
rect 445 17789 463 17853
rect 527 17789 545 17853
rect 609 17789 627 17853
rect 691 17789 709 17853
rect 773 17789 791 17853
rect 855 17789 873 17853
rect 937 17789 955 17853
rect 1019 17789 1037 17853
rect 1101 17789 1119 17853
rect 1183 17789 1201 17853
rect 1265 17789 1283 17853
rect 1347 17789 1365 17853
rect 1429 17789 1447 17853
rect 1511 17789 1529 17853
rect 1593 17789 1611 17853
rect 1675 17789 1693 17853
rect 1757 17789 1775 17853
rect 1839 17789 1857 17853
rect 1921 17789 1939 17853
rect 2003 17789 2021 17853
rect 2085 17789 2103 17853
rect 2167 17789 2185 17853
rect 2249 17789 2267 17853
rect 2331 17789 2349 17853
rect 2413 17789 2431 17853
rect 2495 17789 2513 17853
rect 2577 17789 2594 17853
rect 2658 17789 2675 17853
rect 2739 17789 2756 17853
rect 2820 17789 2821 17853
rect 0 17771 2821 17789
rect 0 17707 135 17771
rect 199 17707 217 17771
rect 281 17707 299 17771
rect 363 17707 381 17771
rect 445 17707 463 17771
rect 527 17707 545 17771
rect 609 17707 627 17771
rect 691 17707 709 17771
rect 773 17707 791 17771
rect 855 17707 873 17771
rect 937 17707 955 17771
rect 1019 17707 1037 17771
rect 1101 17707 1119 17771
rect 1183 17707 1201 17771
rect 1265 17707 1283 17771
rect 1347 17707 1365 17771
rect 1429 17707 1447 17771
rect 1511 17707 1529 17771
rect 1593 17707 1611 17771
rect 1675 17707 1693 17771
rect 1757 17707 1775 17771
rect 1839 17707 1857 17771
rect 1921 17707 1939 17771
rect 2003 17707 2021 17771
rect 2085 17707 2103 17771
rect 2167 17707 2185 17771
rect 2249 17707 2267 17771
rect 2331 17707 2349 17771
rect 2413 17707 2431 17771
rect 2495 17707 2513 17771
rect 2577 17707 2594 17771
rect 2658 17707 2675 17771
rect 2739 17707 2756 17771
rect 2820 17707 2821 17771
rect 0 17689 2821 17707
rect 0 17625 135 17689
rect 199 17625 217 17689
rect 281 17625 299 17689
rect 363 17625 381 17689
rect 445 17625 463 17689
rect 527 17625 545 17689
rect 609 17625 627 17689
rect 691 17625 709 17689
rect 773 17625 791 17689
rect 855 17625 873 17689
rect 937 17625 955 17689
rect 1019 17625 1037 17689
rect 1101 17625 1119 17689
rect 1183 17625 1201 17689
rect 1265 17625 1283 17689
rect 1347 17625 1365 17689
rect 1429 17625 1447 17689
rect 1511 17625 1529 17689
rect 1593 17625 1611 17689
rect 1675 17625 1693 17689
rect 1757 17625 1775 17689
rect 1839 17625 1857 17689
rect 1921 17625 1939 17689
rect 2003 17625 2021 17689
rect 2085 17625 2103 17689
rect 2167 17625 2185 17689
rect 2249 17625 2267 17689
rect 2331 17625 2349 17689
rect 2413 17625 2431 17689
rect 2495 17625 2513 17689
rect 2577 17625 2594 17689
rect 2658 17625 2675 17689
rect 2739 17625 2756 17689
rect 2820 17625 2821 17689
rect 2854 18163 3250 18164
rect 2854 18099 2856 18163
rect 2920 18099 2938 18163
rect 3002 18099 3020 18163
rect 3084 18099 3102 18163
rect 3166 18099 3184 18163
rect 3248 18099 3250 18163
rect 2854 18077 3250 18099
rect 2854 18013 2856 18077
rect 2920 18013 2938 18077
rect 3002 18013 3020 18077
rect 3084 18013 3102 18077
rect 3166 18013 3184 18077
rect 3248 18013 3250 18077
rect 2854 17991 3250 18013
rect 2854 17927 2856 17991
rect 2920 17927 2938 17991
rect 3002 17927 3020 17991
rect 3084 17927 3102 17991
rect 3166 17927 3184 17991
rect 3248 17927 3250 17991
rect 2854 17905 3250 17927
rect 11801 18163 12197 18164
rect 11801 18099 11803 18163
rect 11867 18099 11885 18163
rect 11949 18099 11967 18163
rect 12031 18099 12049 18163
rect 12113 18099 12131 18163
rect 12195 18099 12197 18163
rect 11801 18077 12197 18099
rect 11801 18013 11803 18077
rect 11867 18013 11885 18077
rect 11949 18013 11967 18077
rect 12031 18013 12049 18077
rect 12113 18013 12131 18077
rect 12195 18013 12197 18077
rect 11801 17991 12197 18013
rect 11801 17927 11803 17991
rect 11867 17927 11885 17991
rect 11949 17927 11967 17991
rect 12031 17927 12049 17991
rect 12113 17927 12131 17991
rect 12195 17927 12197 17991
rect 2854 17841 2856 17905
rect 2920 17841 2938 17905
rect 3002 17841 3020 17905
rect 3084 17841 3102 17905
rect 3166 17841 3184 17905
rect 3248 17841 3250 17905
rect 2854 17819 3250 17841
rect 2854 17755 2856 17819
rect 2920 17755 2938 17819
rect 3002 17755 3020 17819
rect 3084 17755 3102 17819
rect 3166 17755 3184 17819
rect 3248 17755 3250 17819
rect 2854 17734 3250 17755
rect 2854 17670 2856 17734
rect 2920 17670 2938 17734
rect 3002 17670 3020 17734
rect 3084 17670 3102 17734
rect 3166 17670 3184 17734
rect 3248 17670 3250 17734
rect 3283 17905 3505 17906
rect 3283 17841 3284 17905
rect 3348 17841 3440 17905
rect 3504 17841 3505 17905
rect 3283 17821 3505 17841
rect 3283 17757 3284 17821
rect 3348 17757 3440 17821
rect 3504 17757 3505 17821
rect 3283 17738 3505 17757
rect 3283 17674 3284 17738
rect 3348 17674 3440 17738
rect 3504 17674 3505 17738
rect 3283 17673 3505 17674
rect 11546 17905 11768 17906
rect 11546 17841 11547 17905
rect 11611 17841 11703 17905
rect 11767 17841 11768 17905
rect 11546 17821 11768 17841
rect 11546 17757 11547 17821
rect 11611 17757 11703 17821
rect 11767 17757 11768 17821
rect 11546 17738 11768 17757
rect 11546 17674 11547 17738
rect 11611 17674 11703 17738
rect 11767 17674 11768 17738
rect 11546 17673 11768 17674
rect 11801 17905 12197 17927
rect 11801 17841 11803 17905
rect 11867 17841 11885 17905
rect 11949 17841 11967 17905
rect 12031 17841 12049 17905
rect 12113 17841 12131 17905
rect 12195 17841 12197 17905
rect 11801 17819 12197 17841
rect 11801 17755 11803 17819
rect 11867 17755 11885 17819
rect 11949 17755 11967 17819
rect 12031 17755 12049 17819
rect 12113 17755 12131 17819
rect 12195 17755 12197 17819
rect 11801 17734 12197 17755
rect 2854 17669 3250 17670
rect 11801 17670 11803 17734
rect 11867 17670 11885 17734
rect 11949 17670 11967 17734
rect 12031 17670 12049 17734
rect 12113 17670 12131 17734
rect 12195 17670 12197 17734
rect 11801 17669 12197 17670
rect 12230 18117 12231 18181
rect 12295 18117 12312 18181
rect 12376 18117 12393 18181
rect 12457 18117 12474 18181
rect 12538 18117 12556 18181
rect 12620 18117 12638 18181
rect 12702 18117 12720 18181
rect 12784 18117 12802 18181
rect 12866 18117 12884 18181
rect 12948 18117 12966 18181
rect 13030 18117 13048 18181
rect 13112 18117 13130 18181
rect 13194 18117 13212 18181
rect 13276 18117 13294 18181
rect 13358 18117 13376 18181
rect 13440 18117 13458 18181
rect 13522 18117 13540 18181
rect 13604 18117 13622 18181
rect 13686 18117 13704 18181
rect 13768 18117 13786 18181
rect 13850 18117 13868 18181
rect 13932 18117 13950 18181
rect 14014 18117 14032 18181
rect 14096 18117 14114 18181
rect 14178 18117 14196 18181
rect 14260 18117 14278 18181
rect 14342 18117 14360 18181
rect 14424 18117 14442 18181
rect 14506 18117 14524 18181
rect 14588 18117 14606 18181
rect 14670 18117 14688 18181
rect 14752 18117 14770 18181
rect 14834 18117 14852 18181
rect 14916 18117 15000 18181
rect 12230 18099 15000 18117
rect 12230 18035 12231 18099
rect 12295 18035 12312 18099
rect 12376 18035 12393 18099
rect 12457 18035 12474 18099
rect 12538 18035 12556 18099
rect 12620 18035 12638 18099
rect 12702 18035 12720 18099
rect 12784 18035 12802 18099
rect 12866 18035 12884 18099
rect 12948 18035 12966 18099
rect 13030 18035 13048 18099
rect 13112 18035 13130 18099
rect 13194 18035 13212 18099
rect 13276 18035 13294 18099
rect 13358 18035 13376 18099
rect 13440 18035 13458 18099
rect 13522 18035 13540 18099
rect 13604 18035 13622 18099
rect 13686 18035 13704 18099
rect 13768 18035 13786 18099
rect 13850 18035 13868 18099
rect 13932 18035 13950 18099
rect 14014 18035 14032 18099
rect 14096 18035 14114 18099
rect 14178 18035 14196 18099
rect 14260 18035 14278 18099
rect 14342 18035 14360 18099
rect 14424 18035 14442 18099
rect 14506 18035 14524 18099
rect 14588 18035 14606 18099
rect 14670 18035 14688 18099
rect 14752 18035 14770 18099
rect 14834 18035 14852 18099
rect 14916 18035 15000 18099
rect 12230 18017 15000 18035
rect 12230 17953 12231 18017
rect 12295 17953 12312 18017
rect 12376 17953 12393 18017
rect 12457 17953 12474 18017
rect 12538 17953 12556 18017
rect 12620 17953 12638 18017
rect 12702 17953 12720 18017
rect 12784 17953 12802 18017
rect 12866 17953 12884 18017
rect 12948 17953 12966 18017
rect 13030 17953 13048 18017
rect 13112 17953 13130 18017
rect 13194 17953 13212 18017
rect 13276 17953 13294 18017
rect 13358 17953 13376 18017
rect 13440 17953 13458 18017
rect 13522 17953 13540 18017
rect 13604 17953 13622 18017
rect 13686 17953 13704 18017
rect 13768 17953 13786 18017
rect 13850 17953 13868 18017
rect 13932 17953 13950 18017
rect 14014 17953 14032 18017
rect 14096 17953 14114 18017
rect 14178 17953 14196 18017
rect 14260 17953 14278 18017
rect 14342 17953 14360 18017
rect 14424 17953 14442 18017
rect 14506 17953 14524 18017
rect 14588 17953 14606 18017
rect 14670 17953 14688 18017
rect 14752 17953 14770 18017
rect 14834 17953 14852 18017
rect 14916 17953 15000 18017
rect 12230 17935 15000 17953
rect 12230 17871 12231 17935
rect 12295 17871 12312 17935
rect 12376 17871 12393 17935
rect 12457 17871 12474 17935
rect 12538 17871 12556 17935
rect 12620 17871 12638 17935
rect 12702 17871 12720 17935
rect 12784 17871 12802 17935
rect 12866 17871 12884 17935
rect 12948 17871 12966 17935
rect 13030 17871 13048 17935
rect 13112 17871 13130 17935
rect 13194 17871 13212 17935
rect 13276 17871 13294 17935
rect 13358 17871 13376 17935
rect 13440 17871 13458 17935
rect 13522 17871 13540 17935
rect 13604 17871 13622 17935
rect 13686 17871 13704 17935
rect 13768 17871 13786 17935
rect 13850 17871 13868 17935
rect 13932 17871 13950 17935
rect 14014 17871 14032 17935
rect 14096 17871 14114 17935
rect 14178 17871 14196 17935
rect 14260 17871 14278 17935
rect 14342 17871 14360 17935
rect 14424 17871 14442 17935
rect 14506 17871 14524 17935
rect 14588 17871 14606 17935
rect 14670 17871 14688 17935
rect 14752 17871 14770 17935
rect 14834 17871 14852 17935
rect 14916 17871 15000 17935
rect 12230 17853 15000 17871
rect 12230 17789 12231 17853
rect 12295 17789 12312 17853
rect 12376 17789 12393 17853
rect 12457 17789 12474 17853
rect 12538 17789 12556 17853
rect 12620 17789 12638 17853
rect 12702 17789 12720 17853
rect 12784 17789 12802 17853
rect 12866 17789 12884 17853
rect 12948 17789 12966 17853
rect 13030 17789 13048 17853
rect 13112 17789 13130 17853
rect 13194 17789 13212 17853
rect 13276 17789 13294 17853
rect 13358 17789 13376 17853
rect 13440 17789 13458 17853
rect 13522 17789 13540 17853
rect 13604 17789 13622 17853
rect 13686 17789 13704 17853
rect 13768 17789 13786 17853
rect 13850 17789 13868 17853
rect 13932 17789 13950 17853
rect 14014 17789 14032 17853
rect 14096 17789 14114 17853
rect 14178 17789 14196 17853
rect 14260 17789 14278 17853
rect 14342 17789 14360 17853
rect 14424 17789 14442 17853
rect 14506 17789 14524 17853
rect 14588 17789 14606 17853
rect 14670 17789 14688 17853
rect 14752 17789 14770 17853
rect 14834 17789 14852 17853
rect 14916 17789 15000 17853
rect 12230 17771 15000 17789
rect 12230 17707 12231 17771
rect 12295 17707 12312 17771
rect 12376 17707 12393 17771
rect 12457 17707 12474 17771
rect 12538 17707 12556 17771
rect 12620 17707 12638 17771
rect 12702 17707 12720 17771
rect 12784 17707 12802 17771
rect 12866 17707 12884 17771
rect 12948 17707 12966 17771
rect 13030 17707 13048 17771
rect 13112 17707 13130 17771
rect 13194 17707 13212 17771
rect 13276 17707 13294 17771
rect 13358 17707 13376 17771
rect 13440 17707 13458 17771
rect 13522 17707 13540 17771
rect 13604 17707 13622 17771
rect 13686 17707 13704 17771
rect 13768 17707 13786 17771
rect 13850 17707 13868 17771
rect 13932 17707 13950 17771
rect 14014 17707 14032 17771
rect 14096 17707 14114 17771
rect 14178 17707 14196 17771
rect 14260 17707 14278 17771
rect 14342 17707 14360 17771
rect 14424 17707 14442 17771
rect 14506 17707 14524 17771
rect 14588 17707 14606 17771
rect 14670 17707 14688 17771
rect 14752 17707 14770 17771
rect 14834 17707 14852 17771
rect 14916 17707 15000 17771
rect 12230 17689 15000 17707
rect 0 17607 2821 17625
rect 0 17543 135 17607
rect 199 17543 217 17607
rect 281 17543 299 17607
rect 363 17543 381 17607
rect 445 17543 463 17607
rect 527 17543 545 17607
rect 609 17543 627 17607
rect 691 17543 709 17607
rect 773 17543 791 17607
rect 855 17543 873 17607
rect 937 17543 955 17607
rect 1019 17543 1037 17607
rect 1101 17543 1119 17607
rect 1183 17543 1201 17607
rect 1265 17543 1283 17607
rect 1347 17543 1365 17607
rect 1429 17543 1447 17607
rect 1511 17543 1529 17607
rect 1593 17543 1611 17607
rect 1675 17543 1693 17607
rect 1757 17543 1775 17607
rect 1839 17543 1857 17607
rect 1921 17543 1939 17607
rect 2003 17543 2021 17607
rect 2085 17543 2103 17607
rect 2167 17543 2185 17607
rect 2249 17543 2267 17607
rect 2331 17543 2349 17607
rect 2413 17543 2431 17607
rect 2495 17543 2513 17607
rect 2577 17543 2594 17607
rect 2658 17543 2675 17607
rect 2739 17543 2756 17607
rect 2820 17543 2821 17607
rect 0 17525 2821 17543
rect 0 17461 135 17525
rect 199 17461 217 17525
rect 281 17461 299 17525
rect 363 17461 381 17525
rect 445 17461 463 17525
rect 527 17461 545 17525
rect 609 17461 627 17525
rect 691 17461 709 17525
rect 773 17461 791 17525
rect 855 17461 873 17525
rect 937 17461 955 17525
rect 1019 17461 1037 17525
rect 1101 17461 1119 17525
rect 1183 17461 1201 17525
rect 1265 17461 1283 17525
rect 1347 17461 1365 17525
rect 1429 17461 1447 17525
rect 1511 17461 1529 17525
rect 1593 17461 1611 17525
rect 1675 17461 1693 17525
rect 1757 17461 1775 17525
rect 1839 17461 1857 17525
rect 1921 17461 1939 17525
rect 2003 17461 2021 17525
rect 2085 17461 2103 17525
rect 2167 17461 2185 17525
rect 2249 17461 2267 17525
rect 2331 17461 2349 17525
rect 2413 17461 2431 17525
rect 2495 17461 2513 17525
rect 2577 17461 2594 17525
rect 2658 17461 2675 17525
rect 2739 17461 2756 17525
rect 2820 17461 2821 17525
rect 0 17443 2821 17461
rect 0 17379 135 17443
rect 199 17379 217 17443
rect 281 17379 299 17443
rect 363 17379 381 17443
rect 445 17379 463 17443
rect 527 17379 545 17443
rect 609 17379 627 17443
rect 691 17379 709 17443
rect 773 17379 791 17443
rect 855 17379 873 17443
rect 937 17379 955 17443
rect 1019 17379 1037 17443
rect 1101 17379 1119 17443
rect 1183 17379 1201 17443
rect 1265 17379 1283 17443
rect 1347 17379 1365 17443
rect 1429 17379 1447 17443
rect 1511 17379 1529 17443
rect 1593 17379 1611 17443
rect 1675 17379 1693 17443
rect 1757 17379 1775 17443
rect 1839 17379 1857 17443
rect 1921 17379 1939 17443
rect 2003 17379 2021 17443
rect 2085 17379 2103 17443
rect 2167 17379 2185 17443
rect 2249 17379 2267 17443
rect 2331 17379 2349 17443
rect 2413 17379 2431 17443
rect 2495 17379 2513 17443
rect 2577 17379 2594 17443
rect 2658 17379 2675 17443
rect 2739 17379 2756 17443
rect 2820 17379 2821 17443
rect 0 17361 2821 17379
rect 0 17297 135 17361
rect 199 17297 217 17361
rect 281 17297 299 17361
rect 363 17297 381 17361
rect 445 17297 463 17361
rect 527 17297 545 17361
rect 609 17297 627 17361
rect 691 17297 709 17361
rect 773 17297 791 17361
rect 855 17297 873 17361
rect 937 17297 955 17361
rect 1019 17297 1037 17361
rect 1101 17297 1119 17361
rect 1183 17297 1201 17361
rect 1265 17297 1283 17361
rect 1347 17297 1365 17361
rect 1429 17297 1447 17361
rect 1511 17297 1529 17361
rect 1593 17297 1611 17361
rect 1675 17297 1693 17361
rect 1757 17297 1775 17361
rect 1839 17297 1857 17361
rect 1921 17297 1939 17361
rect 2003 17297 2021 17361
rect 2085 17297 2103 17361
rect 2167 17297 2185 17361
rect 2249 17297 2267 17361
rect 2331 17297 2349 17361
rect 2413 17297 2431 17361
rect 2495 17297 2513 17361
rect 2577 17297 2594 17361
rect 2658 17297 2675 17361
rect 2739 17297 2756 17361
rect 2820 17297 2821 17361
rect 0 17279 2821 17297
rect 0 17215 135 17279
rect 199 17215 217 17279
rect 281 17215 299 17279
rect 363 17215 381 17279
rect 445 17215 463 17279
rect 527 17215 545 17279
rect 609 17215 627 17279
rect 691 17215 709 17279
rect 773 17215 791 17279
rect 855 17215 873 17279
rect 937 17215 955 17279
rect 1019 17215 1037 17279
rect 1101 17215 1119 17279
rect 1183 17215 1201 17279
rect 1265 17215 1283 17279
rect 1347 17215 1365 17279
rect 1429 17215 1447 17279
rect 1511 17215 1529 17279
rect 1593 17215 1611 17279
rect 1675 17215 1693 17279
rect 1757 17215 1775 17279
rect 1839 17215 1857 17279
rect 1921 17215 1939 17279
rect 2003 17215 2021 17279
rect 2085 17215 2103 17279
rect 2167 17215 2185 17279
rect 2249 17215 2267 17279
rect 2331 17215 2349 17279
rect 2413 17215 2431 17279
rect 2495 17215 2513 17279
rect 2577 17215 2594 17279
rect 2658 17215 2675 17279
rect 2739 17215 2756 17279
rect 2820 17215 2821 17279
rect 0 17197 2821 17215
rect 0 17133 135 17197
rect 199 17133 217 17197
rect 281 17133 299 17197
rect 363 17133 381 17197
rect 445 17133 463 17197
rect 527 17133 545 17197
rect 609 17133 627 17197
rect 691 17133 709 17197
rect 773 17133 791 17197
rect 855 17133 873 17197
rect 937 17133 955 17197
rect 1019 17133 1037 17197
rect 1101 17133 1119 17197
rect 1183 17133 1201 17197
rect 1265 17133 1283 17197
rect 1347 17133 1365 17197
rect 1429 17133 1447 17197
rect 1511 17133 1529 17197
rect 1593 17133 1611 17197
rect 1675 17133 1693 17197
rect 1757 17133 1775 17197
rect 1839 17133 1857 17197
rect 1921 17133 1939 17197
rect 2003 17133 2021 17197
rect 2085 17133 2103 17197
rect 2167 17133 2185 17197
rect 2249 17133 2267 17197
rect 2331 17133 2349 17197
rect 2413 17133 2431 17197
rect 2495 17133 2513 17197
rect 2577 17133 2594 17197
rect 2658 17133 2675 17197
rect 2739 17133 2756 17197
rect 2820 17133 2821 17197
rect 0 17115 2821 17133
rect 0 17051 135 17115
rect 199 17051 217 17115
rect 281 17051 299 17115
rect 363 17051 381 17115
rect 445 17051 463 17115
rect 527 17051 545 17115
rect 609 17051 627 17115
rect 691 17051 709 17115
rect 773 17051 791 17115
rect 855 17051 873 17115
rect 937 17051 955 17115
rect 1019 17051 1037 17115
rect 1101 17051 1119 17115
rect 1183 17051 1201 17115
rect 1265 17051 1283 17115
rect 1347 17051 1365 17115
rect 1429 17051 1447 17115
rect 1511 17051 1529 17115
rect 1593 17051 1611 17115
rect 1675 17051 1693 17115
rect 1757 17051 1775 17115
rect 1839 17051 1857 17115
rect 1921 17051 1939 17115
rect 2003 17051 2021 17115
rect 2085 17051 2103 17115
rect 2167 17051 2185 17115
rect 2249 17051 2267 17115
rect 2331 17051 2349 17115
rect 2413 17051 2431 17115
rect 2495 17051 2513 17115
rect 2577 17051 2594 17115
rect 2658 17051 2675 17115
rect 2739 17051 2756 17115
rect 2820 17051 2821 17115
rect 0 17033 2821 17051
rect 0 16969 135 17033
rect 199 16969 217 17033
rect 281 16969 299 17033
rect 363 16969 381 17033
rect 445 16969 463 17033
rect 527 16969 545 17033
rect 609 16969 627 17033
rect 691 16969 709 17033
rect 773 16969 791 17033
rect 855 16969 873 17033
rect 937 16969 955 17033
rect 1019 16969 1037 17033
rect 1101 16969 1119 17033
rect 1183 16969 1201 17033
rect 1265 16969 1283 17033
rect 1347 16969 1365 17033
rect 1429 16969 1447 17033
rect 1511 16969 1529 17033
rect 1593 16969 1611 17033
rect 1675 16969 1693 17033
rect 1757 16969 1775 17033
rect 1839 16969 1857 17033
rect 1921 16969 1939 17033
rect 2003 16969 2021 17033
rect 2085 16969 2103 17033
rect 2167 16969 2185 17033
rect 2249 16969 2267 17033
rect 2331 16969 2349 17033
rect 2413 16969 2431 17033
rect 2495 16969 2513 17033
rect 2577 16969 2594 17033
rect 2658 16969 2675 17033
rect 2739 16969 2756 17033
rect 2820 16969 2821 17033
rect 0 16951 2821 16969
rect 0 16887 135 16951
rect 199 16887 217 16951
rect 281 16887 299 16951
rect 363 16887 381 16951
rect 445 16887 463 16951
rect 527 16887 545 16951
rect 609 16887 627 16951
rect 691 16887 709 16951
rect 773 16887 791 16951
rect 855 16887 873 16951
rect 937 16887 955 16951
rect 1019 16887 1037 16951
rect 1101 16887 1119 16951
rect 1183 16887 1201 16951
rect 1265 16887 1283 16951
rect 1347 16887 1365 16951
rect 1429 16887 1447 16951
rect 1511 16887 1529 16951
rect 1593 16887 1611 16951
rect 1675 16887 1693 16951
rect 1757 16887 1775 16951
rect 1839 16887 1857 16951
rect 1921 16887 1939 16951
rect 2003 16887 2021 16951
rect 2085 16887 2103 16951
rect 2167 16887 2185 16951
rect 2249 16887 2267 16951
rect 2331 16887 2349 16951
rect 2413 16887 2431 16951
rect 2495 16887 2513 16951
rect 2577 16887 2594 16951
rect 2658 16887 2675 16951
rect 2739 16887 2756 16951
rect 2820 16887 2821 16951
rect 0 16869 2821 16887
rect 0 16805 135 16869
rect 199 16805 217 16869
rect 281 16805 299 16869
rect 363 16805 381 16869
rect 445 16805 463 16869
rect 527 16805 545 16869
rect 609 16805 627 16869
rect 691 16805 709 16869
rect 773 16805 791 16869
rect 855 16805 873 16869
rect 937 16805 955 16869
rect 1019 16805 1037 16869
rect 1101 16805 1119 16869
rect 1183 16805 1201 16869
rect 1265 16805 1283 16869
rect 1347 16805 1365 16869
rect 1429 16805 1447 16869
rect 1511 16805 1529 16869
rect 1593 16805 1611 16869
rect 1675 16805 1693 16869
rect 1757 16805 1775 16869
rect 1839 16805 1857 16869
rect 1921 16805 1939 16869
rect 2003 16805 2021 16869
rect 2085 16805 2103 16869
rect 2167 16805 2185 16869
rect 2249 16805 2267 16869
rect 2331 16805 2349 16869
rect 2413 16805 2431 16869
rect 2495 16805 2513 16869
rect 2577 16805 2594 16869
rect 2658 16805 2675 16869
rect 2739 16805 2756 16869
rect 2820 16805 2821 16869
rect 0 16787 2821 16805
rect 0 16723 135 16787
rect 199 16723 217 16787
rect 281 16723 299 16787
rect 363 16723 381 16787
rect 445 16723 463 16787
rect 527 16723 545 16787
rect 609 16723 627 16787
rect 691 16723 709 16787
rect 773 16723 791 16787
rect 855 16723 873 16787
rect 937 16723 955 16787
rect 1019 16723 1037 16787
rect 1101 16723 1119 16787
rect 1183 16723 1201 16787
rect 1265 16723 1283 16787
rect 1347 16723 1365 16787
rect 1429 16723 1447 16787
rect 1511 16723 1529 16787
rect 1593 16723 1611 16787
rect 1675 16723 1693 16787
rect 1757 16723 1775 16787
rect 1839 16723 1857 16787
rect 1921 16723 1939 16787
rect 2003 16723 2021 16787
rect 2085 16723 2103 16787
rect 2167 16723 2185 16787
rect 2249 16723 2267 16787
rect 2331 16723 2349 16787
rect 2413 16723 2431 16787
rect 2495 16723 2513 16787
rect 2577 16723 2594 16787
rect 2658 16723 2675 16787
rect 2739 16723 2756 16787
rect 2820 16723 2821 16787
rect 0 16705 2821 16723
rect 0 16641 135 16705
rect 199 16641 217 16705
rect 281 16641 299 16705
rect 363 16641 381 16705
rect 445 16641 463 16705
rect 527 16641 545 16705
rect 609 16641 627 16705
rect 691 16641 709 16705
rect 773 16641 791 16705
rect 855 16641 873 16705
rect 937 16641 955 16705
rect 1019 16641 1037 16705
rect 1101 16641 1119 16705
rect 1183 16641 1201 16705
rect 1265 16641 1283 16705
rect 1347 16641 1365 16705
rect 1429 16641 1447 16705
rect 1511 16641 1529 16705
rect 1593 16641 1611 16705
rect 1675 16641 1693 16705
rect 1757 16641 1775 16705
rect 1839 16641 1857 16705
rect 1921 16641 1939 16705
rect 2003 16641 2021 16705
rect 2085 16641 2103 16705
rect 2167 16641 2185 16705
rect 2249 16641 2267 16705
rect 2331 16641 2349 16705
rect 2413 16641 2431 16705
rect 2495 16641 2513 16705
rect 2577 16641 2594 16705
rect 2658 16641 2675 16705
rect 2739 16641 2756 16705
rect 2820 16641 2821 16705
rect 0 16623 2821 16641
rect 0 16559 135 16623
rect 199 16559 217 16623
rect 281 16559 299 16623
rect 363 16559 381 16623
rect 445 16559 463 16623
rect 527 16559 545 16623
rect 609 16559 627 16623
rect 691 16559 709 16623
rect 773 16559 791 16623
rect 855 16559 873 16623
rect 937 16559 955 16623
rect 1019 16559 1037 16623
rect 1101 16559 1119 16623
rect 1183 16559 1201 16623
rect 1265 16559 1283 16623
rect 1347 16559 1365 16623
rect 1429 16559 1447 16623
rect 1511 16559 1529 16623
rect 1593 16559 1611 16623
rect 1675 16559 1693 16623
rect 1757 16559 1775 16623
rect 1839 16559 1857 16623
rect 1921 16559 1939 16623
rect 2003 16559 2021 16623
rect 2085 16559 2103 16623
rect 2167 16559 2185 16623
rect 2249 16559 2267 16623
rect 2331 16559 2349 16623
rect 2413 16559 2431 16623
rect 2495 16559 2513 16623
rect 2577 16559 2594 16623
rect 2658 16559 2675 16623
rect 2739 16559 2756 16623
rect 2820 16559 2821 16623
rect 2875 17627 3771 17628
rect 2875 17563 2881 17627
rect 2945 17563 2963 17627
rect 3027 17563 3045 17627
rect 3109 17563 3127 17627
rect 3191 17563 3209 17627
rect 3273 17563 3291 17627
rect 3355 17563 3373 17627
rect 3437 17563 3455 17627
rect 3519 17563 3537 17627
rect 3601 17563 3619 17627
rect 3683 17563 3701 17627
rect 3765 17563 3771 17627
rect 2875 17546 3771 17563
rect 2875 17482 2881 17546
rect 2945 17482 2963 17546
rect 3027 17482 3045 17546
rect 3109 17482 3127 17546
rect 3191 17482 3209 17546
rect 3273 17482 3291 17546
rect 3355 17482 3373 17546
rect 3437 17482 3455 17546
rect 3519 17482 3537 17546
rect 3601 17482 3619 17546
rect 3683 17482 3701 17546
rect 3765 17482 3771 17546
rect 2875 17465 3771 17482
rect 2875 17401 2881 17465
rect 2945 17401 2963 17465
rect 3027 17401 3045 17465
rect 3109 17401 3127 17465
rect 3191 17401 3209 17465
rect 3273 17401 3291 17465
rect 3355 17401 3373 17465
rect 3437 17401 3455 17465
rect 3519 17401 3537 17465
rect 3601 17401 3619 17465
rect 3683 17401 3701 17465
rect 3765 17401 3771 17465
rect 11280 17627 12176 17628
rect 11280 17563 11286 17627
rect 11350 17563 11368 17627
rect 11432 17563 11450 17627
rect 11514 17563 11532 17627
rect 11596 17563 11614 17627
rect 11678 17563 11696 17627
rect 11760 17563 11778 17627
rect 11842 17563 11860 17627
rect 11924 17563 11942 17627
rect 12006 17563 12024 17627
rect 12088 17563 12106 17627
rect 12170 17563 12176 17627
rect 11280 17546 12176 17563
rect 11280 17482 11286 17546
rect 11350 17482 11368 17546
rect 11432 17482 11450 17546
rect 11514 17482 11532 17546
rect 11596 17482 11614 17546
rect 11678 17482 11696 17546
rect 11760 17482 11778 17546
rect 11842 17482 11860 17546
rect 11924 17482 11942 17546
rect 12006 17482 12024 17546
rect 12088 17482 12106 17546
rect 12170 17482 12176 17546
rect 11280 17465 12176 17482
rect 2875 17384 3771 17401
rect 2875 17320 2881 17384
rect 2945 17320 2963 17384
rect 3027 17320 3045 17384
rect 3109 17320 3127 17384
rect 3191 17320 3209 17384
rect 3273 17320 3291 17384
rect 3355 17320 3373 17384
rect 3437 17320 3455 17384
rect 3519 17320 3537 17384
rect 3601 17320 3619 17384
rect 3683 17320 3701 17384
rect 3765 17320 3771 17384
rect 2875 17303 3771 17320
rect 2875 17239 2881 17303
rect 2945 17239 2963 17303
rect 3027 17239 3045 17303
rect 3109 17239 3127 17303
rect 3191 17239 3209 17303
rect 3273 17239 3291 17303
rect 3355 17239 3373 17303
rect 3437 17239 3455 17303
rect 3519 17239 3537 17303
rect 3601 17239 3619 17303
rect 3683 17239 3701 17303
rect 3765 17239 3771 17303
rect 2875 17223 3771 17239
rect 2875 17159 2881 17223
rect 2945 17159 2963 17223
rect 3027 17159 3045 17223
rect 3109 17159 3127 17223
rect 3191 17159 3209 17223
rect 3273 17159 3291 17223
rect 3355 17159 3373 17223
rect 3437 17159 3455 17223
rect 3519 17159 3537 17223
rect 3601 17159 3619 17223
rect 3683 17159 3701 17223
rect 3765 17159 3771 17223
rect 3799 17402 4013 17403
rect 3799 17338 3800 17402
rect 3864 17338 3948 17402
rect 4012 17338 4013 17402
rect 3799 17314 4013 17338
rect 3799 17250 3800 17314
rect 3864 17250 3948 17314
rect 4012 17250 4013 17314
rect 3799 17227 4013 17250
rect 3799 17163 3800 17227
rect 3864 17163 3948 17227
rect 4012 17163 4013 17227
rect 3799 17162 4013 17163
rect 11038 17402 11252 17403
rect 11038 17338 11039 17402
rect 11103 17338 11187 17402
rect 11251 17338 11252 17402
rect 11038 17314 11252 17338
rect 11038 17250 11039 17314
rect 11103 17250 11187 17314
rect 11251 17250 11252 17314
rect 11038 17227 11252 17250
rect 11038 17163 11039 17227
rect 11103 17163 11187 17227
rect 11251 17163 11252 17227
rect 11038 17162 11252 17163
rect 11280 17401 11286 17465
rect 11350 17401 11368 17465
rect 11432 17401 11450 17465
rect 11514 17401 11532 17465
rect 11596 17401 11614 17465
rect 11678 17401 11696 17465
rect 11760 17401 11778 17465
rect 11842 17401 11860 17465
rect 11924 17401 11942 17465
rect 12006 17401 12024 17465
rect 12088 17401 12106 17465
rect 12170 17401 12176 17465
rect 11280 17384 12176 17401
rect 11280 17320 11286 17384
rect 11350 17320 11368 17384
rect 11432 17320 11450 17384
rect 11514 17320 11532 17384
rect 11596 17320 11614 17384
rect 11678 17320 11696 17384
rect 11760 17320 11778 17384
rect 11842 17320 11860 17384
rect 11924 17320 11942 17384
rect 12006 17320 12024 17384
rect 12088 17320 12106 17384
rect 12170 17320 12176 17384
rect 11280 17303 12176 17320
rect 11280 17239 11286 17303
rect 11350 17239 11368 17303
rect 11432 17239 11450 17303
rect 11514 17239 11532 17303
rect 11596 17239 11614 17303
rect 11678 17239 11696 17303
rect 11760 17239 11778 17303
rect 11842 17239 11860 17303
rect 11924 17239 11942 17303
rect 12006 17239 12024 17303
rect 12088 17239 12106 17303
rect 12170 17239 12176 17303
rect 11280 17223 12176 17239
rect 2875 17143 3771 17159
rect 2875 17079 2881 17143
rect 2945 17079 2963 17143
rect 3027 17079 3045 17143
rect 3109 17079 3127 17143
rect 3191 17079 3209 17143
rect 3273 17079 3291 17143
rect 3355 17079 3373 17143
rect 3437 17079 3455 17143
rect 3519 17079 3537 17143
rect 3601 17079 3619 17143
rect 3683 17079 3701 17143
rect 3765 17079 3771 17143
rect 11280 17159 11286 17223
rect 11350 17159 11368 17223
rect 11432 17159 11450 17223
rect 11514 17159 11532 17223
rect 11596 17159 11614 17223
rect 11678 17159 11696 17223
rect 11760 17159 11778 17223
rect 11842 17159 11860 17223
rect 11924 17159 11942 17223
rect 12006 17159 12024 17223
rect 12088 17159 12106 17223
rect 12170 17159 12176 17223
rect 11280 17143 12176 17159
rect 2875 17063 3771 17079
rect 2875 16999 2881 17063
rect 2945 16999 2963 17063
rect 3027 16999 3045 17063
rect 3109 16999 3127 17063
rect 3191 16999 3209 17063
rect 3273 16999 3291 17063
rect 3355 16999 3373 17063
rect 3437 16999 3455 17063
rect 3519 16999 3537 17063
rect 3601 16999 3619 17063
rect 3683 16999 3701 17063
rect 3765 16999 3771 17063
rect 2875 16983 3771 16999
rect 2875 16919 2881 16983
rect 2945 16919 2963 16983
rect 3027 16919 3045 16983
rect 3109 16919 3127 16983
rect 3191 16919 3209 16983
rect 3273 16919 3291 16983
rect 3355 16919 3373 16983
rect 3437 16919 3455 16983
rect 3519 16919 3537 16983
rect 3601 16919 3619 16983
rect 3683 16919 3701 16983
rect 3765 16919 3771 16983
rect 2875 16903 3771 16919
rect 2875 16839 2881 16903
rect 2945 16839 2963 16903
rect 3027 16839 3045 16903
rect 3109 16839 3127 16903
rect 3191 16839 3209 16903
rect 3273 16839 3291 16903
rect 3355 16839 3373 16903
rect 3437 16839 3455 16903
rect 3519 16839 3537 16903
rect 3601 16839 3619 16903
rect 3683 16839 3701 16903
rect 3765 16839 3771 16903
rect 2875 16823 3771 16839
rect 2875 16759 2881 16823
rect 2945 16759 2963 16823
rect 3027 16759 3045 16823
rect 3109 16759 3127 16823
rect 3191 16759 3209 16823
rect 3273 16759 3291 16823
rect 3355 16759 3373 16823
rect 3437 16759 3455 16823
rect 3519 16759 3537 16823
rect 3601 16759 3619 16823
rect 3683 16759 3701 16823
rect 3765 16759 3771 16823
rect 2875 16743 3771 16759
rect 2875 16679 2881 16743
rect 2945 16679 2963 16743
rect 3027 16679 3045 16743
rect 3109 16679 3127 16743
rect 3191 16679 3209 16743
rect 3273 16679 3291 16743
rect 3355 16679 3373 16743
rect 3437 16679 3455 16743
rect 3519 16679 3537 16743
rect 3601 16679 3619 16743
rect 3683 16679 3701 16743
rect 3765 16679 3771 16743
rect 2875 16663 3771 16679
rect 2875 16599 2881 16663
rect 2945 16599 2963 16663
rect 3027 16599 3045 16663
rect 3109 16599 3127 16663
rect 3191 16599 3209 16663
rect 3273 16599 3291 16663
rect 3355 16599 3373 16663
rect 3437 16599 3455 16663
rect 3519 16599 3537 16663
rect 3601 16599 3619 16663
rect 3683 16599 3701 16663
rect 3765 16599 3771 16663
rect 2875 16598 3771 16599
rect 3834 17117 4290 17118
rect 3834 17053 3838 17117
rect 3902 17053 3934 17117
rect 3998 17053 4030 17117
rect 4094 17053 4126 17117
rect 4190 17053 4222 17117
rect 4286 17053 4290 17117
rect 3834 17024 4290 17053
rect 3834 16960 3838 17024
rect 3902 16960 3934 17024
rect 3998 16960 4030 17024
rect 4094 16960 4126 17024
rect 4190 16960 4222 17024
rect 4286 16960 4290 17024
rect 3834 16931 4290 16960
rect 3834 16867 3838 16931
rect 3902 16867 3934 16931
rect 3998 16867 4030 16931
rect 4094 16867 4126 16931
rect 4190 16867 4222 16931
rect 4286 16867 4290 16931
rect 3834 16838 4290 16867
rect 10761 17117 11217 17118
rect 10761 17053 10765 17117
rect 10829 17053 10861 17117
rect 10925 17053 10957 17117
rect 11021 17053 11053 17117
rect 11117 17053 11149 17117
rect 11213 17053 11217 17117
rect 10761 17024 11217 17053
rect 10761 16960 10765 17024
rect 10829 16960 10861 17024
rect 10925 16960 10957 17024
rect 11021 16960 11053 17024
rect 11117 16960 11149 17024
rect 11213 16960 11217 17024
rect 10761 16931 11217 16960
rect 10761 16867 10765 16931
rect 10829 16867 10861 16931
rect 10925 16867 10957 16931
rect 11021 16867 11053 16931
rect 11117 16867 11149 16931
rect 11213 16867 11217 16931
rect 3834 16774 3838 16838
rect 3902 16774 3934 16838
rect 3998 16774 4030 16838
rect 4094 16774 4126 16838
rect 4190 16774 4222 16838
rect 4286 16774 4290 16838
rect 3834 16746 4290 16774
rect 3834 16682 3838 16746
rect 3902 16682 3934 16746
rect 3998 16682 4030 16746
rect 4094 16682 4126 16746
rect 4190 16682 4222 16746
rect 4286 16682 4290 16746
rect 3834 16654 4290 16682
rect 3834 16590 3838 16654
rect 3902 16590 3934 16654
rect 3998 16590 4030 16654
rect 4094 16590 4126 16654
rect 4190 16590 4222 16654
rect 4286 16590 4290 16654
rect 3834 16589 4290 16590
rect 4330 16856 4554 16857
rect 4330 16792 4331 16856
rect 4395 16792 4489 16856
rect 4553 16792 4554 16856
rect 4330 16746 4554 16792
rect 4330 16682 4331 16746
rect 4395 16682 4489 16746
rect 4553 16682 4554 16746
rect 4330 16636 4554 16682
rect 4330 16572 4331 16636
rect 4395 16572 4489 16636
rect 4553 16572 4554 16636
rect 4330 16571 4554 16572
rect 10497 16856 10721 16857
rect 10497 16792 10498 16856
rect 10562 16792 10656 16856
rect 10720 16792 10721 16856
rect 10497 16746 10721 16792
rect 10497 16682 10498 16746
rect 10562 16682 10656 16746
rect 10720 16682 10721 16746
rect 10497 16636 10721 16682
rect 10497 16572 10498 16636
rect 10562 16572 10656 16636
rect 10720 16572 10721 16636
rect 10761 16838 11217 16867
rect 10761 16774 10765 16838
rect 10829 16774 10861 16838
rect 10925 16774 10957 16838
rect 11021 16774 11053 16838
rect 11117 16774 11149 16838
rect 11213 16774 11217 16838
rect 10761 16746 11217 16774
rect 10761 16682 10765 16746
rect 10829 16682 10861 16746
rect 10925 16682 10957 16746
rect 11021 16682 11053 16746
rect 11117 16682 11149 16746
rect 11213 16682 11217 16746
rect 10761 16654 11217 16682
rect 10761 16590 10765 16654
rect 10829 16590 10861 16654
rect 10925 16590 10957 16654
rect 11021 16590 11053 16654
rect 11117 16590 11149 16654
rect 11213 16590 11217 16654
rect 11280 17079 11286 17143
rect 11350 17079 11368 17143
rect 11432 17079 11450 17143
rect 11514 17079 11532 17143
rect 11596 17079 11614 17143
rect 11678 17079 11696 17143
rect 11760 17079 11778 17143
rect 11842 17079 11860 17143
rect 11924 17079 11942 17143
rect 12006 17079 12024 17143
rect 12088 17079 12106 17143
rect 12170 17079 12176 17143
rect 11280 17063 12176 17079
rect 11280 16999 11286 17063
rect 11350 16999 11368 17063
rect 11432 16999 11450 17063
rect 11514 16999 11532 17063
rect 11596 16999 11614 17063
rect 11678 16999 11696 17063
rect 11760 16999 11778 17063
rect 11842 16999 11860 17063
rect 11924 16999 11942 17063
rect 12006 16999 12024 17063
rect 12088 16999 12106 17063
rect 12170 16999 12176 17063
rect 11280 16983 12176 16999
rect 11280 16919 11286 16983
rect 11350 16919 11368 16983
rect 11432 16919 11450 16983
rect 11514 16919 11532 16983
rect 11596 16919 11614 16983
rect 11678 16919 11696 16983
rect 11760 16919 11778 16983
rect 11842 16919 11860 16983
rect 11924 16919 11942 16983
rect 12006 16919 12024 16983
rect 12088 16919 12106 16983
rect 12170 16919 12176 16983
rect 11280 16903 12176 16919
rect 11280 16839 11286 16903
rect 11350 16839 11368 16903
rect 11432 16839 11450 16903
rect 11514 16839 11532 16903
rect 11596 16839 11614 16903
rect 11678 16839 11696 16903
rect 11760 16839 11778 16903
rect 11842 16839 11860 16903
rect 11924 16839 11942 16903
rect 12006 16839 12024 16903
rect 12088 16839 12106 16903
rect 12170 16839 12176 16903
rect 11280 16823 12176 16839
rect 11280 16759 11286 16823
rect 11350 16759 11368 16823
rect 11432 16759 11450 16823
rect 11514 16759 11532 16823
rect 11596 16759 11614 16823
rect 11678 16759 11696 16823
rect 11760 16759 11778 16823
rect 11842 16759 11860 16823
rect 11924 16759 11942 16823
rect 12006 16759 12024 16823
rect 12088 16759 12106 16823
rect 12170 16759 12176 16823
rect 11280 16743 12176 16759
rect 11280 16679 11286 16743
rect 11350 16679 11368 16743
rect 11432 16679 11450 16743
rect 11514 16679 11532 16743
rect 11596 16679 11614 16743
rect 11678 16679 11696 16743
rect 11760 16679 11778 16743
rect 11842 16679 11860 16743
rect 11924 16679 11942 16743
rect 12006 16679 12024 16743
rect 12088 16679 12106 16743
rect 12170 16679 12176 16743
rect 11280 16663 12176 16679
rect 11280 16599 11286 16663
rect 11350 16599 11368 16663
rect 11432 16599 11450 16663
rect 11514 16599 11532 16663
rect 11596 16599 11614 16663
rect 11678 16599 11696 16663
rect 11760 16599 11778 16663
rect 11842 16599 11860 16663
rect 11924 16599 11942 16663
rect 12006 16599 12024 16663
rect 12088 16599 12106 16663
rect 12170 16599 12176 16663
rect 11280 16598 12176 16599
rect 12230 17625 12231 17689
rect 12295 17625 12312 17689
rect 12376 17625 12393 17689
rect 12457 17625 12474 17689
rect 12538 17625 12556 17689
rect 12620 17625 12638 17689
rect 12702 17625 12720 17689
rect 12784 17625 12802 17689
rect 12866 17625 12884 17689
rect 12948 17625 12966 17689
rect 13030 17625 13048 17689
rect 13112 17625 13130 17689
rect 13194 17625 13212 17689
rect 13276 17625 13294 17689
rect 13358 17625 13376 17689
rect 13440 17625 13458 17689
rect 13522 17625 13540 17689
rect 13604 17625 13622 17689
rect 13686 17625 13704 17689
rect 13768 17625 13786 17689
rect 13850 17625 13868 17689
rect 13932 17625 13950 17689
rect 14014 17625 14032 17689
rect 14096 17625 14114 17689
rect 14178 17625 14196 17689
rect 14260 17625 14278 17689
rect 14342 17625 14360 17689
rect 14424 17625 14442 17689
rect 14506 17625 14524 17689
rect 14588 17625 14606 17689
rect 14670 17625 14688 17689
rect 14752 17625 14770 17689
rect 14834 17625 14852 17689
rect 14916 17625 15000 17689
rect 12230 17607 15000 17625
rect 12230 17543 12231 17607
rect 12295 17543 12312 17607
rect 12376 17543 12393 17607
rect 12457 17543 12474 17607
rect 12538 17543 12556 17607
rect 12620 17543 12638 17607
rect 12702 17543 12720 17607
rect 12784 17543 12802 17607
rect 12866 17543 12884 17607
rect 12948 17543 12966 17607
rect 13030 17543 13048 17607
rect 13112 17543 13130 17607
rect 13194 17543 13212 17607
rect 13276 17543 13294 17607
rect 13358 17543 13376 17607
rect 13440 17543 13458 17607
rect 13522 17543 13540 17607
rect 13604 17543 13622 17607
rect 13686 17543 13704 17607
rect 13768 17543 13786 17607
rect 13850 17543 13868 17607
rect 13932 17543 13950 17607
rect 14014 17543 14032 17607
rect 14096 17543 14114 17607
rect 14178 17543 14196 17607
rect 14260 17543 14278 17607
rect 14342 17543 14360 17607
rect 14424 17543 14442 17607
rect 14506 17543 14524 17607
rect 14588 17543 14606 17607
rect 14670 17543 14688 17607
rect 14752 17543 14770 17607
rect 14834 17543 14852 17607
rect 14916 17543 15000 17607
rect 12230 17525 15000 17543
rect 12230 17461 12231 17525
rect 12295 17461 12312 17525
rect 12376 17461 12393 17525
rect 12457 17461 12474 17525
rect 12538 17461 12556 17525
rect 12620 17461 12638 17525
rect 12702 17461 12720 17525
rect 12784 17461 12802 17525
rect 12866 17461 12884 17525
rect 12948 17461 12966 17525
rect 13030 17461 13048 17525
rect 13112 17461 13130 17525
rect 13194 17461 13212 17525
rect 13276 17461 13294 17525
rect 13358 17461 13376 17525
rect 13440 17461 13458 17525
rect 13522 17461 13540 17525
rect 13604 17461 13622 17525
rect 13686 17461 13704 17525
rect 13768 17461 13786 17525
rect 13850 17461 13868 17525
rect 13932 17461 13950 17525
rect 14014 17461 14032 17525
rect 14096 17461 14114 17525
rect 14178 17461 14196 17525
rect 14260 17461 14278 17525
rect 14342 17461 14360 17525
rect 14424 17461 14442 17525
rect 14506 17461 14524 17525
rect 14588 17461 14606 17525
rect 14670 17461 14688 17525
rect 14752 17461 14770 17525
rect 14834 17461 14852 17525
rect 14916 17461 15000 17525
rect 12230 17443 15000 17461
rect 12230 17379 12231 17443
rect 12295 17379 12312 17443
rect 12376 17379 12393 17443
rect 12457 17379 12474 17443
rect 12538 17379 12556 17443
rect 12620 17379 12638 17443
rect 12702 17379 12720 17443
rect 12784 17379 12802 17443
rect 12866 17379 12884 17443
rect 12948 17379 12966 17443
rect 13030 17379 13048 17443
rect 13112 17379 13130 17443
rect 13194 17379 13212 17443
rect 13276 17379 13294 17443
rect 13358 17379 13376 17443
rect 13440 17379 13458 17443
rect 13522 17379 13540 17443
rect 13604 17379 13622 17443
rect 13686 17379 13704 17443
rect 13768 17379 13786 17443
rect 13850 17379 13868 17443
rect 13932 17379 13950 17443
rect 14014 17379 14032 17443
rect 14096 17379 14114 17443
rect 14178 17379 14196 17443
rect 14260 17379 14278 17443
rect 14342 17379 14360 17443
rect 14424 17379 14442 17443
rect 14506 17379 14524 17443
rect 14588 17379 14606 17443
rect 14670 17379 14688 17443
rect 14752 17379 14770 17443
rect 14834 17379 14852 17443
rect 14916 17379 15000 17443
rect 12230 17361 15000 17379
rect 12230 17297 12231 17361
rect 12295 17297 12312 17361
rect 12376 17297 12393 17361
rect 12457 17297 12474 17361
rect 12538 17297 12556 17361
rect 12620 17297 12638 17361
rect 12702 17297 12720 17361
rect 12784 17297 12802 17361
rect 12866 17297 12884 17361
rect 12948 17297 12966 17361
rect 13030 17297 13048 17361
rect 13112 17297 13130 17361
rect 13194 17297 13212 17361
rect 13276 17297 13294 17361
rect 13358 17297 13376 17361
rect 13440 17297 13458 17361
rect 13522 17297 13540 17361
rect 13604 17297 13622 17361
rect 13686 17297 13704 17361
rect 13768 17297 13786 17361
rect 13850 17297 13868 17361
rect 13932 17297 13950 17361
rect 14014 17297 14032 17361
rect 14096 17297 14114 17361
rect 14178 17297 14196 17361
rect 14260 17297 14278 17361
rect 14342 17297 14360 17361
rect 14424 17297 14442 17361
rect 14506 17297 14524 17361
rect 14588 17297 14606 17361
rect 14670 17297 14688 17361
rect 14752 17297 14770 17361
rect 14834 17297 14852 17361
rect 14916 17297 15000 17361
rect 12230 17279 15000 17297
rect 12230 17215 12231 17279
rect 12295 17215 12312 17279
rect 12376 17215 12393 17279
rect 12457 17215 12474 17279
rect 12538 17215 12556 17279
rect 12620 17215 12638 17279
rect 12702 17215 12720 17279
rect 12784 17215 12802 17279
rect 12866 17215 12884 17279
rect 12948 17215 12966 17279
rect 13030 17215 13048 17279
rect 13112 17215 13130 17279
rect 13194 17215 13212 17279
rect 13276 17215 13294 17279
rect 13358 17215 13376 17279
rect 13440 17215 13458 17279
rect 13522 17215 13540 17279
rect 13604 17215 13622 17279
rect 13686 17215 13704 17279
rect 13768 17215 13786 17279
rect 13850 17215 13868 17279
rect 13932 17215 13950 17279
rect 14014 17215 14032 17279
rect 14096 17215 14114 17279
rect 14178 17215 14196 17279
rect 14260 17215 14278 17279
rect 14342 17215 14360 17279
rect 14424 17215 14442 17279
rect 14506 17215 14524 17279
rect 14588 17215 14606 17279
rect 14670 17215 14688 17279
rect 14752 17215 14770 17279
rect 14834 17215 14852 17279
rect 14916 17215 15000 17279
rect 12230 17197 15000 17215
rect 12230 17133 12231 17197
rect 12295 17133 12312 17197
rect 12376 17133 12393 17197
rect 12457 17133 12474 17197
rect 12538 17133 12556 17197
rect 12620 17133 12638 17197
rect 12702 17133 12720 17197
rect 12784 17133 12802 17197
rect 12866 17133 12884 17197
rect 12948 17133 12966 17197
rect 13030 17133 13048 17197
rect 13112 17133 13130 17197
rect 13194 17133 13212 17197
rect 13276 17133 13294 17197
rect 13358 17133 13376 17197
rect 13440 17133 13458 17197
rect 13522 17133 13540 17197
rect 13604 17133 13622 17197
rect 13686 17133 13704 17197
rect 13768 17133 13786 17197
rect 13850 17133 13868 17197
rect 13932 17133 13950 17197
rect 14014 17133 14032 17197
rect 14096 17133 14114 17197
rect 14178 17133 14196 17197
rect 14260 17133 14278 17197
rect 14342 17133 14360 17197
rect 14424 17133 14442 17197
rect 14506 17133 14524 17197
rect 14588 17133 14606 17197
rect 14670 17133 14688 17197
rect 14752 17133 14770 17197
rect 14834 17133 14852 17197
rect 14916 17133 15000 17197
rect 12230 17115 15000 17133
rect 12230 17051 12231 17115
rect 12295 17051 12312 17115
rect 12376 17051 12393 17115
rect 12457 17051 12474 17115
rect 12538 17051 12556 17115
rect 12620 17051 12638 17115
rect 12702 17051 12720 17115
rect 12784 17051 12802 17115
rect 12866 17051 12884 17115
rect 12948 17051 12966 17115
rect 13030 17051 13048 17115
rect 13112 17051 13130 17115
rect 13194 17051 13212 17115
rect 13276 17051 13294 17115
rect 13358 17051 13376 17115
rect 13440 17051 13458 17115
rect 13522 17051 13540 17115
rect 13604 17051 13622 17115
rect 13686 17051 13704 17115
rect 13768 17051 13786 17115
rect 13850 17051 13868 17115
rect 13932 17051 13950 17115
rect 14014 17051 14032 17115
rect 14096 17051 14114 17115
rect 14178 17051 14196 17115
rect 14260 17051 14278 17115
rect 14342 17051 14360 17115
rect 14424 17051 14442 17115
rect 14506 17051 14524 17115
rect 14588 17051 14606 17115
rect 14670 17051 14688 17115
rect 14752 17051 14770 17115
rect 14834 17051 14852 17115
rect 14916 17051 15000 17115
rect 12230 17033 15000 17051
rect 12230 16969 12231 17033
rect 12295 16969 12312 17033
rect 12376 16969 12393 17033
rect 12457 16969 12474 17033
rect 12538 16969 12556 17033
rect 12620 16969 12638 17033
rect 12702 16969 12720 17033
rect 12784 16969 12802 17033
rect 12866 16969 12884 17033
rect 12948 16969 12966 17033
rect 13030 16969 13048 17033
rect 13112 16969 13130 17033
rect 13194 16969 13212 17033
rect 13276 16969 13294 17033
rect 13358 16969 13376 17033
rect 13440 16969 13458 17033
rect 13522 16969 13540 17033
rect 13604 16969 13622 17033
rect 13686 16969 13704 17033
rect 13768 16969 13786 17033
rect 13850 16969 13868 17033
rect 13932 16969 13950 17033
rect 14014 16969 14032 17033
rect 14096 16969 14114 17033
rect 14178 16969 14196 17033
rect 14260 16969 14278 17033
rect 14342 16969 14360 17033
rect 14424 16969 14442 17033
rect 14506 16969 14524 17033
rect 14588 16969 14606 17033
rect 14670 16969 14688 17033
rect 14752 16969 14770 17033
rect 14834 16969 14852 17033
rect 14916 16969 15000 17033
rect 12230 16951 15000 16969
rect 12230 16887 12231 16951
rect 12295 16887 12312 16951
rect 12376 16887 12393 16951
rect 12457 16887 12474 16951
rect 12538 16887 12556 16951
rect 12620 16887 12638 16951
rect 12702 16887 12720 16951
rect 12784 16887 12802 16951
rect 12866 16887 12884 16951
rect 12948 16887 12966 16951
rect 13030 16887 13048 16951
rect 13112 16887 13130 16951
rect 13194 16887 13212 16951
rect 13276 16887 13294 16951
rect 13358 16887 13376 16951
rect 13440 16887 13458 16951
rect 13522 16887 13540 16951
rect 13604 16887 13622 16951
rect 13686 16887 13704 16951
rect 13768 16887 13786 16951
rect 13850 16887 13868 16951
rect 13932 16887 13950 16951
rect 14014 16887 14032 16951
rect 14096 16887 14114 16951
rect 14178 16887 14196 16951
rect 14260 16887 14278 16951
rect 14342 16887 14360 16951
rect 14424 16887 14442 16951
rect 14506 16887 14524 16951
rect 14588 16887 14606 16951
rect 14670 16887 14688 16951
rect 14752 16887 14770 16951
rect 14834 16887 14852 16951
rect 14916 16887 15000 16951
rect 12230 16869 15000 16887
rect 12230 16805 12231 16869
rect 12295 16805 12312 16869
rect 12376 16805 12393 16869
rect 12457 16805 12474 16869
rect 12538 16805 12556 16869
rect 12620 16805 12638 16869
rect 12702 16805 12720 16869
rect 12784 16805 12802 16869
rect 12866 16805 12884 16869
rect 12948 16805 12966 16869
rect 13030 16805 13048 16869
rect 13112 16805 13130 16869
rect 13194 16805 13212 16869
rect 13276 16805 13294 16869
rect 13358 16805 13376 16869
rect 13440 16805 13458 16869
rect 13522 16805 13540 16869
rect 13604 16805 13622 16869
rect 13686 16805 13704 16869
rect 13768 16805 13786 16869
rect 13850 16805 13868 16869
rect 13932 16805 13950 16869
rect 14014 16805 14032 16869
rect 14096 16805 14114 16869
rect 14178 16805 14196 16869
rect 14260 16805 14278 16869
rect 14342 16805 14360 16869
rect 14424 16805 14442 16869
rect 14506 16805 14524 16869
rect 14588 16805 14606 16869
rect 14670 16805 14688 16869
rect 14752 16805 14770 16869
rect 14834 16805 14852 16869
rect 14916 16805 15000 16869
rect 12230 16787 15000 16805
rect 12230 16723 12231 16787
rect 12295 16723 12312 16787
rect 12376 16723 12393 16787
rect 12457 16723 12474 16787
rect 12538 16723 12556 16787
rect 12620 16723 12638 16787
rect 12702 16723 12720 16787
rect 12784 16723 12802 16787
rect 12866 16723 12884 16787
rect 12948 16723 12966 16787
rect 13030 16723 13048 16787
rect 13112 16723 13130 16787
rect 13194 16723 13212 16787
rect 13276 16723 13294 16787
rect 13358 16723 13376 16787
rect 13440 16723 13458 16787
rect 13522 16723 13540 16787
rect 13604 16723 13622 16787
rect 13686 16723 13704 16787
rect 13768 16723 13786 16787
rect 13850 16723 13868 16787
rect 13932 16723 13950 16787
rect 14014 16723 14032 16787
rect 14096 16723 14114 16787
rect 14178 16723 14196 16787
rect 14260 16723 14278 16787
rect 14342 16723 14360 16787
rect 14424 16723 14442 16787
rect 14506 16723 14524 16787
rect 14588 16723 14606 16787
rect 14670 16723 14688 16787
rect 14752 16723 14770 16787
rect 14834 16723 14852 16787
rect 14916 16723 15000 16787
rect 12230 16705 15000 16723
rect 12230 16641 12231 16705
rect 12295 16641 12312 16705
rect 12376 16641 12393 16705
rect 12457 16641 12474 16705
rect 12538 16641 12556 16705
rect 12620 16641 12638 16705
rect 12702 16641 12720 16705
rect 12784 16641 12802 16705
rect 12866 16641 12884 16705
rect 12948 16641 12966 16705
rect 13030 16641 13048 16705
rect 13112 16641 13130 16705
rect 13194 16641 13212 16705
rect 13276 16641 13294 16705
rect 13358 16641 13376 16705
rect 13440 16641 13458 16705
rect 13522 16641 13540 16705
rect 13604 16641 13622 16705
rect 13686 16641 13704 16705
rect 13768 16641 13786 16705
rect 13850 16641 13868 16705
rect 13932 16641 13950 16705
rect 14014 16641 14032 16705
rect 14096 16641 14114 16705
rect 14178 16641 14196 16705
rect 14260 16641 14278 16705
rect 14342 16641 14360 16705
rect 14424 16641 14442 16705
rect 14506 16641 14524 16705
rect 14588 16641 14606 16705
rect 14670 16641 14688 16705
rect 14752 16641 14770 16705
rect 14834 16641 14852 16705
rect 14916 16641 15000 16705
rect 12230 16623 15000 16641
rect 10761 16589 11217 16590
rect 10497 16571 10721 16572
rect 0 16558 2821 16559
rect 12230 16559 12231 16623
rect 12295 16559 12312 16623
rect 12376 16559 12393 16623
rect 12457 16559 12474 16623
rect 12538 16559 12556 16623
rect 12620 16559 12638 16623
rect 12702 16559 12720 16623
rect 12784 16559 12802 16623
rect 12866 16559 12884 16623
rect 12948 16559 12966 16623
rect 13030 16559 13048 16623
rect 13112 16559 13130 16623
rect 13194 16559 13212 16623
rect 13276 16559 13294 16623
rect 13358 16559 13376 16623
rect 13440 16559 13458 16623
rect 13522 16559 13540 16623
rect 13604 16559 13622 16623
rect 13686 16559 13704 16623
rect 13768 16559 13786 16623
rect 13850 16559 13868 16623
rect 13932 16559 13950 16623
rect 14014 16559 14032 16623
rect 14096 16559 14114 16623
rect 14178 16559 14196 16623
rect 14260 16559 14278 16623
rect 14342 16559 14360 16623
rect 14424 16559 14442 16623
rect 14506 16559 14524 16623
rect 14588 16559 14606 16623
rect 14670 16559 14688 16623
rect 14752 16559 14770 16623
rect 14834 16559 14852 16623
rect 14916 16559 15000 16623
rect 0 16525 254 16558
rect 12230 16557 15000 16559
rect 14746 16525 15000 16557
rect 0 16524 4900 16525
rect 0 16460 157 16524
rect 221 16460 237 16524
rect 301 16460 317 16524
rect 381 16460 397 16524
rect 461 16460 477 16524
rect 541 16460 557 16524
rect 621 16460 637 16524
rect 701 16460 717 16524
rect 781 16460 797 16524
rect 861 16460 877 16524
rect 941 16460 957 16524
rect 1021 16460 1037 16524
rect 1101 16460 1117 16524
rect 1181 16460 1197 16524
rect 1261 16460 1277 16524
rect 1341 16460 1357 16524
rect 1421 16460 1437 16524
rect 1501 16460 1517 16524
rect 1581 16460 1597 16524
rect 1661 16460 1677 16524
rect 1741 16460 1757 16524
rect 1821 16460 1837 16524
rect 1901 16460 1917 16524
rect 1981 16460 1997 16524
rect 2061 16460 2077 16524
rect 2141 16460 2157 16524
rect 2221 16460 2237 16524
rect 2301 16460 2317 16524
rect 2381 16460 2397 16524
rect 2461 16460 2477 16524
rect 2541 16460 2557 16524
rect 2621 16460 2637 16524
rect 2701 16460 2717 16524
rect 2781 16460 2797 16524
rect 2861 16460 2877 16524
rect 2941 16460 2957 16524
rect 3021 16460 3037 16524
rect 3101 16460 3117 16524
rect 3181 16460 3197 16524
rect 3261 16460 3277 16524
rect 3341 16460 3357 16524
rect 3421 16460 3437 16524
rect 3501 16460 3517 16524
rect 3581 16460 3597 16524
rect 3661 16460 3677 16524
rect 3741 16460 3757 16524
rect 3821 16460 3837 16524
rect 3901 16460 3917 16524
rect 3981 16460 3997 16524
rect 4061 16460 4077 16524
rect 4141 16460 4157 16524
rect 4221 16460 4237 16524
rect 4301 16460 4317 16524
rect 4381 16460 4397 16524
rect 4461 16460 4477 16524
rect 4541 16460 4557 16524
rect 4621 16460 4637 16524
rect 4701 16460 4717 16524
rect 4781 16460 4797 16524
rect 4861 16460 4900 16524
rect 0 16443 4900 16460
rect 0 16379 157 16443
rect 221 16379 237 16443
rect 301 16379 317 16443
rect 381 16379 397 16443
rect 461 16379 477 16443
rect 541 16379 557 16443
rect 621 16379 637 16443
rect 701 16379 717 16443
rect 781 16379 797 16443
rect 861 16379 877 16443
rect 941 16379 957 16443
rect 1021 16379 1037 16443
rect 1101 16379 1117 16443
rect 1181 16379 1197 16443
rect 1261 16379 1277 16443
rect 1341 16379 1357 16443
rect 1421 16379 1437 16443
rect 1501 16379 1517 16443
rect 1581 16379 1597 16443
rect 1661 16379 1677 16443
rect 1741 16379 1757 16443
rect 1821 16379 1837 16443
rect 1901 16379 1917 16443
rect 1981 16379 1997 16443
rect 2061 16379 2077 16443
rect 2141 16379 2157 16443
rect 2221 16379 2237 16443
rect 2301 16379 2317 16443
rect 2381 16379 2397 16443
rect 2461 16379 2477 16443
rect 2541 16379 2557 16443
rect 2621 16379 2637 16443
rect 2701 16379 2717 16443
rect 2781 16379 2797 16443
rect 2861 16379 2877 16443
rect 2941 16379 2957 16443
rect 3021 16379 3037 16443
rect 3101 16379 3117 16443
rect 3181 16379 3197 16443
rect 3261 16379 3277 16443
rect 3341 16379 3357 16443
rect 3421 16379 3437 16443
rect 3501 16379 3517 16443
rect 3581 16379 3597 16443
rect 3661 16379 3677 16443
rect 3741 16379 3757 16443
rect 3821 16379 3837 16443
rect 3901 16379 3917 16443
rect 3981 16379 3997 16443
rect 4061 16379 4077 16443
rect 4141 16379 4157 16443
rect 4221 16379 4237 16443
rect 4301 16379 4317 16443
rect 4381 16379 4397 16443
rect 4461 16379 4477 16443
rect 4541 16379 4557 16443
rect 4621 16379 4637 16443
rect 4701 16379 4717 16443
rect 4781 16379 4797 16443
rect 4861 16379 4900 16443
rect 0 16362 4900 16379
rect 0 16298 157 16362
rect 221 16298 237 16362
rect 301 16298 317 16362
rect 381 16298 397 16362
rect 461 16298 477 16362
rect 541 16298 557 16362
rect 621 16298 637 16362
rect 701 16298 717 16362
rect 781 16298 797 16362
rect 861 16298 877 16362
rect 941 16298 957 16362
rect 1021 16298 1037 16362
rect 1101 16298 1117 16362
rect 1181 16298 1197 16362
rect 1261 16298 1277 16362
rect 1341 16298 1357 16362
rect 1421 16298 1437 16362
rect 1501 16298 1517 16362
rect 1581 16298 1597 16362
rect 1661 16298 1677 16362
rect 1741 16298 1757 16362
rect 1821 16298 1837 16362
rect 1901 16298 1917 16362
rect 1981 16298 1997 16362
rect 2061 16298 2077 16362
rect 2141 16298 2157 16362
rect 2221 16298 2237 16362
rect 2301 16298 2317 16362
rect 2381 16298 2397 16362
rect 2461 16298 2477 16362
rect 2541 16298 2557 16362
rect 2621 16298 2637 16362
rect 2701 16298 2717 16362
rect 2781 16298 2797 16362
rect 2861 16298 2877 16362
rect 2941 16298 2957 16362
rect 3021 16298 3037 16362
rect 3101 16298 3117 16362
rect 3181 16298 3197 16362
rect 3261 16298 3277 16362
rect 3341 16298 3357 16362
rect 3421 16298 3437 16362
rect 3501 16298 3517 16362
rect 3581 16298 3597 16362
rect 3661 16298 3677 16362
rect 3741 16298 3757 16362
rect 3821 16298 3837 16362
rect 3901 16298 3917 16362
rect 3981 16298 3997 16362
rect 4061 16298 4077 16362
rect 4141 16298 4157 16362
rect 4221 16298 4237 16362
rect 4301 16298 4317 16362
rect 4381 16298 4397 16362
rect 4461 16298 4477 16362
rect 4541 16298 4557 16362
rect 4621 16298 4637 16362
rect 4701 16298 4717 16362
rect 4781 16298 4797 16362
rect 4861 16298 4900 16362
rect 0 16281 4900 16298
rect 0 16217 157 16281
rect 221 16217 237 16281
rect 301 16217 317 16281
rect 381 16217 397 16281
rect 461 16217 477 16281
rect 541 16217 557 16281
rect 621 16217 637 16281
rect 701 16217 717 16281
rect 781 16217 797 16281
rect 861 16217 877 16281
rect 941 16217 957 16281
rect 1021 16217 1037 16281
rect 1101 16217 1117 16281
rect 1181 16217 1197 16281
rect 1261 16217 1277 16281
rect 1341 16217 1357 16281
rect 1421 16217 1437 16281
rect 1501 16217 1517 16281
rect 1581 16217 1597 16281
rect 1661 16217 1677 16281
rect 1741 16217 1757 16281
rect 1821 16217 1837 16281
rect 1901 16217 1917 16281
rect 1981 16217 1997 16281
rect 2061 16217 2077 16281
rect 2141 16217 2157 16281
rect 2221 16217 2237 16281
rect 2301 16217 2317 16281
rect 2381 16217 2397 16281
rect 2461 16217 2477 16281
rect 2541 16217 2557 16281
rect 2621 16217 2637 16281
rect 2701 16217 2717 16281
rect 2781 16217 2797 16281
rect 2861 16217 2877 16281
rect 2941 16217 2957 16281
rect 3021 16217 3037 16281
rect 3101 16217 3117 16281
rect 3181 16217 3197 16281
rect 3261 16217 3277 16281
rect 3341 16217 3357 16281
rect 3421 16217 3437 16281
rect 3501 16217 3517 16281
rect 3581 16217 3597 16281
rect 3661 16217 3677 16281
rect 3741 16217 3757 16281
rect 3821 16217 3837 16281
rect 3901 16217 3917 16281
rect 3981 16217 3997 16281
rect 4061 16217 4077 16281
rect 4141 16217 4157 16281
rect 4221 16217 4237 16281
rect 4301 16217 4317 16281
rect 4381 16217 4397 16281
rect 4461 16217 4477 16281
rect 4541 16217 4557 16281
rect 4621 16217 4637 16281
rect 4701 16217 4717 16281
rect 4781 16217 4797 16281
rect 4861 16217 4900 16281
rect 0 16200 4900 16217
rect 0 16136 157 16200
rect 221 16136 237 16200
rect 301 16136 317 16200
rect 381 16136 397 16200
rect 461 16136 477 16200
rect 541 16136 557 16200
rect 621 16136 637 16200
rect 701 16136 717 16200
rect 781 16136 797 16200
rect 861 16136 877 16200
rect 941 16136 957 16200
rect 1021 16136 1037 16200
rect 1101 16136 1117 16200
rect 1181 16136 1197 16200
rect 1261 16136 1277 16200
rect 1341 16136 1357 16200
rect 1421 16136 1437 16200
rect 1501 16136 1517 16200
rect 1581 16136 1597 16200
rect 1661 16136 1677 16200
rect 1741 16136 1757 16200
rect 1821 16136 1837 16200
rect 1901 16136 1917 16200
rect 1981 16136 1997 16200
rect 2061 16136 2077 16200
rect 2141 16136 2157 16200
rect 2221 16136 2237 16200
rect 2301 16136 2317 16200
rect 2381 16136 2397 16200
rect 2461 16136 2477 16200
rect 2541 16136 2557 16200
rect 2621 16136 2637 16200
rect 2701 16136 2717 16200
rect 2781 16136 2797 16200
rect 2861 16136 2877 16200
rect 2941 16136 2957 16200
rect 3021 16136 3037 16200
rect 3101 16136 3117 16200
rect 3181 16136 3197 16200
rect 3261 16136 3277 16200
rect 3341 16136 3357 16200
rect 3421 16136 3437 16200
rect 3501 16136 3517 16200
rect 3581 16136 3597 16200
rect 3661 16136 3677 16200
rect 3741 16136 3757 16200
rect 3821 16136 3837 16200
rect 3901 16136 3917 16200
rect 3981 16136 3997 16200
rect 4061 16136 4077 16200
rect 4141 16136 4157 16200
rect 4221 16136 4237 16200
rect 4301 16136 4317 16200
rect 4381 16136 4397 16200
rect 4461 16136 4477 16200
rect 4541 16136 4557 16200
rect 4621 16136 4637 16200
rect 4701 16136 4717 16200
rect 4781 16136 4797 16200
rect 4861 16136 4900 16200
rect 0 16119 4900 16136
rect 0 16055 157 16119
rect 221 16055 237 16119
rect 301 16055 317 16119
rect 381 16055 397 16119
rect 461 16055 477 16119
rect 541 16055 557 16119
rect 621 16055 637 16119
rect 701 16055 717 16119
rect 781 16055 797 16119
rect 861 16055 877 16119
rect 941 16055 957 16119
rect 1021 16055 1037 16119
rect 1101 16055 1117 16119
rect 1181 16055 1197 16119
rect 1261 16055 1277 16119
rect 1341 16055 1357 16119
rect 1421 16055 1437 16119
rect 1501 16055 1517 16119
rect 1581 16055 1597 16119
rect 1661 16055 1677 16119
rect 1741 16055 1757 16119
rect 1821 16055 1837 16119
rect 1901 16055 1917 16119
rect 1981 16055 1997 16119
rect 2061 16055 2077 16119
rect 2141 16055 2157 16119
rect 2221 16055 2237 16119
rect 2301 16055 2317 16119
rect 2381 16055 2397 16119
rect 2461 16055 2477 16119
rect 2541 16055 2557 16119
rect 2621 16055 2637 16119
rect 2701 16055 2717 16119
rect 2781 16055 2797 16119
rect 2861 16055 2877 16119
rect 2941 16055 2957 16119
rect 3021 16055 3037 16119
rect 3101 16055 3117 16119
rect 3181 16055 3197 16119
rect 3261 16055 3277 16119
rect 3341 16055 3357 16119
rect 3421 16055 3437 16119
rect 3501 16055 3517 16119
rect 3581 16055 3597 16119
rect 3661 16055 3677 16119
rect 3741 16055 3757 16119
rect 3821 16055 3837 16119
rect 3901 16055 3917 16119
rect 3981 16055 3997 16119
rect 4061 16055 4077 16119
rect 4141 16055 4157 16119
rect 4221 16055 4237 16119
rect 4301 16055 4317 16119
rect 4381 16055 4397 16119
rect 4461 16055 4477 16119
rect 4541 16055 4557 16119
rect 4621 16055 4637 16119
rect 4701 16055 4717 16119
rect 4781 16055 4797 16119
rect 4861 16055 4900 16119
rect 0 16038 4900 16055
rect 0 15974 157 16038
rect 221 15974 237 16038
rect 301 15974 317 16038
rect 381 15974 397 16038
rect 461 15974 477 16038
rect 541 15974 557 16038
rect 621 15974 637 16038
rect 701 15974 717 16038
rect 781 15974 797 16038
rect 861 15974 877 16038
rect 941 15974 957 16038
rect 1021 15974 1037 16038
rect 1101 15974 1117 16038
rect 1181 15974 1197 16038
rect 1261 15974 1277 16038
rect 1341 15974 1357 16038
rect 1421 15974 1437 16038
rect 1501 15974 1517 16038
rect 1581 15974 1597 16038
rect 1661 15974 1677 16038
rect 1741 15974 1757 16038
rect 1821 15974 1837 16038
rect 1901 15974 1917 16038
rect 1981 15974 1997 16038
rect 2061 15974 2077 16038
rect 2141 15974 2157 16038
rect 2221 15974 2237 16038
rect 2301 15974 2317 16038
rect 2381 15974 2397 16038
rect 2461 15974 2477 16038
rect 2541 15974 2557 16038
rect 2621 15974 2637 16038
rect 2701 15974 2717 16038
rect 2781 15974 2797 16038
rect 2861 15974 2877 16038
rect 2941 15974 2957 16038
rect 3021 15974 3037 16038
rect 3101 15974 3117 16038
rect 3181 15974 3197 16038
rect 3261 15974 3277 16038
rect 3341 15974 3357 16038
rect 3421 15974 3437 16038
rect 3501 15974 3517 16038
rect 3581 15974 3597 16038
rect 3661 15974 3677 16038
rect 3741 15974 3757 16038
rect 3821 15974 3837 16038
rect 3901 15974 3917 16038
rect 3981 15974 3997 16038
rect 4061 15974 4077 16038
rect 4141 15974 4157 16038
rect 4221 15974 4237 16038
rect 4301 15974 4317 16038
rect 4381 15974 4397 16038
rect 4461 15974 4477 16038
rect 4541 15974 4557 16038
rect 4621 15974 4637 16038
rect 4701 15974 4717 16038
rect 4781 15974 4797 16038
rect 4861 15974 4900 16038
rect 0 15957 4900 15974
rect 0 15893 157 15957
rect 221 15893 237 15957
rect 301 15893 317 15957
rect 381 15893 397 15957
rect 461 15893 477 15957
rect 541 15893 557 15957
rect 621 15893 637 15957
rect 701 15893 717 15957
rect 781 15893 797 15957
rect 861 15893 877 15957
rect 941 15893 957 15957
rect 1021 15893 1037 15957
rect 1101 15893 1117 15957
rect 1181 15893 1197 15957
rect 1261 15893 1277 15957
rect 1341 15893 1357 15957
rect 1421 15893 1437 15957
rect 1501 15893 1517 15957
rect 1581 15893 1597 15957
rect 1661 15893 1677 15957
rect 1741 15893 1757 15957
rect 1821 15893 1837 15957
rect 1901 15893 1917 15957
rect 1981 15893 1997 15957
rect 2061 15893 2077 15957
rect 2141 15893 2157 15957
rect 2221 15893 2237 15957
rect 2301 15893 2317 15957
rect 2381 15893 2397 15957
rect 2461 15893 2477 15957
rect 2541 15893 2557 15957
rect 2621 15893 2637 15957
rect 2701 15893 2717 15957
rect 2781 15893 2797 15957
rect 2861 15893 2877 15957
rect 2941 15893 2957 15957
rect 3021 15893 3037 15957
rect 3101 15893 3117 15957
rect 3181 15893 3197 15957
rect 3261 15893 3277 15957
rect 3341 15893 3357 15957
rect 3421 15893 3437 15957
rect 3501 15893 3517 15957
rect 3581 15893 3597 15957
rect 3661 15893 3677 15957
rect 3741 15893 3757 15957
rect 3821 15893 3837 15957
rect 3901 15893 3917 15957
rect 3981 15893 3997 15957
rect 4061 15893 4077 15957
rect 4141 15893 4157 15957
rect 4221 15893 4237 15957
rect 4301 15893 4317 15957
rect 4381 15893 4397 15957
rect 4461 15893 4477 15957
rect 4541 15893 4557 15957
rect 4621 15893 4637 15957
rect 4701 15893 4717 15957
rect 4781 15893 4797 15957
rect 4861 15893 4900 15957
rect 0 15876 4900 15893
rect 0 15812 157 15876
rect 221 15812 237 15876
rect 301 15812 317 15876
rect 381 15812 397 15876
rect 461 15812 477 15876
rect 541 15812 557 15876
rect 621 15812 637 15876
rect 701 15812 717 15876
rect 781 15812 797 15876
rect 861 15812 877 15876
rect 941 15812 957 15876
rect 1021 15812 1037 15876
rect 1101 15812 1117 15876
rect 1181 15812 1197 15876
rect 1261 15812 1277 15876
rect 1341 15812 1357 15876
rect 1421 15812 1437 15876
rect 1501 15812 1517 15876
rect 1581 15812 1597 15876
rect 1661 15812 1677 15876
rect 1741 15812 1757 15876
rect 1821 15812 1837 15876
rect 1901 15812 1917 15876
rect 1981 15812 1997 15876
rect 2061 15812 2077 15876
rect 2141 15812 2157 15876
rect 2221 15812 2237 15876
rect 2301 15812 2317 15876
rect 2381 15812 2397 15876
rect 2461 15812 2477 15876
rect 2541 15812 2557 15876
rect 2621 15812 2637 15876
rect 2701 15812 2717 15876
rect 2781 15812 2797 15876
rect 2861 15812 2877 15876
rect 2941 15812 2957 15876
rect 3021 15812 3037 15876
rect 3101 15812 3117 15876
rect 3181 15812 3197 15876
rect 3261 15812 3277 15876
rect 3341 15812 3357 15876
rect 3421 15812 3437 15876
rect 3501 15812 3517 15876
rect 3581 15812 3597 15876
rect 3661 15812 3677 15876
rect 3741 15812 3757 15876
rect 3821 15812 3837 15876
rect 3901 15812 3917 15876
rect 3981 15812 3997 15876
rect 4061 15812 4077 15876
rect 4141 15812 4157 15876
rect 4221 15812 4237 15876
rect 4301 15812 4317 15876
rect 4381 15812 4397 15876
rect 4461 15812 4477 15876
rect 4541 15812 4557 15876
rect 4621 15812 4637 15876
rect 4701 15812 4717 15876
rect 4781 15812 4797 15876
rect 4861 15812 4900 15876
rect 0 15795 4900 15812
rect 0 15731 157 15795
rect 221 15731 237 15795
rect 301 15731 317 15795
rect 381 15731 397 15795
rect 461 15731 477 15795
rect 541 15731 557 15795
rect 621 15731 637 15795
rect 701 15731 717 15795
rect 781 15731 797 15795
rect 861 15731 877 15795
rect 941 15731 957 15795
rect 1021 15731 1037 15795
rect 1101 15731 1117 15795
rect 1181 15731 1197 15795
rect 1261 15731 1277 15795
rect 1341 15731 1357 15795
rect 1421 15731 1437 15795
rect 1501 15731 1517 15795
rect 1581 15731 1597 15795
rect 1661 15731 1677 15795
rect 1741 15731 1757 15795
rect 1821 15731 1837 15795
rect 1901 15731 1917 15795
rect 1981 15731 1997 15795
rect 2061 15731 2077 15795
rect 2141 15731 2157 15795
rect 2221 15731 2237 15795
rect 2301 15731 2317 15795
rect 2381 15731 2397 15795
rect 2461 15731 2477 15795
rect 2541 15731 2557 15795
rect 2621 15731 2637 15795
rect 2701 15731 2717 15795
rect 2781 15731 2797 15795
rect 2861 15731 2877 15795
rect 2941 15731 2957 15795
rect 3021 15731 3037 15795
rect 3101 15731 3117 15795
rect 3181 15731 3197 15795
rect 3261 15731 3277 15795
rect 3341 15731 3357 15795
rect 3421 15731 3437 15795
rect 3501 15731 3517 15795
rect 3581 15731 3597 15795
rect 3661 15731 3677 15795
rect 3741 15731 3757 15795
rect 3821 15731 3837 15795
rect 3901 15731 3917 15795
rect 3981 15731 3997 15795
rect 4061 15731 4077 15795
rect 4141 15731 4157 15795
rect 4221 15731 4237 15795
rect 4301 15731 4317 15795
rect 4381 15731 4397 15795
rect 4461 15731 4477 15795
rect 4541 15731 4557 15795
rect 4621 15731 4637 15795
rect 4701 15731 4717 15795
rect 4781 15731 4797 15795
rect 4861 15731 4900 15795
rect 0 15714 4900 15731
rect 0 15650 157 15714
rect 221 15650 237 15714
rect 301 15650 317 15714
rect 381 15650 397 15714
rect 461 15650 477 15714
rect 541 15650 557 15714
rect 621 15650 637 15714
rect 701 15650 717 15714
rect 781 15650 797 15714
rect 861 15650 877 15714
rect 941 15650 957 15714
rect 1021 15650 1037 15714
rect 1101 15650 1117 15714
rect 1181 15650 1197 15714
rect 1261 15650 1277 15714
rect 1341 15650 1357 15714
rect 1421 15650 1437 15714
rect 1501 15650 1517 15714
rect 1581 15650 1597 15714
rect 1661 15650 1677 15714
rect 1741 15650 1757 15714
rect 1821 15650 1837 15714
rect 1901 15650 1917 15714
rect 1981 15650 1997 15714
rect 2061 15650 2077 15714
rect 2141 15650 2157 15714
rect 2221 15650 2237 15714
rect 2301 15650 2317 15714
rect 2381 15650 2397 15714
rect 2461 15650 2477 15714
rect 2541 15650 2557 15714
rect 2621 15650 2637 15714
rect 2701 15650 2717 15714
rect 2781 15650 2797 15714
rect 2861 15650 2877 15714
rect 2941 15650 2957 15714
rect 3021 15650 3037 15714
rect 3101 15650 3117 15714
rect 3181 15650 3197 15714
rect 3261 15650 3277 15714
rect 3341 15650 3357 15714
rect 3421 15650 3437 15714
rect 3501 15650 3517 15714
rect 3581 15650 3597 15714
rect 3661 15650 3677 15714
rect 3741 15650 3757 15714
rect 3821 15650 3837 15714
rect 3901 15650 3917 15714
rect 3981 15650 3997 15714
rect 4061 15650 4077 15714
rect 4141 15650 4157 15714
rect 4221 15650 4237 15714
rect 4301 15650 4317 15714
rect 4381 15650 4397 15714
rect 4461 15650 4477 15714
rect 4541 15650 4557 15714
rect 4621 15650 4637 15714
rect 4701 15650 4717 15714
rect 4781 15650 4797 15714
rect 4861 15650 4900 15714
rect 0 15633 4900 15650
rect 0 15569 157 15633
rect 221 15569 237 15633
rect 301 15569 317 15633
rect 381 15569 397 15633
rect 461 15569 477 15633
rect 541 15569 557 15633
rect 621 15569 637 15633
rect 701 15569 717 15633
rect 781 15569 797 15633
rect 861 15569 877 15633
rect 941 15569 957 15633
rect 1021 15569 1037 15633
rect 1101 15569 1117 15633
rect 1181 15569 1197 15633
rect 1261 15569 1277 15633
rect 1341 15569 1357 15633
rect 1421 15569 1437 15633
rect 1501 15569 1517 15633
rect 1581 15569 1597 15633
rect 1661 15569 1677 15633
rect 1741 15569 1757 15633
rect 1821 15569 1837 15633
rect 1901 15569 1917 15633
rect 1981 15569 1997 15633
rect 2061 15569 2077 15633
rect 2141 15569 2157 15633
rect 2221 15569 2237 15633
rect 2301 15569 2317 15633
rect 2381 15569 2397 15633
rect 2461 15569 2477 15633
rect 2541 15569 2557 15633
rect 2621 15569 2637 15633
rect 2701 15569 2717 15633
rect 2781 15569 2797 15633
rect 2861 15569 2877 15633
rect 2941 15569 2957 15633
rect 3021 15569 3037 15633
rect 3101 15569 3117 15633
rect 3181 15569 3197 15633
rect 3261 15569 3277 15633
rect 3341 15569 3357 15633
rect 3421 15569 3437 15633
rect 3501 15569 3517 15633
rect 3581 15569 3597 15633
rect 3661 15569 3677 15633
rect 3741 15569 3757 15633
rect 3821 15569 3837 15633
rect 3901 15569 3917 15633
rect 3981 15569 3997 15633
rect 4061 15569 4077 15633
rect 4141 15569 4157 15633
rect 4221 15569 4237 15633
rect 4301 15569 4317 15633
rect 4381 15569 4397 15633
rect 4461 15569 4477 15633
rect 4541 15569 4557 15633
rect 4621 15569 4637 15633
rect 4701 15569 4717 15633
rect 4781 15569 4797 15633
rect 4861 15569 4900 15633
rect 0 15552 4900 15569
rect 0 15488 157 15552
rect 221 15488 237 15552
rect 301 15488 317 15552
rect 381 15488 397 15552
rect 461 15488 477 15552
rect 541 15488 557 15552
rect 621 15488 637 15552
rect 701 15488 717 15552
rect 781 15488 797 15552
rect 861 15488 877 15552
rect 941 15488 957 15552
rect 1021 15488 1037 15552
rect 1101 15488 1117 15552
rect 1181 15488 1197 15552
rect 1261 15488 1277 15552
rect 1341 15488 1357 15552
rect 1421 15488 1437 15552
rect 1501 15488 1517 15552
rect 1581 15488 1597 15552
rect 1661 15488 1677 15552
rect 1741 15488 1757 15552
rect 1821 15488 1837 15552
rect 1901 15488 1917 15552
rect 1981 15488 1997 15552
rect 2061 15488 2077 15552
rect 2141 15488 2157 15552
rect 2221 15488 2237 15552
rect 2301 15488 2317 15552
rect 2381 15488 2397 15552
rect 2461 15488 2477 15552
rect 2541 15488 2557 15552
rect 2621 15488 2637 15552
rect 2701 15488 2717 15552
rect 2781 15488 2797 15552
rect 2861 15488 2877 15552
rect 2941 15488 2957 15552
rect 3021 15488 3037 15552
rect 3101 15488 3117 15552
rect 3181 15488 3197 15552
rect 3261 15488 3277 15552
rect 3341 15488 3357 15552
rect 3421 15488 3437 15552
rect 3501 15488 3517 15552
rect 3581 15488 3597 15552
rect 3661 15488 3677 15552
rect 3741 15488 3757 15552
rect 3821 15488 3837 15552
rect 3901 15488 3917 15552
rect 3981 15488 3997 15552
rect 4061 15488 4077 15552
rect 4141 15488 4157 15552
rect 4221 15488 4237 15552
rect 4301 15488 4317 15552
rect 4381 15488 4397 15552
rect 4461 15488 4477 15552
rect 4541 15488 4557 15552
rect 4621 15488 4637 15552
rect 4701 15488 4717 15552
rect 4781 15488 4797 15552
rect 4861 15488 4900 15552
rect 0 15471 4900 15488
rect 0 15407 157 15471
rect 221 15407 237 15471
rect 301 15407 317 15471
rect 381 15407 397 15471
rect 461 15407 477 15471
rect 541 15407 557 15471
rect 621 15407 637 15471
rect 701 15407 717 15471
rect 781 15407 797 15471
rect 861 15407 877 15471
rect 941 15407 957 15471
rect 1021 15407 1037 15471
rect 1101 15407 1117 15471
rect 1181 15407 1197 15471
rect 1261 15407 1277 15471
rect 1341 15407 1357 15471
rect 1421 15407 1437 15471
rect 1501 15407 1517 15471
rect 1581 15407 1597 15471
rect 1661 15407 1677 15471
rect 1741 15407 1757 15471
rect 1821 15407 1837 15471
rect 1901 15407 1917 15471
rect 1981 15407 1997 15471
rect 2061 15407 2077 15471
rect 2141 15407 2157 15471
rect 2221 15407 2237 15471
rect 2301 15407 2317 15471
rect 2381 15407 2397 15471
rect 2461 15407 2477 15471
rect 2541 15407 2557 15471
rect 2621 15407 2637 15471
rect 2701 15407 2717 15471
rect 2781 15407 2797 15471
rect 2861 15407 2877 15471
rect 2941 15407 2957 15471
rect 3021 15407 3037 15471
rect 3101 15407 3117 15471
rect 3181 15407 3197 15471
rect 3261 15407 3277 15471
rect 3341 15407 3357 15471
rect 3421 15407 3437 15471
rect 3501 15407 3517 15471
rect 3581 15407 3597 15471
rect 3661 15407 3677 15471
rect 3741 15407 3757 15471
rect 3821 15407 3837 15471
rect 3901 15407 3917 15471
rect 3981 15407 3997 15471
rect 4061 15407 4077 15471
rect 4141 15407 4157 15471
rect 4221 15407 4237 15471
rect 4301 15407 4317 15471
rect 4381 15407 4397 15471
rect 4461 15407 4477 15471
rect 4541 15407 4557 15471
rect 4621 15407 4637 15471
rect 4701 15407 4717 15471
rect 4781 15407 4797 15471
rect 4861 15407 4900 15471
rect 0 15390 4900 15407
rect 0 15326 157 15390
rect 221 15326 237 15390
rect 301 15326 317 15390
rect 381 15326 397 15390
rect 461 15326 477 15390
rect 541 15326 557 15390
rect 621 15326 637 15390
rect 701 15326 717 15390
rect 781 15326 797 15390
rect 861 15326 877 15390
rect 941 15326 957 15390
rect 1021 15326 1037 15390
rect 1101 15326 1117 15390
rect 1181 15326 1197 15390
rect 1261 15326 1277 15390
rect 1341 15326 1357 15390
rect 1421 15326 1437 15390
rect 1501 15326 1517 15390
rect 1581 15326 1597 15390
rect 1661 15326 1677 15390
rect 1741 15326 1757 15390
rect 1821 15326 1837 15390
rect 1901 15326 1917 15390
rect 1981 15326 1997 15390
rect 2061 15326 2077 15390
rect 2141 15326 2157 15390
rect 2221 15326 2237 15390
rect 2301 15326 2317 15390
rect 2381 15326 2397 15390
rect 2461 15326 2477 15390
rect 2541 15326 2557 15390
rect 2621 15326 2637 15390
rect 2701 15326 2717 15390
rect 2781 15326 2797 15390
rect 2861 15326 2877 15390
rect 2941 15326 2957 15390
rect 3021 15326 3037 15390
rect 3101 15326 3117 15390
rect 3181 15326 3197 15390
rect 3261 15326 3277 15390
rect 3341 15326 3357 15390
rect 3421 15326 3437 15390
rect 3501 15326 3517 15390
rect 3581 15326 3597 15390
rect 3661 15326 3677 15390
rect 3741 15326 3757 15390
rect 3821 15326 3837 15390
rect 3901 15326 3917 15390
rect 3981 15326 3997 15390
rect 4061 15326 4077 15390
rect 4141 15326 4157 15390
rect 4221 15326 4237 15390
rect 4301 15326 4317 15390
rect 4381 15326 4397 15390
rect 4461 15326 4477 15390
rect 4541 15326 4557 15390
rect 4621 15326 4637 15390
rect 4701 15326 4717 15390
rect 4781 15326 4797 15390
rect 4861 15326 4900 15390
rect 0 15309 4900 15326
rect 0 15245 157 15309
rect 221 15245 237 15309
rect 301 15245 317 15309
rect 381 15245 397 15309
rect 461 15245 477 15309
rect 541 15245 557 15309
rect 621 15245 637 15309
rect 701 15245 717 15309
rect 781 15245 797 15309
rect 861 15245 877 15309
rect 941 15245 957 15309
rect 1021 15245 1037 15309
rect 1101 15245 1117 15309
rect 1181 15245 1197 15309
rect 1261 15245 1277 15309
rect 1341 15245 1357 15309
rect 1421 15245 1437 15309
rect 1501 15245 1517 15309
rect 1581 15245 1597 15309
rect 1661 15245 1677 15309
rect 1741 15245 1757 15309
rect 1821 15245 1837 15309
rect 1901 15245 1917 15309
rect 1981 15245 1997 15309
rect 2061 15245 2077 15309
rect 2141 15245 2157 15309
rect 2221 15245 2237 15309
rect 2301 15245 2317 15309
rect 2381 15245 2397 15309
rect 2461 15245 2477 15309
rect 2541 15245 2557 15309
rect 2621 15245 2637 15309
rect 2701 15245 2717 15309
rect 2781 15245 2797 15309
rect 2861 15245 2877 15309
rect 2941 15245 2957 15309
rect 3021 15245 3037 15309
rect 3101 15245 3117 15309
rect 3181 15245 3197 15309
rect 3261 15245 3277 15309
rect 3341 15245 3357 15309
rect 3421 15245 3437 15309
rect 3501 15245 3517 15309
rect 3581 15245 3597 15309
rect 3661 15245 3677 15309
rect 3741 15245 3757 15309
rect 3821 15245 3837 15309
rect 3901 15245 3917 15309
rect 3981 15245 3997 15309
rect 4061 15245 4077 15309
rect 4141 15245 4157 15309
rect 4221 15245 4237 15309
rect 4301 15245 4317 15309
rect 4381 15245 4397 15309
rect 4461 15245 4477 15309
rect 4541 15245 4557 15309
rect 4621 15245 4637 15309
rect 4701 15245 4717 15309
rect 4781 15245 4797 15309
rect 4861 15245 4900 15309
rect 0 15228 4900 15245
rect 0 15164 157 15228
rect 221 15164 237 15228
rect 301 15164 317 15228
rect 381 15164 397 15228
rect 461 15164 477 15228
rect 541 15164 557 15228
rect 621 15164 637 15228
rect 701 15164 717 15228
rect 781 15164 797 15228
rect 861 15164 877 15228
rect 941 15164 957 15228
rect 1021 15164 1037 15228
rect 1101 15164 1117 15228
rect 1181 15164 1197 15228
rect 1261 15164 1277 15228
rect 1341 15164 1357 15228
rect 1421 15164 1437 15228
rect 1501 15164 1517 15228
rect 1581 15164 1597 15228
rect 1661 15164 1677 15228
rect 1741 15164 1757 15228
rect 1821 15164 1837 15228
rect 1901 15164 1917 15228
rect 1981 15164 1997 15228
rect 2061 15164 2077 15228
rect 2141 15164 2157 15228
rect 2221 15164 2237 15228
rect 2301 15164 2317 15228
rect 2381 15164 2397 15228
rect 2461 15164 2477 15228
rect 2541 15164 2557 15228
rect 2621 15164 2637 15228
rect 2701 15164 2717 15228
rect 2781 15164 2797 15228
rect 2861 15164 2877 15228
rect 2941 15164 2957 15228
rect 3021 15164 3037 15228
rect 3101 15164 3117 15228
rect 3181 15164 3197 15228
rect 3261 15164 3277 15228
rect 3341 15164 3357 15228
rect 3421 15164 3437 15228
rect 3501 15164 3517 15228
rect 3581 15164 3597 15228
rect 3661 15164 3677 15228
rect 3741 15164 3757 15228
rect 3821 15164 3837 15228
rect 3901 15164 3917 15228
rect 3981 15164 3997 15228
rect 4061 15164 4077 15228
rect 4141 15164 4157 15228
rect 4221 15164 4237 15228
rect 4301 15164 4317 15228
rect 4381 15164 4397 15228
rect 4461 15164 4477 15228
rect 4541 15164 4557 15228
rect 4621 15164 4637 15228
rect 4701 15164 4717 15228
rect 4781 15164 4797 15228
rect 4861 15164 4900 15228
rect 0 15147 4900 15164
rect 0 15083 157 15147
rect 221 15083 237 15147
rect 301 15083 317 15147
rect 381 15083 397 15147
rect 461 15083 477 15147
rect 541 15083 557 15147
rect 621 15083 637 15147
rect 701 15083 717 15147
rect 781 15083 797 15147
rect 861 15083 877 15147
rect 941 15083 957 15147
rect 1021 15083 1037 15147
rect 1101 15083 1117 15147
rect 1181 15083 1197 15147
rect 1261 15083 1277 15147
rect 1341 15083 1357 15147
rect 1421 15083 1437 15147
rect 1501 15083 1517 15147
rect 1581 15083 1597 15147
rect 1661 15083 1677 15147
rect 1741 15083 1757 15147
rect 1821 15083 1837 15147
rect 1901 15083 1917 15147
rect 1981 15083 1997 15147
rect 2061 15083 2077 15147
rect 2141 15083 2157 15147
rect 2221 15083 2237 15147
rect 2301 15083 2317 15147
rect 2381 15083 2397 15147
rect 2461 15083 2477 15147
rect 2541 15083 2557 15147
rect 2621 15083 2637 15147
rect 2701 15083 2717 15147
rect 2781 15083 2797 15147
rect 2861 15083 2877 15147
rect 2941 15083 2957 15147
rect 3021 15083 3037 15147
rect 3101 15083 3117 15147
rect 3181 15083 3197 15147
rect 3261 15083 3277 15147
rect 3341 15083 3357 15147
rect 3421 15083 3437 15147
rect 3501 15083 3517 15147
rect 3581 15083 3597 15147
rect 3661 15083 3677 15147
rect 3741 15083 3757 15147
rect 3821 15083 3837 15147
rect 3901 15083 3917 15147
rect 3981 15083 3997 15147
rect 4061 15083 4077 15147
rect 4141 15083 4157 15147
rect 4221 15083 4237 15147
rect 4301 15083 4317 15147
rect 4381 15083 4397 15147
rect 4461 15083 4477 15147
rect 4541 15083 4557 15147
rect 4621 15083 4637 15147
rect 4701 15083 4717 15147
rect 4781 15083 4797 15147
rect 4861 15083 4900 15147
rect 0 15066 4900 15083
rect 0 15002 157 15066
rect 221 15002 237 15066
rect 301 15002 317 15066
rect 381 15002 397 15066
rect 461 15002 477 15066
rect 541 15002 557 15066
rect 621 15002 637 15066
rect 701 15002 717 15066
rect 781 15002 797 15066
rect 861 15002 877 15066
rect 941 15002 957 15066
rect 1021 15002 1037 15066
rect 1101 15002 1117 15066
rect 1181 15002 1197 15066
rect 1261 15002 1277 15066
rect 1341 15002 1357 15066
rect 1421 15002 1437 15066
rect 1501 15002 1517 15066
rect 1581 15002 1597 15066
rect 1661 15002 1677 15066
rect 1741 15002 1757 15066
rect 1821 15002 1837 15066
rect 1901 15002 1917 15066
rect 1981 15002 1997 15066
rect 2061 15002 2077 15066
rect 2141 15002 2157 15066
rect 2221 15002 2237 15066
rect 2301 15002 2317 15066
rect 2381 15002 2397 15066
rect 2461 15002 2477 15066
rect 2541 15002 2557 15066
rect 2621 15002 2637 15066
rect 2701 15002 2717 15066
rect 2781 15002 2797 15066
rect 2861 15002 2877 15066
rect 2941 15002 2957 15066
rect 3021 15002 3037 15066
rect 3101 15002 3117 15066
rect 3181 15002 3197 15066
rect 3261 15002 3277 15066
rect 3341 15002 3357 15066
rect 3421 15002 3437 15066
rect 3501 15002 3517 15066
rect 3581 15002 3597 15066
rect 3661 15002 3677 15066
rect 3741 15002 3757 15066
rect 3821 15002 3837 15066
rect 3901 15002 3917 15066
rect 3981 15002 3997 15066
rect 4061 15002 4077 15066
rect 4141 15002 4157 15066
rect 4221 15002 4237 15066
rect 4301 15002 4317 15066
rect 4381 15002 4397 15066
rect 4461 15002 4477 15066
rect 4541 15002 4557 15066
rect 4621 15002 4637 15066
rect 4701 15002 4717 15066
rect 4781 15002 4797 15066
rect 4861 15002 4900 15066
rect 0 14985 4900 15002
rect 0 14921 157 14985
rect 221 14921 237 14985
rect 301 14921 317 14985
rect 381 14921 397 14985
rect 461 14921 477 14985
rect 541 14921 557 14985
rect 621 14921 637 14985
rect 701 14921 717 14985
rect 781 14921 797 14985
rect 861 14921 877 14985
rect 941 14921 957 14985
rect 1021 14921 1037 14985
rect 1101 14921 1117 14985
rect 1181 14921 1197 14985
rect 1261 14921 1277 14985
rect 1341 14921 1357 14985
rect 1421 14921 1437 14985
rect 1501 14921 1517 14985
rect 1581 14921 1597 14985
rect 1661 14921 1677 14985
rect 1741 14921 1757 14985
rect 1821 14921 1837 14985
rect 1901 14921 1917 14985
rect 1981 14921 1997 14985
rect 2061 14921 2077 14985
rect 2141 14921 2157 14985
rect 2221 14921 2237 14985
rect 2301 14921 2317 14985
rect 2381 14921 2397 14985
rect 2461 14921 2477 14985
rect 2541 14921 2557 14985
rect 2621 14921 2637 14985
rect 2701 14921 2717 14985
rect 2781 14921 2797 14985
rect 2861 14921 2877 14985
rect 2941 14921 2957 14985
rect 3021 14921 3037 14985
rect 3101 14921 3117 14985
rect 3181 14921 3197 14985
rect 3261 14921 3277 14985
rect 3341 14921 3357 14985
rect 3421 14921 3437 14985
rect 3501 14921 3517 14985
rect 3581 14921 3597 14985
rect 3661 14921 3677 14985
rect 3741 14921 3757 14985
rect 3821 14921 3837 14985
rect 3901 14921 3917 14985
rect 3981 14921 3997 14985
rect 4061 14921 4077 14985
rect 4141 14921 4157 14985
rect 4221 14921 4237 14985
rect 4301 14921 4317 14985
rect 4381 14921 4397 14985
rect 4461 14921 4477 14985
rect 4541 14921 4557 14985
rect 4621 14921 4637 14985
rect 4701 14921 4717 14985
rect 4781 14921 4797 14985
rect 4861 14921 4900 14985
rect 0 14904 4900 14921
rect 0 14840 157 14904
rect 221 14840 237 14904
rect 301 14840 317 14904
rect 381 14840 397 14904
rect 461 14840 477 14904
rect 541 14840 557 14904
rect 621 14840 637 14904
rect 701 14840 717 14904
rect 781 14840 797 14904
rect 861 14840 877 14904
rect 941 14840 957 14904
rect 1021 14840 1037 14904
rect 1101 14840 1117 14904
rect 1181 14840 1197 14904
rect 1261 14840 1277 14904
rect 1341 14840 1357 14904
rect 1421 14840 1437 14904
rect 1501 14840 1517 14904
rect 1581 14840 1597 14904
rect 1661 14840 1677 14904
rect 1741 14840 1757 14904
rect 1821 14840 1837 14904
rect 1901 14840 1917 14904
rect 1981 14840 1997 14904
rect 2061 14840 2077 14904
rect 2141 14840 2157 14904
rect 2221 14840 2237 14904
rect 2301 14840 2317 14904
rect 2381 14840 2397 14904
rect 2461 14840 2477 14904
rect 2541 14840 2557 14904
rect 2621 14840 2637 14904
rect 2701 14840 2717 14904
rect 2781 14840 2797 14904
rect 2861 14840 2877 14904
rect 2941 14840 2957 14904
rect 3021 14840 3037 14904
rect 3101 14840 3117 14904
rect 3181 14840 3197 14904
rect 3261 14840 3277 14904
rect 3341 14840 3357 14904
rect 3421 14840 3437 14904
rect 3501 14840 3517 14904
rect 3581 14840 3597 14904
rect 3661 14840 3677 14904
rect 3741 14840 3757 14904
rect 3821 14840 3837 14904
rect 3901 14840 3917 14904
rect 3981 14840 3997 14904
rect 4061 14840 4077 14904
rect 4141 14840 4157 14904
rect 4221 14840 4237 14904
rect 4301 14840 4317 14904
rect 4381 14840 4397 14904
rect 4461 14840 4477 14904
rect 4541 14840 4557 14904
rect 4621 14840 4637 14904
rect 4701 14840 4717 14904
rect 4781 14840 4797 14904
rect 4861 14840 4900 14904
rect 0 14823 4900 14840
rect 0 14759 157 14823
rect 221 14759 237 14823
rect 301 14759 317 14823
rect 381 14759 397 14823
rect 461 14759 477 14823
rect 541 14759 557 14823
rect 621 14759 637 14823
rect 701 14759 717 14823
rect 781 14759 797 14823
rect 861 14759 877 14823
rect 941 14759 957 14823
rect 1021 14759 1037 14823
rect 1101 14759 1117 14823
rect 1181 14759 1197 14823
rect 1261 14759 1277 14823
rect 1341 14759 1357 14823
rect 1421 14759 1437 14823
rect 1501 14759 1517 14823
rect 1581 14759 1597 14823
rect 1661 14759 1677 14823
rect 1741 14759 1757 14823
rect 1821 14759 1837 14823
rect 1901 14759 1917 14823
rect 1981 14759 1997 14823
rect 2061 14759 2077 14823
rect 2141 14759 2157 14823
rect 2221 14759 2237 14823
rect 2301 14759 2317 14823
rect 2381 14759 2397 14823
rect 2461 14759 2477 14823
rect 2541 14759 2557 14823
rect 2621 14759 2637 14823
rect 2701 14759 2717 14823
rect 2781 14759 2797 14823
rect 2861 14759 2877 14823
rect 2941 14759 2957 14823
rect 3021 14759 3037 14823
rect 3101 14759 3117 14823
rect 3181 14759 3197 14823
rect 3261 14759 3277 14823
rect 3341 14759 3357 14823
rect 3421 14759 3437 14823
rect 3501 14759 3517 14823
rect 3581 14759 3597 14823
rect 3661 14759 3677 14823
rect 3741 14759 3757 14823
rect 3821 14759 3837 14823
rect 3901 14759 3917 14823
rect 3981 14759 3997 14823
rect 4061 14759 4077 14823
rect 4141 14759 4157 14823
rect 4221 14759 4237 14823
rect 4301 14759 4317 14823
rect 4381 14759 4397 14823
rect 4461 14759 4477 14823
rect 4541 14759 4557 14823
rect 4621 14759 4637 14823
rect 4701 14759 4717 14823
rect 4781 14759 4797 14823
rect 4861 14759 4900 14823
rect 0 14742 4900 14759
rect 0 14678 157 14742
rect 221 14678 237 14742
rect 301 14678 317 14742
rect 381 14678 397 14742
rect 461 14678 477 14742
rect 541 14678 557 14742
rect 621 14678 637 14742
rect 701 14678 717 14742
rect 781 14678 797 14742
rect 861 14678 877 14742
rect 941 14678 957 14742
rect 1021 14678 1037 14742
rect 1101 14678 1117 14742
rect 1181 14678 1197 14742
rect 1261 14678 1277 14742
rect 1341 14678 1357 14742
rect 1421 14678 1437 14742
rect 1501 14678 1517 14742
rect 1581 14678 1597 14742
rect 1661 14678 1677 14742
rect 1741 14678 1757 14742
rect 1821 14678 1837 14742
rect 1901 14678 1917 14742
rect 1981 14678 1997 14742
rect 2061 14678 2077 14742
rect 2141 14678 2157 14742
rect 2221 14678 2237 14742
rect 2301 14678 2317 14742
rect 2381 14678 2397 14742
rect 2461 14678 2477 14742
rect 2541 14678 2557 14742
rect 2621 14678 2637 14742
rect 2701 14678 2717 14742
rect 2781 14678 2797 14742
rect 2861 14678 2877 14742
rect 2941 14678 2957 14742
rect 3021 14678 3037 14742
rect 3101 14678 3117 14742
rect 3181 14678 3197 14742
rect 3261 14678 3277 14742
rect 3341 14678 3357 14742
rect 3421 14678 3437 14742
rect 3501 14678 3517 14742
rect 3581 14678 3597 14742
rect 3661 14678 3677 14742
rect 3741 14678 3757 14742
rect 3821 14678 3837 14742
rect 3901 14678 3917 14742
rect 3981 14678 3997 14742
rect 4061 14678 4077 14742
rect 4141 14678 4157 14742
rect 4221 14678 4237 14742
rect 4301 14678 4317 14742
rect 4381 14678 4397 14742
rect 4461 14678 4477 14742
rect 4541 14678 4557 14742
rect 4621 14678 4637 14742
rect 4701 14678 4717 14742
rect 4781 14678 4797 14742
rect 4861 14678 4900 14742
rect 0 14661 4900 14678
rect 0 14597 157 14661
rect 221 14597 237 14661
rect 301 14597 317 14661
rect 381 14597 397 14661
rect 461 14597 477 14661
rect 541 14597 557 14661
rect 621 14597 637 14661
rect 701 14597 717 14661
rect 781 14597 797 14661
rect 861 14597 877 14661
rect 941 14597 957 14661
rect 1021 14597 1037 14661
rect 1101 14597 1117 14661
rect 1181 14597 1197 14661
rect 1261 14597 1277 14661
rect 1341 14597 1357 14661
rect 1421 14597 1437 14661
rect 1501 14597 1517 14661
rect 1581 14597 1597 14661
rect 1661 14597 1677 14661
rect 1741 14597 1757 14661
rect 1821 14597 1837 14661
rect 1901 14597 1917 14661
rect 1981 14597 1997 14661
rect 2061 14597 2077 14661
rect 2141 14597 2157 14661
rect 2221 14597 2237 14661
rect 2301 14597 2317 14661
rect 2381 14597 2397 14661
rect 2461 14597 2477 14661
rect 2541 14597 2557 14661
rect 2621 14597 2637 14661
rect 2701 14597 2717 14661
rect 2781 14597 2797 14661
rect 2861 14597 2877 14661
rect 2941 14597 2957 14661
rect 3021 14597 3037 14661
rect 3101 14597 3117 14661
rect 3181 14597 3197 14661
rect 3261 14597 3277 14661
rect 3341 14597 3357 14661
rect 3421 14597 3437 14661
rect 3501 14597 3517 14661
rect 3581 14597 3597 14661
rect 3661 14597 3677 14661
rect 3741 14597 3757 14661
rect 3821 14597 3837 14661
rect 3901 14597 3917 14661
rect 3981 14597 3997 14661
rect 4061 14597 4077 14661
rect 4141 14597 4157 14661
rect 4221 14597 4237 14661
rect 4301 14597 4317 14661
rect 4381 14597 4397 14661
rect 4461 14597 4477 14661
rect 4541 14597 4557 14661
rect 4621 14597 4637 14661
rect 4701 14597 4717 14661
rect 4781 14597 4797 14661
rect 4861 14597 4900 14661
rect 0 14579 4900 14597
rect 0 14515 157 14579
rect 221 14515 237 14579
rect 301 14515 317 14579
rect 381 14515 397 14579
rect 461 14515 477 14579
rect 541 14515 557 14579
rect 621 14515 637 14579
rect 701 14515 717 14579
rect 781 14515 797 14579
rect 861 14515 877 14579
rect 941 14515 957 14579
rect 1021 14515 1037 14579
rect 1101 14515 1117 14579
rect 1181 14515 1197 14579
rect 1261 14515 1277 14579
rect 1341 14515 1357 14579
rect 1421 14515 1437 14579
rect 1501 14515 1517 14579
rect 1581 14515 1597 14579
rect 1661 14515 1677 14579
rect 1741 14515 1757 14579
rect 1821 14515 1837 14579
rect 1901 14515 1917 14579
rect 1981 14515 1997 14579
rect 2061 14515 2077 14579
rect 2141 14515 2157 14579
rect 2221 14515 2237 14579
rect 2301 14515 2317 14579
rect 2381 14515 2397 14579
rect 2461 14515 2477 14579
rect 2541 14515 2557 14579
rect 2621 14515 2637 14579
rect 2701 14515 2717 14579
rect 2781 14515 2797 14579
rect 2861 14515 2877 14579
rect 2941 14515 2957 14579
rect 3021 14515 3037 14579
rect 3101 14515 3117 14579
rect 3181 14515 3197 14579
rect 3261 14515 3277 14579
rect 3341 14515 3357 14579
rect 3421 14515 3437 14579
rect 3501 14515 3517 14579
rect 3581 14515 3597 14579
rect 3661 14515 3677 14579
rect 3741 14515 3757 14579
rect 3821 14515 3837 14579
rect 3901 14515 3917 14579
rect 3981 14515 3997 14579
rect 4061 14515 4077 14579
rect 4141 14515 4157 14579
rect 4221 14515 4237 14579
rect 4301 14515 4317 14579
rect 4381 14515 4397 14579
rect 4461 14515 4477 14579
rect 4541 14515 4557 14579
rect 4621 14515 4637 14579
rect 4701 14515 4717 14579
rect 4781 14515 4797 14579
rect 4861 14515 4900 14579
rect 0 14497 4900 14515
rect 0 14433 157 14497
rect 221 14433 237 14497
rect 301 14433 317 14497
rect 381 14433 397 14497
rect 461 14433 477 14497
rect 541 14433 557 14497
rect 621 14433 637 14497
rect 701 14433 717 14497
rect 781 14433 797 14497
rect 861 14433 877 14497
rect 941 14433 957 14497
rect 1021 14433 1037 14497
rect 1101 14433 1117 14497
rect 1181 14433 1197 14497
rect 1261 14433 1277 14497
rect 1341 14433 1357 14497
rect 1421 14433 1437 14497
rect 1501 14433 1517 14497
rect 1581 14433 1597 14497
rect 1661 14433 1677 14497
rect 1741 14433 1757 14497
rect 1821 14433 1837 14497
rect 1901 14433 1917 14497
rect 1981 14433 1997 14497
rect 2061 14433 2077 14497
rect 2141 14433 2157 14497
rect 2221 14433 2237 14497
rect 2301 14433 2317 14497
rect 2381 14433 2397 14497
rect 2461 14433 2477 14497
rect 2541 14433 2557 14497
rect 2621 14433 2637 14497
rect 2701 14433 2717 14497
rect 2781 14433 2797 14497
rect 2861 14433 2877 14497
rect 2941 14433 2957 14497
rect 3021 14433 3037 14497
rect 3101 14433 3117 14497
rect 3181 14433 3197 14497
rect 3261 14433 3277 14497
rect 3341 14433 3357 14497
rect 3421 14433 3437 14497
rect 3501 14433 3517 14497
rect 3581 14433 3597 14497
rect 3661 14433 3677 14497
rect 3741 14433 3757 14497
rect 3821 14433 3837 14497
rect 3901 14433 3917 14497
rect 3981 14433 3997 14497
rect 4061 14433 4077 14497
rect 4141 14433 4157 14497
rect 4221 14433 4237 14497
rect 4301 14433 4317 14497
rect 4381 14433 4397 14497
rect 4461 14433 4477 14497
rect 4541 14433 4557 14497
rect 4621 14433 4637 14497
rect 4701 14433 4717 14497
rect 4781 14433 4797 14497
rect 4861 14433 4900 14497
rect 0 14415 4900 14433
rect 0 14351 157 14415
rect 221 14351 237 14415
rect 301 14351 317 14415
rect 381 14351 397 14415
rect 461 14351 477 14415
rect 541 14351 557 14415
rect 621 14351 637 14415
rect 701 14351 717 14415
rect 781 14351 797 14415
rect 861 14351 877 14415
rect 941 14351 957 14415
rect 1021 14351 1037 14415
rect 1101 14351 1117 14415
rect 1181 14351 1197 14415
rect 1261 14351 1277 14415
rect 1341 14351 1357 14415
rect 1421 14351 1437 14415
rect 1501 14351 1517 14415
rect 1581 14351 1597 14415
rect 1661 14351 1677 14415
rect 1741 14351 1757 14415
rect 1821 14351 1837 14415
rect 1901 14351 1917 14415
rect 1981 14351 1997 14415
rect 2061 14351 2077 14415
rect 2141 14351 2157 14415
rect 2221 14351 2237 14415
rect 2301 14351 2317 14415
rect 2381 14351 2397 14415
rect 2461 14351 2477 14415
rect 2541 14351 2557 14415
rect 2621 14351 2637 14415
rect 2701 14351 2717 14415
rect 2781 14351 2797 14415
rect 2861 14351 2877 14415
rect 2941 14351 2957 14415
rect 3021 14351 3037 14415
rect 3101 14351 3117 14415
rect 3181 14351 3197 14415
rect 3261 14351 3277 14415
rect 3341 14351 3357 14415
rect 3421 14351 3437 14415
rect 3501 14351 3517 14415
rect 3581 14351 3597 14415
rect 3661 14351 3677 14415
rect 3741 14351 3757 14415
rect 3821 14351 3837 14415
rect 3901 14351 3917 14415
rect 3981 14351 3997 14415
rect 4061 14351 4077 14415
rect 4141 14351 4157 14415
rect 4221 14351 4237 14415
rect 4301 14351 4317 14415
rect 4381 14351 4397 14415
rect 4461 14351 4477 14415
rect 4541 14351 4557 14415
rect 4621 14351 4637 14415
rect 4701 14351 4717 14415
rect 4781 14351 4797 14415
rect 4861 14351 4900 14415
rect 0 14333 4900 14351
rect 0 14269 157 14333
rect 221 14269 237 14333
rect 301 14269 317 14333
rect 381 14269 397 14333
rect 461 14269 477 14333
rect 541 14269 557 14333
rect 621 14269 637 14333
rect 701 14269 717 14333
rect 781 14269 797 14333
rect 861 14269 877 14333
rect 941 14269 957 14333
rect 1021 14269 1037 14333
rect 1101 14269 1117 14333
rect 1181 14269 1197 14333
rect 1261 14269 1277 14333
rect 1341 14269 1357 14333
rect 1421 14269 1437 14333
rect 1501 14269 1517 14333
rect 1581 14269 1597 14333
rect 1661 14269 1677 14333
rect 1741 14269 1757 14333
rect 1821 14269 1837 14333
rect 1901 14269 1917 14333
rect 1981 14269 1997 14333
rect 2061 14269 2077 14333
rect 2141 14269 2157 14333
rect 2221 14269 2237 14333
rect 2301 14269 2317 14333
rect 2381 14269 2397 14333
rect 2461 14269 2477 14333
rect 2541 14269 2557 14333
rect 2621 14269 2637 14333
rect 2701 14269 2717 14333
rect 2781 14269 2797 14333
rect 2861 14269 2877 14333
rect 2941 14269 2957 14333
rect 3021 14269 3037 14333
rect 3101 14269 3117 14333
rect 3181 14269 3197 14333
rect 3261 14269 3277 14333
rect 3341 14269 3357 14333
rect 3421 14269 3437 14333
rect 3501 14269 3517 14333
rect 3581 14269 3597 14333
rect 3661 14269 3677 14333
rect 3741 14269 3757 14333
rect 3821 14269 3837 14333
rect 3901 14269 3917 14333
rect 3981 14269 3997 14333
rect 4061 14269 4077 14333
rect 4141 14269 4157 14333
rect 4221 14269 4237 14333
rect 4301 14269 4317 14333
rect 4381 14269 4397 14333
rect 4461 14269 4477 14333
rect 4541 14269 4557 14333
rect 4621 14269 4637 14333
rect 4701 14269 4717 14333
rect 4781 14269 4797 14333
rect 4861 14269 4900 14333
rect 0 14251 4900 14269
rect 0 14187 157 14251
rect 221 14187 237 14251
rect 301 14187 317 14251
rect 381 14187 397 14251
rect 461 14187 477 14251
rect 541 14187 557 14251
rect 621 14187 637 14251
rect 701 14187 717 14251
rect 781 14187 797 14251
rect 861 14187 877 14251
rect 941 14187 957 14251
rect 1021 14187 1037 14251
rect 1101 14187 1117 14251
rect 1181 14187 1197 14251
rect 1261 14187 1277 14251
rect 1341 14187 1357 14251
rect 1421 14187 1437 14251
rect 1501 14187 1517 14251
rect 1581 14187 1597 14251
rect 1661 14187 1677 14251
rect 1741 14187 1757 14251
rect 1821 14187 1837 14251
rect 1901 14187 1917 14251
rect 1981 14187 1997 14251
rect 2061 14187 2077 14251
rect 2141 14187 2157 14251
rect 2221 14187 2237 14251
rect 2301 14187 2317 14251
rect 2381 14187 2397 14251
rect 2461 14187 2477 14251
rect 2541 14187 2557 14251
rect 2621 14187 2637 14251
rect 2701 14187 2717 14251
rect 2781 14187 2797 14251
rect 2861 14187 2877 14251
rect 2941 14187 2957 14251
rect 3021 14187 3037 14251
rect 3101 14187 3117 14251
rect 3181 14187 3197 14251
rect 3261 14187 3277 14251
rect 3341 14187 3357 14251
rect 3421 14187 3437 14251
rect 3501 14187 3517 14251
rect 3581 14187 3597 14251
rect 3661 14187 3677 14251
rect 3741 14187 3757 14251
rect 3821 14187 3837 14251
rect 3901 14187 3917 14251
rect 3981 14187 3997 14251
rect 4061 14187 4077 14251
rect 4141 14187 4157 14251
rect 4221 14187 4237 14251
rect 4301 14187 4317 14251
rect 4381 14187 4397 14251
rect 4461 14187 4477 14251
rect 4541 14187 4557 14251
rect 4621 14187 4637 14251
rect 4701 14187 4717 14251
rect 4781 14187 4797 14251
rect 4861 14187 4900 14251
rect 0 14169 4900 14187
rect 0 14105 157 14169
rect 221 14105 237 14169
rect 301 14105 317 14169
rect 381 14105 397 14169
rect 461 14105 477 14169
rect 541 14105 557 14169
rect 621 14105 637 14169
rect 701 14105 717 14169
rect 781 14105 797 14169
rect 861 14105 877 14169
rect 941 14105 957 14169
rect 1021 14105 1037 14169
rect 1101 14105 1117 14169
rect 1181 14105 1197 14169
rect 1261 14105 1277 14169
rect 1341 14105 1357 14169
rect 1421 14105 1437 14169
rect 1501 14105 1517 14169
rect 1581 14105 1597 14169
rect 1661 14105 1677 14169
rect 1741 14105 1757 14169
rect 1821 14105 1837 14169
rect 1901 14105 1917 14169
rect 1981 14105 1997 14169
rect 2061 14105 2077 14169
rect 2141 14105 2157 14169
rect 2221 14105 2237 14169
rect 2301 14105 2317 14169
rect 2381 14105 2397 14169
rect 2461 14105 2477 14169
rect 2541 14105 2557 14169
rect 2621 14105 2637 14169
rect 2701 14105 2717 14169
rect 2781 14105 2797 14169
rect 2861 14105 2877 14169
rect 2941 14105 2957 14169
rect 3021 14105 3037 14169
rect 3101 14105 3117 14169
rect 3181 14105 3197 14169
rect 3261 14105 3277 14169
rect 3341 14105 3357 14169
rect 3421 14105 3437 14169
rect 3501 14105 3517 14169
rect 3581 14105 3597 14169
rect 3661 14105 3677 14169
rect 3741 14105 3757 14169
rect 3821 14105 3837 14169
rect 3901 14105 3917 14169
rect 3981 14105 3997 14169
rect 4061 14105 4077 14169
rect 4141 14105 4157 14169
rect 4221 14105 4237 14169
rect 4301 14105 4317 14169
rect 4381 14105 4397 14169
rect 4461 14105 4477 14169
rect 4541 14105 4557 14169
rect 4621 14105 4637 14169
rect 4701 14105 4717 14169
rect 4781 14105 4797 14169
rect 4861 14105 4900 14169
rect 0 14087 4900 14105
rect 0 14023 157 14087
rect 221 14023 237 14087
rect 301 14023 317 14087
rect 381 14023 397 14087
rect 461 14023 477 14087
rect 541 14023 557 14087
rect 621 14023 637 14087
rect 701 14023 717 14087
rect 781 14023 797 14087
rect 861 14023 877 14087
rect 941 14023 957 14087
rect 1021 14023 1037 14087
rect 1101 14023 1117 14087
rect 1181 14023 1197 14087
rect 1261 14023 1277 14087
rect 1341 14023 1357 14087
rect 1421 14023 1437 14087
rect 1501 14023 1517 14087
rect 1581 14023 1597 14087
rect 1661 14023 1677 14087
rect 1741 14023 1757 14087
rect 1821 14023 1837 14087
rect 1901 14023 1917 14087
rect 1981 14023 1997 14087
rect 2061 14023 2077 14087
rect 2141 14023 2157 14087
rect 2221 14023 2237 14087
rect 2301 14023 2317 14087
rect 2381 14023 2397 14087
rect 2461 14023 2477 14087
rect 2541 14023 2557 14087
rect 2621 14023 2637 14087
rect 2701 14023 2717 14087
rect 2781 14023 2797 14087
rect 2861 14023 2877 14087
rect 2941 14023 2957 14087
rect 3021 14023 3037 14087
rect 3101 14023 3117 14087
rect 3181 14023 3197 14087
rect 3261 14023 3277 14087
rect 3341 14023 3357 14087
rect 3421 14023 3437 14087
rect 3501 14023 3517 14087
rect 3581 14023 3597 14087
rect 3661 14023 3677 14087
rect 3741 14023 3757 14087
rect 3821 14023 3837 14087
rect 3901 14023 3917 14087
rect 3981 14023 3997 14087
rect 4061 14023 4077 14087
rect 4141 14023 4157 14087
rect 4221 14023 4237 14087
rect 4301 14023 4317 14087
rect 4381 14023 4397 14087
rect 4461 14023 4477 14087
rect 4541 14023 4557 14087
rect 4621 14023 4637 14087
rect 4701 14023 4717 14087
rect 4781 14023 4797 14087
rect 4861 14023 4900 14087
rect 0 14005 4900 14023
rect 0 13941 157 14005
rect 221 13941 237 14005
rect 301 13941 317 14005
rect 381 13941 397 14005
rect 461 13941 477 14005
rect 541 13941 557 14005
rect 621 13941 637 14005
rect 701 13941 717 14005
rect 781 13941 797 14005
rect 861 13941 877 14005
rect 941 13941 957 14005
rect 1021 13941 1037 14005
rect 1101 13941 1117 14005
rect 1181 13941 1197 14005
rect 1261 13941 1277 14005
rect 1341 13941 1357 14005
rect 1421 13941 1437 14005
rect 1501 13941 1517 14005
rect 1581 13941 1597 14005
rect 1661 13941 1677 14005
rect 1741 13941 1757 14005
rect 1821 13941 1837 14005
rect 1901 13941 1917 14005
rect 1981 13941 1997 14005
rect 2061 13941 2077 14005
rect 2141 13941 2157 14005
rect 2221 13941 2237 14005
rect 2301 13941 2317 14005
rect 2381 13941 2397 14005
rect 2461 13941 2477 14005
rect 2541 13941 2557 14005
rect 2621 13941 2637 14005
rect 2701 13941 2717 14005
rect 2781 13941 2797 14005
rect 2861 13941 2877 14005
rect 2941 13941 2957 14005
rect 3021 13941 3037 14005
rect 3101 13941 3117 14005
rect 3181 13941 3197 14005
rect 3261 13941 3277 14005
rect 3341 13941 3357 14005
rect 3421 13941 3437 14005
rect 3501 13941 3517 14005
rect 3581 13941 3597 14005
rect 3661 13941 3677 14005
rect 3741 13941 3757 14005
rect 3821 13941 3837 14005
rect 3901 13941 3917 14005
rect 3981 13941 3997 14005
rect 4061 13941 4077 14005
rect 4141 13941 4157 14005
rect 4221 13941 4237 14005
rect 4301 13941 4317 14005
rect 4381 13941 4397 14005
rect 4461 13941 4477 14005
rect 4541 13941 4557 14005
rect 4621 13941 4637 14005
rect 4701 13941 4717 14005
rect 4781 13941 4797 14005
rect 4861 13941 4900 14005
rect 0 13923 4900 13941
rect 0 13859 157 13923
rect 221 13859 237 13923
rect 301 13859 317 13923
rect 381 13859 397 13923
rect 461 13859 477 13923
rect 541 13859 557 13923
rect 621 13859 637 13923
rect 701 13859 717 13923
rect 781 13859 797 13923
rect 861 13859 877 13923
rect 941 13859 957 13923
rect 1021 13859 1037 13923
rect 1101 13859 1117 13923
rect 1181 13859 1197 13923
rect 1261 13859 1277 13923
rect 1341 13859 1357 13923
rect 1421 13859 1437 13923
rect 1501 13859 1517 13923
rect 1581 13859 1597 13923
rect 1661 13859 1677 13923
rect 1741 13859 1757 13923
rect 1821 13859 1837 13923
rect 1901 13859 1917 13923
rect 1981 13859 1997 13923
rect 2061 13859 2077 13923
rect 2141 13859 2157 13923
rect 2221 13859 2237 13923
rect 2301 13859 2317 13923
rect 2381 13859 2397 13923
rect 2461 13859 2477 13923
rect 2541 13859 2557 13923
rect 2621 13859 2637 13923
rect 2701 13859 2717 13923
rect 2781 13859 2797 13923
rect 2861 13859 2877 13923
rect 2941 13859 2957 13923
rect 3021 13859 3037 13923
rect 3101 13859 3117 13923
rect 3181 13859 3197 13923
rect 3261 13859 3277 13923
rect 3341 13859 3357 13923
rect 3421 13859 3437 13923
rect 3501 13859 3517 13923
rect 3581 13859 3597 13923
rect 3661 13859 3677 13923
rect 3741 13859 3757 13923
rect 3821 13859 3837 13923
rect 3901 13859 3917 13923
rect 3981 13859 3997 13923
rect 4061 13859 4077 13923
rect 4141 13859 4157 13923
rect 4221 13859 4237 13923
rect 4301 13859 4317 13923
rect 4381 13859 4397 13923
rect 4461 13859 4477 13923
rect 4541 13859 4557 13923
rect 4621 13859 4637 13923
rect 4701 13859 4717 13923
rect 4781 13859 4797 13923
rect 4861 13859 4900 13923
rect 0 13841 4900 13859
rect 0 13777 157 13841
rect 221 13777 237 13841
rect 301 13777 317 13841
rect 381 13777 397 13841
rect 461 13777 477 13841
rect 541 13777 557 13841
rect 621 13777 637 13841
rect 701 13777 717 13841
rect 781 13777 797 13841
rect 861 13777 877 13841
rect 941 13777 957 13841
rect 1021 13777 1037 13841
rect 1101 13777 1117 13841
rect 1181 13777 1197 13841
rect 1261 13777 1277 13841
rect 1341 13777 1357 13841
rect 1421 13777 1437 13841
rect 1501 13777 1517 13841
rect 1581 13777 1597 13841
rect 1661 13777 1677 13841
rect 1741 13777 1757 13841
rect 1821 13777 1837 13841
rect 1901 13777 1917 13841
rect 1981 13777 1997 13841
rect 2061 13777 2077 13841
rect 2141 13777 2157 13841
rect 2221 13777 2237 13841
rect 2301 13777 2317 13841
rect 2381 13777 2397 13841
rect 2461 13777 2477 13841
rect 2541 13777 2557 13841
rect 2621 13777 2637 13841
rect 2701 13777 2717 13841
rect 2781 13777 2797 13841
rect 2861 13777 2877 13841
rect 2941 13777 2957 13841
rect 3021 13777 3037 13841
rect 3101 13777 3117 13841
rect 3181 13777 3197 13841
rect 3261 13777 3277 13841
rect 3341 13777 3357 13841
rect 3421 13777 3437 13841
rect 3501 13777 3517 13841
rect 3581 13777 3597 13841
rect 3661 13777 3677 13841
rect 3741 13777 3757 13841
rect 3821 13777 3837 13841
rect 3901 13777 3917 13841
rect 3981 13777 3997 13841
rect 4061 13777 4077 13841
rect 4141 13777 4157 13841
rect 4221 13777 4237 13841
rect 4301 13777 4317 13841
rect 4381 13777 4397 13841
rect 4461 13777 4477 13841
rect 4541 13777 4557 13841
rect 4621 13777 4637 13841
rect 4701 13777 4717 13841
rect 4781 13777 4797 13841
rect 4861 13777 4900 13841
rect 0 13759 4900 13777
rect 0 13695 157 13759
rect 221 13695 237 13759
rect 301 13695 317 13759
rect 381 13695 397 13759
rect 461 13695 477 13759
rect 541 13695 557 13759
rect 621 13695 637 13759
rect 701 13695 717 13759
rect 781 13695 797 13759
rect 861 13695 877 13759
rect 941 13695 957 13759
rect 1021 13695 1037 13759
rect 1101 13695 1117 13759
rect 1181 13695 1197 13759
rect 1261 13695 1277 13759
rect 1341 13695 1357 13759
rect 1421 13695 1437 13759
rect 1501 13695 1517 13759
rect 1581 13695 1597 13759
rect 1661 13695 1677 13759
rect 1741 13695 1757 13759
rect 1821 13695 1837 13759
rect 1901 13695 1917 13759
rect 1981 13695 1997 13759
rect 2061 13695 2077 13759
rect 2141 13695 2157 13759
rect 2221 13695 2237 13759
rect 2301 13695 2317 13759
rect 2381 13695 2397 13759
rect 2461 13695 2477 13759
rect 2541 13695 2557 13759
rect 2621 13695 2637 13759
rect 2701 13695 2717 13759
rect 2781 13695 2797 13759
rect 2861 13695 2877 13759
rect 2941 13695 2957 13759
rect 3021 13695 3037 13759
rect 3101 13695 3117 13759
rect 3181 13695 3197 13759
rect 3261 13695 3277 13759
rect 3341 13695 3357 13759
rect 3421 13695 3437 13759
rect 3501 13695 3517 13759
rect 3581 13695 3597 13759
rect 3661 13695 3677 13759
rect 3741 13695 3757 13759
rect 3821 13695 3837 13759
rect 3901 13695 3917 13759
rect 3981 13695 3997 13759
rect 4061 13695 4077 13759
rect 4141 13695 4157 13759
rect 4221 13695 4237 13759
rect 4301 13695 4317 13759
rect 4381 13695 4397 13759
rect 4461 13695 4477 13759
rect 4541 13695 4557 13759
rect 4621 13695 4637 13759
rect 4701 13695 4717 13759
rect 4781 13695 4797 13759
rect 4861 13695 4900 13759
rect 0 13677 4900 13695
rect 0 13613 157 13677
rect 221 13613 237 13677
rect 301 13613 317 13677
rect 381 13613 397 13677
rect 461 13613 477 13677
rect 541 13613 557 13677
rect 621 13613 637 13677
rect 701 13613 717 13677
rect 781 13613 797 13677
rect 861 13613 877 13677
rect 941 13613 957 13677
rect 1021 13613 1037 13677
rect 1101 13613 1117 13677
rect 1181 13613 1197 13677
rect 1261 13613 1277 13677
rect 1341 13613 1357 13677
rect 1421 13613 1437 13677
rect 1501 13613 1517 13677
rect 1581 13613 1597 13677
rect 1661 13613 1677 13677
rect 1741 13613 1757 13677
rect 1821 13613 1837 13677
rect 1901 13613 1917 13677
rect 1981 13613 1997 13677
rect 2061 13613 2077 13677
rect 2141 13613 2157 13677
rect 2221 13613 2237 13677
rect 2301 13613 2317 13677
rect 2381 13613 2397 13677
rect 2461 13613 2477 13677
rect 2541 13613 2557 13677
rect 2621 13613 2637 13677
rect 2701 13613 2717 13677
rect 2781 13613 2797 13677
rect 2861 13613 2877 13677
rect 2941 13613 2957 13677
rect 3021 13613 3037 13677
rect 3101 13613 3117 13677
rect 3181 13613 3197 13677
rect 3261 13613 3277 13677
rect 3341 13613 3357 13677
rect 3421 13613 3437 13677
rect 3501 13613 3517 13677
rect 3581 13613 3597 13677
rect 3661 13613 3677 13677
rect 3741 13613 3757 13677
rect 3821 13613 3837 13677
rect 3901 13613 3917 13677
rect 3981 13613 3997 13677
rect 4061 13613 4077 13677
rect 4141 13613 4157 13677
rect 4221 13613 4237 13677
rect 4301 13613 4317 13677
rect 4381 13613 4397 13677
rect 4461 13613 4477 13677
rect 4541 13613 4557 13677
rect 4621 13613 4637 13677
rect 4701 13613 4717 13677
rect 4781 13613 4797 13677
rect 4861 13613 4900 13677
rect 0 13612 4900 13613
rect 10151 16524 15000 16525
rect 10151 16460 10190 16524
rect 10254 16460 10270 16524
rect 10334 16460 10350 16524
rect 10414 16460 10430 16524
rect 10494 16460 10510 16524
rect 10574 16460 10590 16524
rect 10654 16460 10670 16524
rect 10734 16460 10750 16524
rect 10814 16460 10830 16524
rect 10894 16460 10910 16524
rect 10974 16460 10990 16524
rect 11054 16460 11070 16524
rect 11134 16460 11150 16524
rect 11214 16460 11230 16524
rect 11294 16460 11310 16524
rect 11374 16460 11390 16524
rect 11454 16460 11470 16524
rect 11534 16460 11550 16524
rect 11614 16460 11630 16524
rect 11694 16460 11710 16524
rect 11774 16460 11790 16524
rect 11854 16460 11870 16524
rect 11934 16460 11950 16524
rect 12014 16460 12030 16524
rect 12094 16460 12110 16524
rect 12174 16460 12190 16524
rect 12254 16460 12270 16524
rect 12334 16460 12350 16524
rect 12414 16460 12430 16524
rect 12494 16460 12510 16524
rect 12574 16460 12590 16524
rect 12654 16460 12670 16524
rect 12734 16460 12750 16524
rect 12814 16460 12830 16524
rect 12894 16460 12910 16524
rect 12974 16460 12990 16524
rect 13054 16460 13070 16524
rect 13134 16460 13150 16524
rect 13214 16460 13230 16524
rect 13294 16460 13310 16524
rect 13374 16460 13390 16524
rect 13454 16460 13470 16524
rect 13534 16460 13550 16524
rect 13614 16460 13630 16524
rect 13694 16460 13710 16524
rect 13774 16460 13790 16524
rect 13854 16460 13870 16524
rect 13934 16460 13950 16524
rect 14014 16460 14030 16524
rect 14094 16460 14110 16524
rect 14174 16460 14190 16524
rect 14254 16460 14270 16524
rect 14334 16460 14350 16524
rect 14414 16460 14430 16524
rect 14494 16460 14510 16524
rect 14574 16460 14590 16524
rect 14654 16460 14670 16524
rect 14734 16460 14750 16524
rect 14814 16460 14830 16524
rect 14894 16460 15000 16524
rect 10151 16443 15000 16460
rect 10151 16379 10190 16443
rect 10254 16379 10270 16443
rect 10334 16379 10350 16443
rect 10414 16379 10430 16443
rect 10494 16379 10510 16443
rect 10574 16379 10590 16443
rect 10654 16379 10670 16443
rect 10734 16379 10750 16443
rect 10814 16379 10830 16443
rect 10894 16379 10910 16443
rect 10974 16379 10990 16443
rect 11054 16379 11070 16443
rect 11134 16379 11150 16443
rect 11214 16379 11230 16443
rect 11294 16379 11310 16443
rect 11374 16379 11390 16443
rect 11454 16379 11470 16443
rect 11534 16379 11550 16443
rect 11614 16379 11630 16443
rect 11694 16379 11710 16443
rect 11774 16379 11790 16443
rect 11854 16379 11870 16443
rect 11934 16379 11950 16443
rect 12014 16379 12030 16443
rect 12094 16379 12110 16443
rect 12174 16379 12190 16443
rect 12254 16379 12270 16443
rect 12334 16379 12350 16443
rect 12414 16379 12430 16443
rect 12494 16379 12510 16443
rect 12574 16379 12590 16443
rect 12654 16379 12670 16443
rect 12734 16379 12750 16443
rect 12814 16379 12830 16443
rect 12894 16379 12910 16443
rect 12974 16379 12990 16443
rect 13054 16379 13070 16443
rect 13134 16379 13150 16443
rect 13214 16379 13230 16443
rect 13294 16379 13310 16443
rect 13374 16379 13390 16443
rect 13454 16379 13470 16443
rect 13534 16379 13550 16443
rect 13614 16379 13630 16443
rect 13694 16379 13710 16443
rect 13774 16379 13790 16443
rect 13854 16379 13870 16443
rect 13934 16379 13950 16443
rect 14014 16379 14030 16443
rect 14094 16379 14110 16443
rect 14174 16379 14190 16443
rect 14254 16379 14270 16443
rect 14334 16379 14350 16443
rect 14414 16379 14430 16443
rect 14494 16379 14510 16443
rect 14574 16379 14590 16443
rect 14654 16379 14670 16443
rect 14734 16379 14750 16443
rect 14814 16379 14830 16443
rect 14894 16379 15000 16443
rect 10151 16362 15000 16379
rect 10151 16298 10190 16362
rect 10254 16298 10270 16362
rect 10334 16298 10350 16362
rect 10414 16298 10430 16362
rect 10494 16298 10510 16362
rect 10574 16298 10590 16362
rect 10654 16298 10670 16362
rect 10734 16298 10750 16362
rect 10814 16298 10830 16362
rect 10894 16298 10910 16362
rect 10974 16298 10990 16362
rect 11054 16298 11070 16362
rect 11134 16298 11150 16362
rect 11214 16298 11230 16362
rect 11294 16298 11310 16362
rect 11374 16298 11390 16362
rect 11454 16298 11470 16362
rect 11534 16298 11550 16362
rect 11614 16298 11630 16362
rect 11694 16298 11710 16362
rect 11774 16298 11790 16362
rect 11854 16298 11870 16362
rect 11934 16298 11950 16362
rect 12014 16298 12030 16362
rect 12094 16298 12110 16362
rect 12174 16298 12190 16362
rect 12254 16298 12270 16362
rect 12334 16298 12350 16362
rect 12414 16298 12430 16362
rect 12494 16298 12510 16362
rect 12574 16298 12590 16362
rect 12654 16298 12670 16362
rect 12734 16298 12750 16362
rect 12814 16298 12830 16362
rect 12894 16298 12910 16362
rect 12974 16298 12990 16362
rect 13054 16298 13070 16362
rect 13134 16298 13150 16362
rect 13214 16298 13230 16362
rect 13294 16298 13310 16362
rect 13374 16298 13390 16362
rect 13454 16298 13470 16362
rect 13534 16298 13550 16362
rect 13614 16298 13630 16362
rect 13694 16298 13710 16362
rect 13774 16298 13790 16362
rect 13854 16298 13870 16362
rect 13934 16298 13950 16362
rect 14014 16298 14030 16362
rect 14094 16298 14110 16362
rect 14174 16298 14190 16362
rect 14254 16298 14270 16362
rect 14334 16298 14350 16362
rect 14414 16298 14430 16362
rect 14494 16298 14510 16362
rect 14574 16298 14590 16362
rect 14654 16298 14670 16362
rect 14734 16298 14750 16362
rect 14814 16298 14830 16362
rect 14894 16298 15000 16362
rect 10151 16281 15000 16298
rect 10151 16217 10190 16281
rect 10254 16217 10270 16281
rect 10334 16217 10350 16281
rect 10414 16217 10430 16281
rect 10494 16217 10510 16281
rect 10574 16217 10590 16281
rect 10654 16217 10670 16281
rect 10734 16217 10750 16281
rect 10814 16217 10830 16281
rect 10894 16217 10910 16281
rect 10974 16217 10990 16281
rect 11054 16217 11070 16281
rect 11134 16217 11150 16281
rect 11214 16217 11230 16281
rect 11294 16217 11310 16281
rect 11374 16217 11390 16281
rect 11454 16217 11470 16281
rect 11534 16217 11550 16281
rect 11614 16217 11630 16281
rect 11694 16217 11710 16281
rect 11774 16217 11790 16281
rect 11854 16217 11870 16281
rect 11934 16217 11950 16281
rect 12014 16217 12030 16281
rect 12094 16217 12110 16281
rect 12174 16217 12190 16281
rect 12254 16217 12270 16281
rect 12334 16217 12350 16281
rect 12414 16217 12430 16281
rect 12494 16217 12510 16281
rect 12574 16217 12590 16281
rect 12654 16217 12670 16281
rect 12734 16217 12750 16281
rect 12814 16217 12830 16281
rect 12894 16217 12910 16281
rect 12974 16217 12990 16281
rect 13054 16217 13070 16281
rect 13134 16217 13150 16281
rect 13214 16217 13230 16281
rect 13294 16217 13310 16281
rect 13374 16217 13390 16281
rect 13454 16217 13470 16281
rect 13534 16217 13550 16281
rect 13614 16217 13630 16281
rect 13694 16217 13710 16281
rect 13774 16217 13790 16281
rect 13854 16217 13870 16281
rect 13934 16217 13950 16281
rect 14014 16217 14030 16281
rect 14094 16217 14110 16281
rect 14174 16217 14190 16281
rect 14254 16217 14270 16281
rect 14334 16217 14350 16281
rect 14414 16217 14430 16281
rect 14494 16217 14510 16281
rect 14574 16217 14590 16281
rect 14654 16217 14670 16281
rect 14734 16217 14750 16281
rect 14814 16217 14830 16281
rect 14894 16217 15000 16281
rect 10151 16200 15000 16217
rect 10151 16136 10190 16200
rect 10254 16136 10270 16200
rect 10334 16136 10350 16200
rect 10414 16136 10430 16200
rect 10494 16136 10510 16200
rect 10574 16136 10590 16200
rect 10654 16136 10670 16200
rect 10734 16136 10750 16200
rect 10814 16136 10830 16200
rect 10894 16136 10910 16200
rect 10974 16136 10990 16200
rect 11054 16136 11070 16200
rect 11134 16136 11150 16200
rect 11214 16136 11230 16200
rect 11294 16136 11310 16200
rect 11374 16136 11390 16200
rect 11454 16136 11470 16200
rect 11534 16136 11550 16200
rect 11614 16136 11630 16200
rect 11694 16136 11710 16200
rect 11774 16136 11790 16200
rect 11854 16136 11870 16200
rect 11934 16136 11950 16200
rect 12014 16136 12030 16200
rect 12094 16136 12110 16200
rect 12174 16136 12190 16200
rect 12254 16136 12270 16200
rect 12334 16136 12350 16200
rect 12414 16136 12430 16200
rect 12494 16136 12510 16200
rect 12574 16136 12590 16200
rect 12654 16136 12670 16200
rect 12734 16136 12750 16200
rect 12814 16136 12830 16200
rect 12894 16136 12910 16200
rect 12974 16136 12990 16200
rect 13054 16136 13070 16200
rect 13134 16136 13150 16200
rect 13214 16136 13230 16200
rect 13294 16136 13310 16200
rect 13374 16136 13390 16200
rect 13454 16136 13470 16200
rect 13534 16136 13550 16200
rect 13614 16136 13630 16200
rect 13694 16136 13710 16200
rect 13774 16136 13790 16200
rect 13854 16136 13870 16200
rect 13934 16136 13950 16200
rect 14014 16136 14030 16200
rect 14094 16136 14110 16200
rect 14174 16136 14190 16200
rect 14254 16136 14270 16200
rect 14334 16136 14350 16200
rect 14414 16136 14430 16200
rect 14494 16136 14510 16200
rect 14574 16136 14590 16200
rect 14654 16136 14670 16200
rect 14734 16136 14750 16200
rect 14814 16136 14830 16200
rect 14894 16136 15000 16200
rect 10151 16119 15000 16136
rect 10151 16055 10190 16119
rect 10254 16055 10270 16119
rect 10334 16055 10350 16119
rect 10414 16055 10430 16119
rect 10494 16055 10510 16119
rect 10574 16055 10590 16119
rect 10654 16055 10670 16119
rect 10734 16055 10750 16119
rect 10814 16055 10830 16119
rect 10894 16055 10910 16119
rect 10974 16055 10990 16119
rect 11054 16055 11070 16119
rect 11134 16055 11150 16119
rect 11214 16055 11230 16119
rect 11294 16055 11310 16119
rect 11374 16055 11390 16119
rect 11454 16055 11470 16119
rect 11534 16055 11550 16119
rect 11614 16055 11630 16119
rect 11694 16055 11710 16119
rect 11774 16055 11790 16119
rect 11854 16055 11870 16119
rect 11934 16055 11950 16119
rect 12014 16055 12030 16119
rect 12094 16055 12110 16119
rect 12174 16055 12190 16119
rect 12254 16055 12270 16119
rect 12334 16055 12350 16119
rect 12414 16055 12430 16119
rect 12494 16055 12510 16119
rect 12574 16055 12590 16119
rect 12654 16055 12670 16119
rect 12734 16055 12750 16119
rect 12814 16055 12830 16119
rect 12894 16055 12910 16119
rect 12974 16055 12990 16119
rect 13054 16055 13070 16119
rect 13134 16055 13150 16119
rect 13214 16055 13230 16119
rect 13294 16055 13310 16119
rect 13374 16055 13390 16119
rect 13454 16055 13470 16119
rect 13534 16055 13550 16119
rect 13614 16055 13630 16119
rect 13694 16055 13710 16119
rect 13774 16055 13790 16119
rect 13854 16055 13870 16119
rect 13934 16055 13950 16119
rect 14014 16055 14030 16119
rect 14094 16055 14110 16119
rect 14174 16055 14190 16119
rect 14254 16055 14270 16119
rect 14334 16055 14350 16119
rect 14414 16055 14430 16119
rect 14494 16055 14510 16119
rect 14574 16055 14590 16119
rect 14654 16055 14670 16119
rect 14734 16055 14750 16119
rect 14814 16055 14830 16119
rect 14894 16055 15000 16119
rect 10151 16038 15000 16055
rect 10151 15974 10190 16038
rect 10254 15974 10270 16038
rect 10334 15974 10350 16038
rect 10414 15974 10430 16038
rect 10494 15974 10510 16038
rect 10574 15974 10590 16038
rect 10654 15974 10670 16038
rect 10734 15974 10750 16038
rect 10814 15974 10830 16038
rect 10894 15974 10910 16038
rect 10974 15974 10990 16038
rect 11054 15974 11070 16038
rect 11134 15974 11150 16038
rect 11214 15974 11230 16038
rect 11294 15974 11310 16038
rect 11374 15974 11390 16038
rect 11454 15974 11470 16038
rect 11534 15974 11550 16038
rect 11614 15974 11630 16038
rect 11694 15974 11710 16038
rect 11774 15974 11790 16038
rect 11854 15974 11870 16038
rect 11934 15974 11950 16038
rect 12014 15974 12030 16038
rect 12094 15974 12110 16038
rect 12174 15974 12190 16038
rect 12254 15974 12270 16038
rect 12334 15974 12350 16038
rect 12414 15974 12430 16038
rect 12494 15974 12510 16038
rect 12574 15974 12590 16038
rect 12654 15974 12670 16038
rect 12734 15974 12750 16038
rect 12814 15974 12830 16038
rect 12894 15974 12910 16038
rect 12974 15974 12990 16038
rect 13054 15974 13070 16038
rect 13134 15974 13150 16038
rect 13214 15974 13230 16038
rect 13294 15974 13310 16038
rect 13374 15974 13390 16038
rect 13454 15974 13470 16038
rect 13534 15974 13550 16038
rect 13614 15974 13630 16038
rect 13694 15974 13710 16038
rect 13774 15974 13790 16038
rect 13854 15974 13870 16038
rect 13934 15974 13950 16038
rect 14014 15974 14030 16038
rect 14094 15974 14110 16038
rect 14174 15974 14190 16038
rect 14254 15974 14270 16038
rect 14334 15974 14350 16038
rect 14414 15974 14430 16038
rect 14494 15974 14510 16038
rect 14574 15974 14590 16038
rect 14654 15974 14670 16038
rect 14734 15974 14750 16038
rect 14814 15974 14830 16038
rect 14894 15974 15000 16038
rect 10151 15957 15000 15974
rect 10151 15893 10190 15957
rect 10254 15893 10270 15957
rect 10334 15893 10350 15957
rect 10414 15893 10430 15957
rect 10494 15893 10510 15957
rect 10574 15893 10590 15957
rect 10654 15893 10670 15957
rect 10734 15893 10750 15957
rect 10814 15893 10830 15957
rect 10894 15893 10910 15957
rect 10974 15893 10990 15957
rect 11054 15893 11070 15957
rect 11134 15893 11150 15957
rect 11214 15893 11230 15957
rect 11294 15893 11310 15957
rect 11374 15893 11390 15957
rect 11454 15893 11470 15957
rect 11534 15893 11550 15957
rect 11614 15893 11630 15957
rect 11694 15893 11710 15957
rect 11774 15893 11790 15957
rect 11854 15893 11870 15957
rect 11934 15893 11950 15957
rect 12014 15893 12030 15957
rect 12094 15893 12110 15957
rect 12174 15893 12190 15957
rect 12254 15893 12270 15957
rect 12334 15893 12350 15957
rect 12414 15893 12430 15957
rect 12494 15893 12510 15957
rect 12574 15893 12590 15957
rect 12654 15893 12670 15957
rect 12734 15893 12750 15957
rect 12814 15893 12830 15957
rect 12894 15893 12910 15957
rect 12974 15893 12990 15957
rect 13054 15893 13070 15957
rect 13134 15893 13150 15957
rect 13214 15893 13230 15957
rect 13294 15893 13310 15957
rect 13374 15893 13390 15957
rect 13454 15893 13470 15957
rect 13534 15893 13550 15957
rect 13614 15893 13630 15957
rect 13694 15893 13710 15957
rect 13774 15893 13790 15957
rect 13854 15893 13870 15957
rect 13934 15893 13950 15957
rect 14014 15893 14030 15957
rect 14094 15893 14110 15957
rect 14174 15893 14190 15957
rect 14254 15893 14270 15957
rect 14334 15893 14350 15957
rect 14414 15893 14430 15957
rect 14494 15893 14510 15957
rect 14574 15893 14590 15957
rect 14654 15893 14670 15957
rect 14734 15893 14750 15957
rect 14814 15893 14830 15957
rect 14894 15893 15000 15957
rect 10151 15876 15000 15893
rect 10151 15812 10190 15876
rect 10254 15812 10270 15876
rect 10334 15812 10350 15876
rect 10414 15812 10430 15876
rect 10494 15812 10510 15876
rect 10574 15812 10590 15876
rect 10654 15812 10670 15876
rect 10734 15812 10750 15876
rect 10814 15812 10830 15876
rect 10894 15812 10910 15876
rect 10974 15812 10990 15876
rect 11054 15812 11070 15876
rect 11134 15812 11150 15876
rect 11214 15812 11230 15876
rect 11294 15812 11310 15876
rect 11374 15812 11390 15876
rect 11454 15812 11470 15876
rect 11534 15812 11550 15876
rect 11614 15812 11630 15876
rect 11694 15812 11710 15876
rect 11774 15812 11790 15876
rect 11854 15812 11870 15876
rect 11934 15812 11950 15876
rect 12014 15812 12030 15876
rect 12094 15812 12110 15876
rect 12174 15812 12190 15876
rect 12254 15812 12270 15876
rect 12334 15812 12350 15876
rect 12414 15812 12430 15876
rect 12494 15812 12510 15876
rect 12574 15812 12590 15876
rect 12654 15812 12670 15876
rect 12734 15812 12750 15876
rect 12814 15812 12830 15876
rect 12894 15812 12910 15876
rect 12974 15812 12990 15876
rect 13054 15812 13070 15876
rect 13134 15812 13150 15876
rect 13214 15812 13230 15876
rect 13294 15812 13310 15876
rect 13374 15812 13390 15876
rect 13454 15812 13470 15876
rect 13534 15812 13550 15876
rect 13614 15812 13630 15876
rect 13694 15812 13710 15876
rect 13774 15812 13790 15876
rect 13854 15812 13870 15876
rect 13934 15812 13950 15876
rect 14014 15812 14030 15876
rect 14094 15812 14110 15876
rect 14174 15812 14190 15876
rect 14254 15812 14270 15876
rect 14334 15812 14350 15876
rect 14414 15812 14430 15876
rect 14494 15812 14510 15876
rect 14574 15812 14590 15876
rect 14654 15812 14670 15876
rect 14734 15812 14750 15876
rect 14814 15812 14830 15876
rect 14894 15812 15000 15876
rect 10151 15795 15000 15812
rect 10151 15731 10190 15795
rect 10254 15731 10270 15795
rect 10334 15731 10350 15795
rect 10414 15731 10430 15795
rect 10494 15731 10510 15795
rect 10574 15731 10590 15795
rect 10654 15731 10670 15795
rect 10734 15731 10750 15795
rect 10814 15731 10830 15795
rect 10894 15731 10910 15795
rect 10974 15731 10990 15795
rect 11054 15731 11070 15795
rect 11134 15731 11150 15795
rect 11214 15731 11230 15795
rect 11294 15731 11310 15795
rect 11374 15731 11390 15795
rect 11454 15731 11470 15795
rect 11534 15731 11550 15795
rect 11614 15731 11630 15795
rect 11694 15731 11710 15795
rect 11774 15731 11790 15795
rect 11854 15731 11870 15795
rect 11934 15731 11950 15795
rect 12014 15731 12030 15795
rect 12094 15731 12110 15795
rect 12174 15731 12190 15795
rect 12254 15731 12270 15795
rect 12334 15731 12350 15795
rect 12414 15731 12430 15795
rect 12494 15731 12510 15795
rect 12574 15731 12590 15795
rect 12654 15731 12670 15795
rect 12734 15731 12750 15795
rect 12814 15731 12830 15795
rect 12894 15731 12910 15795
rect 12974 15731 12990 15795
rect 13054 15731 13070 15795
rect 13134 15731 13150 15795
rect 13214 15731 13230 15795
rect 13294 15731 13310 15795
rect 13374 15731 13390 15795
rect 13454 15731 13470 15795
rect 13534 15731 13550 15795
rect 13614 15731 13630 15795
rect 13694 15731 13710 15795
rect 13774 15731 13790 15795
rect 13854 15731 13870 15795
rect 13934 15731 13950 15795
rect 14014 15731 14030 15795
rect 14094 15731 14110 15795
rect 14174 15731 14190 15795
rect 14254 15731 14270 15795
rect 14334 15731 14350 15795
rect 14414 15731 14430 15795
rect 14494 15731 14510 15795
rect 14574 15731 14590 15795
rect 14654 15731 14670 15795
rect 14734 15731 14750 15795
rect 14814 15731 14830 15795
rect 14894 15731 15000 15795
rect 10151 15714 15000 15731
rect 10151 15650 10190 15714
rect 10254 15650 10270 15714
rect 10334 15650 10350 15714
rect 10414 15650 10430 15714
rect 10494 15650 10510 15714
rect 10574 15650 10590 15714
rect 10654 15650 10670 15714
rect 10734 15650 10750 15714
rect 10814 15650 10830 15714
rect 10894 15650 10910 15714
rect 10974 15650 10990 15714
rect 11054 15650 11070 15714
rect 11134 15650 11150 15714
rect 11214 15650 11230 15714
rect 11294 15650 11310 15714
rect 11374 15650 11390 15714
rect 11454 15650 11470 15714
rect 11534 15650 11550 15714
rect 11614 15650 11630 15714
rect 11694 15650 11710 15714
rect 11774 15650 11790 15714
rect 11854 15650 11870 15714
rect 11934 15650 11950 15714
rect 12014 15650 12030 15714
rect 12094 15650 12110 15714
rect 12174 15650 12190 15714
rect 12254 15650 12270 15714
rect 12334 15650 12350 15714
rect 12414 15650 12430 15714
rect 12494 15650 12510 15714
rect 12574 15650 12590 15714
rect 12654 15650 12670 15714
rect 12734 15650 12750 15714
rect 12814 15650 12830 15714
rect 12894 15650 12910 15714
rect 12974 15650 12990 15714
rect 13054 15650 13070 15714
rect 13134 15650 13150 15714
rect 13214 15650 13230 15714
rect 13294 15650 13310 15714
rect 13374 15650 13390 15714
rect 13454 15650 13470 15714
rect 13534 15650 13550 15714
rect 13614 15650 13630 15714
rect 13694 15650 13710 15714
rect 13774 15650 13790 15714
rect 13854 15650 13870 15714
rect 13934 15650 13950 15714
rect 14014 15650 14030 15714
rect 14094 15650 14110 15714
rect 14174 15650 14190 15714
rect 14254 15650 14270 15714
rect 14334 15650 14350 15714
rect 14414 15650 14430 15714
rect 14494 15650 14510 15714
rect 14574 15650 14590 15714
rect 14654 15650 14670 15714
rect 14734 15650 14750 15714
rect 14814 15650 14830 15714
rect 14894 15650 15000 15714
rect 10151 15633 15000 15650
rect 10151 15569 10190 15633
rect 10254 15569 10270 15633
rect 10334 15569 10350 15633
rect 10414 15569 10430 15633
rect 10494 15569 10510 15633
rect 10574 15569 10590 15633
rect 10654 15569 10670 15633
rect 10734 15569 10750 15633
rect 10814 15569 10830 15633
rect 10894 15569 10910 15633
rect 10974 15569 10990 15633
rect 11054 15569 11070 15633
rect 11134 15569 11150 15633
rect 11214 15569 11230 15633
rect 11294 15569 11310 15633
rect 11374 15569 11390 15633
rect 11454 15569 11470 15633
rect 11534 15569 11550 15633
rect 11614 15569 11630 15633
rect 11694 15569 11710 15633
rect 11774 15569 11790 15633
rect 11854 15569 11870 15633
rect 11934 15569 11950 15633
rect 12014 15569 12030 15633
rect 12094 15569 12110 15633
rect 12174 15569 12190 15633
rect 12254 15569 12270 15633
rect 12334 15569 12350 15633
rect 12414 15569 12430 15633
rect 12494 15569 12510 15633
rect 12574 15569 12590 15633
rect 12654 15569 12670 15633
rect 12734 15569 12750 15633
rect 12814 15569 12830 15633
rect 12894 15569 12910 15633
rect 12974 15569 12990 15633
rect 13054 15569 13070 15633
rect 13134 15569 13150 15633
rect 13214 15569 13230 15633
rect 13294 15569 13310 15633
rect 13374 15569 13390 15633
rect 13454 15569 13470 15633
rect 13534 15569 13550 15633
rect 13614 15569 13630 15633
rect 13694 15569 13710 15633
rect 13774 15569 13790 15633
rect 13854 15569 13870 15633
rect 13934 15569 13950 15633
rect 14014 15569 14030 15633
rect 14094 15569 14110 15633
rect 14174 15569 14190 15633
rect 14254 15569 14270 15633
rect 14334 15569 14350 15633
rect 14414 15569 14430 15633
rect 14494 15569 14510 15633
rect 14574 15569 14590 15633
rect 14654 15569 14670 15633
rect 14734 15569 14750 15633
rect 14814 15569 14830 15633
rect 14894 15569 15000 15633
rect 10151 15552 15000 15569
rect 10151 15488 10190 15552
rect 10254 15488 10270 15552
rect 10334 15488 10350 15552
rect 10414 15488 10430 15552
rect 10494 15488 10510 15552
rect 10574 15488 10590 15552
rect 10654 15488 10670 15552
rect 10734 15488 10750 15552
rect 10814 15488 10830 15552
rect 10894 15488 10910 15552
rect 10974 15488 10990 15552
rect 11054 15488 11070 15552
rect 11134 15488 11150 15552
rect 11214 15488 11230 15552
rect 11294 15488 11310 15552
rect 11374 15488 11390 15552
rect 11454 15488 11470 15552
rect 11534 15488 11550 15552
rect 11614 15488 11630 15552
rect 11694 15488 11710 15552
rect 11774 15488 11790 15552
rect 11854 15488 11870 15552
rect 11934 15488 11950 15552
rect 12014 15488 12030 15552
rect 12094 15488 12110 15552
rect 12174 15488 12190 15552
rect 12254 15488 12270 15552
rect 12334 15488 12350 15552
rect 12414 15488 12430 15552
rect 12494 15488 12510 15552
rect 12574 15488 12590 15552
rect 12654 15488 12670 15552
rect 12734 15488 12750 15552
rect 12814 15488 12830 15552
rect 12894 15488 12910 15552
rect 12974 15488 12990 15552
rect 13054 15488 13070 15552
rect 13134 15488 13150 15552
rect 13214 15488 13230 15552
rect 13294 15488 13310 15552
rect 13374 15488 13390 15552
rect 13454 15488 13470 15552
rect 13534 15488 13550 15552
rect 13614 15488 13630 15552
rect 13694 15488 13710 15552
rect 13774 15488 13790 15552
rect 13854 15488 13870 15552
rect 13934 15488 13950 15552
rect 14014 15488 14030 15552
rect 14094 15488 14110 15552
rect 14174 15488 14190 15552
rect 14254 15488 14270 15552
rect 14334 15488 14350 15552
rect 14414 15488 14430 15552
rect 14494 15488 14510 15552
rect 14574 15488 14590 15552
rect 14654 15488 14670 15552
rect 14734 15488 14750 15552
rect 14814 15488 14830 15552
rect 14894 15488 15000 15552
rect 10151 15471 15000 15488
rect 10151 15407 10190 15471
rect 10254 15407 10270 15471
rect 10334 15407 10350 15471
rect 10414 15407 10430 15471
rect 10494 15407 10510 15471
rect 10574 15407 10590 15471
rect 10654 15407 10670 15471
rect 10734 15407 10750 15471
rect 10814 15407 10830 15471
rect 10894 15407 10910 15471
rect 10974 15407 10990 15471
rect 11054 15407 11070 15471
rect 11134 15407 11150 15471
rect 11214 15407 11230 15471
rect 11294 15407 11310 15471
rect 11374 15407 11390 15471
rect 11454 15407 11470 15471
rect 11534 15407 11550 15471
rect 11614 15407 11630 15471
rect 11694 15407 11710 15471
rect 11774 15407 11790 15471
rect 11854 15407 11870 15471
rect 11934 15407 11950 15471
rect 12014 15407 12030 15471
rect 12094 15407 12110 15471
rect 12174 15407 12190 15471
rect 12254 15407 12270 15471
rect 12334 15407 12350 15471
rect 12414 15407 12430 15471
rect 12494 15407 12510 15471
rect 12574 15407 12590 15471
rect 12654 15407 12670 15471
rect 12734 15407 12750 15471
rect 12814 15407 12830 15471
rect 12894 15407 12910 15471
rect 12974 15407 12990 15471
rect 13054 15407 13070 15471
rect 13134 15407 13150 15471
rect 13214 15407 13230 15471
rect 13294 15407 13310 15471
rect 13374 15407 13390 15471
rect 13454 15407 13470 15471
rect 13534 15407 13550 15471
rect 13614 15407 13630 15471
rect 13694 15407 13710 15471
rect 13774 15407 13790 15471
rect 13854 15407 13870 15471
rect 13934 15407 13950 15471
rect 14014 15407 14030 15471
rect 14094 15407 14110 15471
rect 14174 15407 14190 15471
rect 14254 15407 14270 15471
rect 14334 15407 14350 15471
rect 14414 15407 14430 15471
rect 14494 15407 14510 15471
rect 14574 15407 14590 15471
rect 14654 15407 14670 15471
rect 14734 15407 14750 15471
rect 14814 15407 14830 15471
rect 14894 15407 15000 15471
rect 10151 15390 15000 15407
rect 10151 15326 10190 15390
rect 10254 15326 10270 15390
rect 10334 15326 10350 15390
rect 10414 15326 10430 15390
rect 10494 15326 10510 15390
rect 10574 15326 10590 15390
rect 10654 15326 10670 15390
rect 10734 15326 10750 15390
rect 10814 15326 10830 15390
rect 10894 15326 10910 15390
rect 10974 15326 10990 15390
rect 11054 15326 11070 15390
rect 11134 15326 11150 15390
rect 11214 15326 11230 15390
rect 11294 15326 11310 15390
rect 11374 15326 11390 15390
rect 11454 15326 11470 15390
rect 11534 15326 11550 15390
rect 11614 15326 11630 15390
rect 11694 15326 11710 15390
rect 11774 15326 11790 15390
rect 11854 15326 11870 15390
rect 11934 15326 11950 15390
rect 12014 15326 12030 15390
rect 12094 15326 12110 15390
rect 12174 15326 12190 15390
rect 12254 15326 12270 15390
rect 12334 15326 12350 15390
rect 12414 15326 12430 15390
rect 12494 15326 12510 15390
rect 12574 15326 12590 15390
rect 12654 15326 12670 15390
rect 12734 15326 12750 15390
rect 12814 15326 12830 15390
rect 12894 15326 12910 15390
rect 12974 15326 12990 15390
rect 13054 15326 13070 15390
rect 13134 15326 13150 15390
rect 13214 15326 13230 15390
rect 13294 15326 13310 15390
rect 13374 15326 13390 15390
rect 13454 15326 13470 15390
rect 13534 15326 13550 15390
rect 13614 15326 13630 15390
rect 13694 15326 13710 15390
rect 13774 15326 13790 15390
rect 13854 15326 13870 15390
rect 13934 15326 13950 15390
rect 14014 15326 14030 15390
rect 14094 15326 14110 15390
rect 14174 15326 14190 15390
rect 14254 15326 14270 15390
rect 14334 15326 14350 15390
rect 14414 15326 14430 15390
rect 14494 15326 14510 15390
rect 14574 15326 14590 15390
rect 14654 15326 14670 15390
rect 14734 15326 14750 15390
rect 14814 15326 14830 15390
rect 14894 15326 15000 15390
rect 10151 15309 15000 15326
rect 10151 15245 10190 15309
rect 10254 15245 10270 15309
rect 10334 15245 10350 15309
rect 10414 15245 10430 15309
rect 10494 15245 10510 15309
rect 10574 15245 10590 15309
rect 10654 15245 10670 15309
rect 10734 15245 10750 15309
rect 10814 15245 10830 15309
rect 10894 15245 10910 15309
rect 10974 15245 10990 15309
rect 11054 15245 11070 15309
rect 11134 15245 11150 15309
rect 11214 15245 11230 15309
rect 11294 15245 11310 15309
rect 11374 15245 11390 15309
rect 11454 15245 11470 15309
rect 11534 15245 11550 15309
rect 11614 15245 11630 15309
rect 11694 15245 11710 15309
rect 11774 15245 11790 15309
rect 11854 15245 11870 15309
rect 11934 15245 11950 15309
rect 12014 15245 12030 15309
rect 12094 15245 12110 15309
rect 12174 15245 12190 15309
rect 12254 15245 12270 15309
rect 12334 15245 12350 15309
rect 12414 15245 12430 15309
rect 12494 15245 12510 15309
rect 12574 15245 12590 15309
rect 12654 15245 12670 15309
rect 12734 15245 12750 15309
rect 12814 15245 12830 15309
rect 12894 15245 12910 15309
rect 12974 15245 12990 15309
rect 13054 15245 13070 15309
rect 13134 15245 13150 15309
rect 13214 15245 13230 15309
rect 13294 15245 13310 15309
rect 13374 15245 13390 15309
rect 13454 15245 13470 15309
rect 13534 15245 13550 15309
rect 13614 15245 13630 15309
rect 13694 15245 13710 15309
rect 13774 15245 13790 15309
rect 13854 15245 13870 15309
rect 13934 15245 13950 15309
rect 14014 15245 14030 15309
rect 14094 15245 14110 15309
rect 14174 15245 14190 15309
rect 14254 15245 14270 15309
rect 14334 15245 14350 15309
rect 14414 15245 14430 15309
rect 14494 15245 14510 15309
rect 14574 15245 14590 15309
rect 14654 15245 14670 15309
rect 14734 15245 14750 15309
rect 14814 15245 14830 15309
rect 14894 15245 15000 15309
rect 10151 15228 15000 15245
rect 10151 15164 10190 15228
rect 10254 15164 10270 15228
rect 10334 15164 10350 15228
rect 10414 15164 10430 15228
rect 10494 15164 10510 15228
rect 10574 15164 10590 15228
rect 10654 15164 10670 15228
rect 10734 15164 10750 15228
rect 10814 15164 10830 15228
rect 10894 15164 10910 15228
rect 10974 15164 10990 15228
rect 11054 15164 11070 15228
rect 11134 15164 11150 15228
rect 11214 15164 11230 15228
rect 11294 15164 11310 15228
rect 11374 15164 11390 15228
rect 11454 15164 11470 15228
rect 11534 15164 11550 15228
rect 11614 15164 11630 15228
rect 11694 15164 11710 15228
rect 11774 15164 11790 15228
rect 11854 15164 11870 15228
rect 11934 15164 11950 15228
rect 12014 15164 12030 15228
rect 12094 15164 12110 15228
rect 12174 15164 12190 15228
rect 12254 15164 12270 15228
rect 12334 15164 12350 15228
rect 12414 15164 12430 15228
rect 12494 15164 12510 15228
rect 12574 15164 12590 15228
rect 12654 15164 12670 15228
rect 12734 15164 12750 15228
rect 12814 15164 12830 15228
rect 12894 15164 12910 15228
rect 12974 15164 12990 15228
rect 13054 15164 13070 15228
rect 13134 15164 13150 15228
rect 13214 15164 13230 15228
rect 13294 15164 13310 15228
rect 13374 15164 13390 15228
rect 13454 15164 13470 15228
rect 13534 15164 13550 15228
rect 13614 15164 13630 15228
rect 13694 15164 13710 15228
rect 13774 15164 13790 15228
rect 13854 15164 13870 15228
rect 13934 15164 13950 15228
rect 14014 15164 14030 15228
rect 14094 15164 14110 15228
rect 14174 15164 14190 15228
rect 14254 15164 14270 15228
rect 14334 15164 14350 15228
rect 14414 15164 14430 15228
rect 14494 15164 14510 15228
rect 14574 15164 14590 15228
rect 14654 15164 14670 15228
rect 14734 15164 14750 15228
rect 14814 15164 14830 15228
rect 14894 15164 15000 15228
rect 10151 15147 15000 15164
rect 10151 15083 10190 15147
rect 10254 15083 10270 15147
rect 10334 15083 10350 15147
rect 10414 15083 10430 15147
rect 10494 15083 10510 15147
rect 10574 15083 10590 15147
rect 10654 15083 10670 15147
rect 10734 15083 10750 15147
rect 10814 15083 10830 15147
rect 10894 15083 10910 15147
rect 10974 15083 10990 15147
rect 11054 15083 11070 15147
rect 11134 15083 11150 15147
rect 11214 15083 11230 15147
rect 11294 15083 11310 15147
rect 11374 15083 11390 15147
rect 11454 15083 11470 15147
rect 11534 15083 11550 15147
rect 11614 15083 11630 15147
rect 11694 15083 11710 15147
rect 11774 15083 11790 15147
rect 11854 15083 11870 15147
rect 11934 15083 11950 15147
rect 12014 15083 12030 15147
rect 12094 15083 12110 15147
rect 12174 15083 12190 15147
rect 12254 15083 12270 15147
rect 12334 15083 12350 15147
rect 12414 15083 12430 15147
rect 12494 15083 12510 15147
rect 12574 15083 12590 15147
rect 12654 15083 12670 15147
rect 12734 15083 12750 15147
rect 12814 15083 12830 15147
rect 12894 15083 12910 15147
rect 12974 15083 12990 15147
rect 13054 15083 13070 15147
rect 13134 15083 13150 15147
rect 13214 15083 13230 15147
rect 13294 15083 13310 15147
rect 13374 15083 13390 15147
rect 13454 15083 13470 15147
rect 13534 15083 13550 15147
rect 13614 15083 13630 15147
rect 13694 15083 13710 15147
rect 13774 15083 13790 15147
rect 13854 15083 13870 15147
rect 13934 15083 13950 15147
rect 14014 15083 14030 15147
rect 14094 15083 14110 15147
rect 14174 15083 14190 15147
rect 14254 15083 14270 15147
rect 14334 15083 14350 15147
rect 14414 15083 14430 15147
rect 14494 15083 14510 15147
rect 14574 15083 14590 15147
rect 14654 15083 14670 15147
rect 14734 15083 14750 15147
rect 14814 15083 14830 15147
rect 14894 15083 15000 15147
rect 10151 15066 15000 15083
rect 10151 15002 10190 15066
rect 10254 15002 10270 15066
rect 10334 15002 10350 15066
rect 10414 15002 10430 15066
rect 10494 15002 10510 15066
rect 10574 15002 10590 15066
rect 10654 15002 10670 15066
rect 10734 15002 10750 15066
rect 10814 15002 10830 15066
rect 10894 15002 10910 15066
rect 10974 15002 10990 15066
rect 11054 15002 11070 15066
rect 11134 15002 11150 15066
rect 11214 15002 11230 15066
rect 11294 15002 11310 15066
rect 11374 15002 11390 15066
rect 11454 15002 11470 15066
rect 11534 15002 11550 15066
rect 11614 15002 11630 15066
rect 11694 15002 11710 15066
rect 11774 15002 11790 15066
rect 11854 15002 11870 15066
rect 11934 15002 11950 15066
rect 12014 15002 12030 15066
rect 12094 15002 12110 15066
rect 12174 15002 12190 15066
rect 12254 15002 12270 15066
rect 12334 15002 12350 15066
rect 12414 15002 12430 15066
rect 12494 15002 12510 15066
rect 12574 15002 12590 15066
rect 12654 15002 12670 15066
rect 12734 15002 12750 15066
rect 12814 15002 12830 15066
rect 12894 15002 12910 15066
rect 12974 15002 12990 15066
rect 13054 15002 13070 15066
rect 13134 15002 13150 15066
rect 13214 15002 13230 15066
rect 13294 15002 13310 15066
rect 13374 15002 13390 15066
rect 13454 15002 13470 15066
rect 13534 15002 13550 15066
rect 13614 15002 13630 15066
rect 13694 15002 13710 15066
rect 13774 15002 13790 15066
rect 13854 15002 13870 15066
rect 13934 15002 13950 15066
rect 14014 15002 14030 15066
rect 14094 15002 14110 15066
rect 14174 15002 14190 15066
rect 14254 15002 14270 15066
rect 14334 15002 14350 15066
rect 14414 15002 14430 15066
rect 14494 15002 14510 15066
rect 14574 15002 14590 15066
rect 14654 15002 14670 15066
rect 14734 15002 14750 15066
rect 14814 15002 14830 15066
rect 14894 15002 15000 15066
rect 10151 14985 15000 15002
rect 10151 14921 10190 14985
rect 10254 14921 10270 14985
rect 10334 14921 10350 14985
rect 10414 14921 10430 14985
rect 10494 14921 10510 14985
rect 10574 14921 10590 14985
rect 10654 14921 10670 14985
rect 10734 14921 10750 14985
rect 10814 14921 10830 14985
rect 10894 14921 10910 14985
rect 10974 14921 10990 14985
rect 11054 14921 11070 14985
rect 11134 14921 11150 14985
rect 11214 14921 11230 14985
rect 11294 14921 11310 14985
rect 11374 14921 11390 14985
rect 11454 14921 11470 14985
rect 11534 14921 11550 14985
rect 11614 14921 11630 14985
rect 11694 14921 11710 14985
rect 11774 14921 11790 14985
rect 11854 14921 11870 14985
rect 11934 14921 11950 14985
rect 12014 14921 12030 14985
rect 12094 14921 12110 14985
rect 12174 14921 12190 14985
rect 12254 14921 12270 14985
rect 12334 14921 12350 14985
rect 12414 14921 12430 14985
rect 12494 14921 12510 14985
rect 12574 14921 12590 14985
rect 12654 14921 12670 14985
rect 12734 14921 12750 14985
rect 12814 14921 12830 14985
rect 12894 14921 12910 14985
rect 12974 14921 12990 14985
rect 13054 14921 13070 14985
rect 13134 14921 13150 14985
rect 13214 14921 13230 14985
rect 13294 14921 13310 14985
rect 13374 14921 13390 14985
rect 13454 14921 13470 14985
rect 13534 14921 13550 14985
rect 13614 14921 13630 14985
rect 13694 14921 13710 14985
rect 13774 14921 13790 14985
rect 13854 14921 13870 14985
rect 13934 14921 13950 14985
rect 14014 14921 14030 14985
rect 14094 14921 14110 14985
rect 14174 14921 14190 14985
rect 14254 14921 14270 14985
rect 14334 14921 14350 14985
rect 14414 14921 14430 14985
rect 14494 14921 14510 14985
rect 14574 14921 14590 14985
rect 14654 14921 14670 14985
rect 14734 14921 14750 14985
rect 14814 14921 14830 14985
rect 14894 14921 15000 14985
rect 10151 14904 15000 14921
rect 10151 14840 10190 14904
rect 10254 14840 10270 14904
rect 10334 14840 10350 14904
rect 10414 14840 10430 14904
rect 10494 14840 10510 14904
rect 10574 14840 10590 14904
rect 10654 14840 10670 14904
rect 10734 14840 10750 14904
rect 10814 14840 10830 14904
rect 10894 14840 10910 14904
rect 10974 14840 10990 14904
rect 11054 14840 11070 14904
rect 11134 14840 11150 14904
rect 11214 14840 11230 14904
rect 11294 14840 11310 14904
rect 11374 14840 11390 14904
rect 11454 14840 11470 14904
rect 11534 14840 11550 14904
rect 11614 14840 11630 14904
rect 11694 14840 11710 14904
rect 11774 14840 11790 14904
rect 11854 14840 11870 14904
rect 11934 14840 11950 14904
rect 12014 14840 12030 14904
rect 12094 14840 12110 14904
rect 12174 14840 12190 14904
rect 12254 14840 12270 14904
rect 12334 14840 12350 14904
rect 12414 14840 12430 14904
rect 12494 14840 12510 14904
rect 12574 14840 12590 14904
rect 12654 14840 12670 14904
rect 12734 14840 12750 14904
rect 12814 14840 12830 14904
rect 12894 14840 12910 14904
rect 12974 14840 12990 14904
rect 13054 14840 13070 14904
rect 13134 14840 13150 14904
rect 13214 14840 13230 14904
rect 13294 14840 13310 14904
rect 13374 14840 13390 14904
rect 13454 14840 13470 14904
rect 13534 14840 13550 14904
rect 13614 14840 13630 14904
rect 13694 14840 13710 14904
rect 13774 14840 13790 14904
rect 13854 14840 13870 14904
rect 13934 14840 13950 14904
rect 14014 14840 14030 14904
rect 14094 14840 14110 14904
rect 14174 14840 14190 14904
rect 14254 14840 14270 14904
rect 14334 14840 14350 14904
rect 14414 14840 14430 14904
rect 14494 14840 14510 14904
rect 14574 14840 14590 14904
rect 14654 14840 14670 14904
rect 14734 14840 14750 14904
rect 14814 14840 14830 14904
rect 14894 14840 15000 14904
rect 10151 14823 15000 14840
rect 10151 14759 10190 14823
rect 10254 14759 10270 14823
rect 10334 14759 10350 14823
rect 10414 14759 10430 14823
rect 10494 14759 10510 14823
rect 10574 14759 10590 14823
rect 10654 14759 10670 14823
rect 10734 14759 10750 14823
rect 10814 14759 10830 14823
rect 10894 14759 10910 14823
rect 10974 14759 10990 14823
rect 11054 14759 11070 14823
rect 11134 14759 11150 14823
rect 11214 14759 11230 14823
rect 11294 14759 11310 14823
rect 11374 14759 11390 14823
rect 11454 14759 11470 14823
rect 11534 14759 11550 14823
rect 11614 14759 11630 14823
rect 11694 14759 11710 14823
rect 11774 14759 11790 14823
rect 11854 14759 11870 14823
rect 11934 14759 11950 14823
rect 12014 14759 12030 14823
rect 12094 14759 12110 14823
rect 12174 14759 12190 14823
rect 12254 14759 12270 14823
rect 12334 14759 12350 14823
rect 12414 14759 12430 14823
rect 12494 14759 12510 14823
rect 12574 14759 12590 14823
rect 12654 14759 12670 14823
rect 12734 14759 12750 14823
rect 12814 14759 12830 14823
rect 12894 14759 12910 14823
rect 12974 14759 12990 14823
rect 13054 14759 13070 14823
rect 13134 14759 13150 14823
rect 13214 14759 13230 14823
rect 13294 14759 13310 14823
rect 13374 14759 13390 14823
rect 13454 14759 13470 14823
rect 13534 14759 13550 14823
rect 13614 14759 13630 14823
rect 13694 14759 13710 14823
rect 13774 14759 13790 14823
rect 13854 14759 13870 14823
rect 13934 14759 13950 14823
rect 14014 14759 14030 14823
rect 14094 14759 14110 14823
rect 14174 14759 14190 14823
rect 14254 14759 14270 14823
rect 14334 14759 14350 14823
rect 14414 14759 14430 14823
rect 14494 14759 14510 14823
rect 14574 14759 14590 14823
rect 14654 14759 14670 14823
rect 14734 14759 14750 14823
rect 14814 14759 14830 14823
rect 14894 14759 15000 14823
rect 10151 14742 15000 14759
rect 10151 14678 10190 14742
rect 10254 14678 10270 14742
rect 10334 14678 10350 14742
rect 10414 14678 10430 14742
rect 10494 14678 10510 14742
rect 10574 14678 10590 14742
rect 10654 14678 10670 14742
rect 10734 14678 10750 14742
rect 10814 14678 10830 14742
rect 10894 14678 10910 14742
rect 10974 14678 10990 14742
rect 11054 14678 11070 14742
rect 11134 14678 11150 14742
rect 11214 14678 11230 14742
rect 11294 14678 11310 14742
rect 11374 14678 11390 14742
rect 11454 14678 11470 14742
rect 11534 14678 11550 14742
rect 11614 14678 11630 14742
rect 11694 14678 11710 14742
rect 11774 14678 11790 14742
rect 11854 14678 11870 14742
rect 11934 14678 11950 14742
rect 12014 14678 12030 14742
rect 12094 14678 12110 14742
rect 12174 14678 12190 14742
rect 12254 14678 12270 14742
rect 12334 14678 12350 14742
rect 12414 14678 12430 14742
rect 12494 14678 12510 14742
rect 12574 14678 12590 14742
rect 12654 14678 12670 14742
rect 12734 14678 12750 14742
rect 12814 14678 12830 14742
rect 12894 14678 12910 14742
rect 12974 14678 12990 14742
rect 13054 14678 13070 14742
rect 13134 14678 13150 14742
rect 13214 14678 13230 14742
rect 13294 14678 13310 14742
rect 13374 14678 13390 14742
rect 13454 14678 13470 14742
rect 13534 14678 13550 14742
rect 13614 14678 13630 14742
rect 13694 14678 13710 14742
rect 13774 14678 13790 14742
rect 13854 14678 13870 14742
rect 13934 14678 13950 14742
rect 14014 14678 14030 14742
rect 14094 14678 14110 14742
rect 14174 14678 14190 14742
rect 14254 14678 14270 14742
rect 14334 14678 14350 14742
rect 14414 14678 14430 14742
rect 14494 14678 14510 14742
rect 14574 14678 14590 14742
rect 14654 14678 14670 14742
rect 14734 14678 14750 14742
rect 14814 14678 14830 14742
rect 14894 14678 15000 14742
rect 10151 14661 15000 14678
rect 10151 14597 10190 14661
rect 10254 14597 10270 14661
rect 10334 14597 10350 14661
rect 10414 14597 10430 14661
rect 10494 14597 10510 14661
rect 10574 14597 10590 14661
rect 10654 14597 10670 14661
rect 10734 14597 10750 14661
rect 10814 14597 10830 14661
rect 10894 14597 10910 14661
rect 10974 14597 10990 14661
rect 11054 14597 11070 14661
rect 11134 14597 11150 14661
rect 11214 14597 11230 14661
rect 11294 14597 11310 14661
rect 11374 14597 11390 14661
rect 11454 14597 11470 14661
rect 11534 14597 11550 14661
rect 11614 14597 11630 14661
rect 11694 14597 11710 14661
rect 11774 14597 11790 14661
rect 11854 14597 11870 14661
rect 11934 14597 11950 14661
rect 12014 14597 12030 14661
rect 12094 14597 12110 14661
rect 12174 14597 12190 14661
rect 12254 14597 12270 14661
rect 12334 14597 12350 14661
rect 12414 14597 12430 14661
rect 12494 14597 12510 14661
rect 12574 14597 12590 14661
rect 12654 14597 12670 14661
rect 12734 14597 12750 14661
rect 12814 14597 12830 14661
rect 12894 14597 12910 14661
rect 12974 14597 12990 14661
rect 13054 14597 13070 14661
rect 13134 14597 13150 14661
rect 13214 14597 13230 14661
rect 13294 14597 13310 14661
rect 13374 14597 13390 14661
rect 13454 14597 13470 14661
rect 13534 14597 13550 14661
rect 13614 14597 13630 14661
rect 13694 14597 13710 14661
rect 13774 14597 13790 14661
rect 13854 14597 13870 14661
rect 13934 14597 13950 14661
rect 14014 14597 14030 14661
rect 14094 14597 14110 14661
rect 14174 14597 14190 14661
rect 14254 14597 14270 14661
rect 14334 14597 14350 14661
rect 14414 14597 14430 14661
rect 14494 14597 14510 14661
rect 14574 14597 14590 14661
rect 14654 14597 14670 14661
rect 14734 14597 14750 14661
rect 14814 14597 14830 14661
rect 14894 14597 15000 14661
rect 10151 14579 15000 14597
rect 10151 14515 10190 14579
rect 10254 14515 10270 14579
rect 10334 14515 10350 14579
rect 10414 14515 10430 14579
rect 10494 14515 10510 14579
rect 10574 14515 10590 14579
rect 10654 14515 10670 14579
rect 10734 14515 10750 14579
rect 10814 14515 10830 14579
rect 10894 14515 10910 14579
rect 10974 14515 10990 14579
rect 11054 14515 11070 14579
rect 11134 14515 11150 14579
rect 11214 14515 11230 14579
rect 11294 14515 11310 14579
rect 11374 14515 11390 14579
rect 11454 14515 11470 14579
rect 11534 14515 11550 14579
rect 11614 14515 11630 14579
rect 11694 14515 11710 14579
rect 11774 14515 11790 14579
rect 11854 14515 11870 14579
rect 11934 14515 11950 14579
rect 12014 14515 12030 14579
rect 12094 14515 12110 14579
rect 12174 14515 12190 14579
rect 12254 14515 12270 14579
rect 12334 14515 12350 14579
rect 12414 14515 12430 14579
rect 12494 14515 12510 14579
rect 12574 14515 12590 14579
rect 12654 14515 12670 14579
rect 12734 14515 12750 14579
rect 12814 14515 12830 14579
rect 12894 14515 12910 14579
rect 12974 14515 12990 14579
rect 13054 14515 13070 14579
rect 13134 14515 13150 14579
rect 13214 14515 13230 14579
rect 13294 14515 13310 14579
rect 13374 14515 13390 14579
rect 13454 14515 13470 14579
rect 13534 14515 13550 14579
rect 13614 14515 13630 14579
rect 13694 14515 13710 14579
rect 13774 14515 13790 14579
rect 13854 14515 13870 14579
rect 13934 14515 13950 14579
rect 14014 14515 14030 14579
rect 14094 14515 14110 14579
rect 14174 14515 14190 14579
rect 14254 14515 14270 14579
rect 14334 14515 14350 14579
rect 14414 14515 14430 14579
rect 14494 14515 14510 14579
rect 14574 14515 14590 14579
rect 14654 14515 14670 14579
rect 14734 14515 14750 14579
rect 14814 14515 14830 14579
rect 14894 14515 15000 14579
rect 10151 14497 15000 14515
rect 10151 14433 10190 14497
rect 10254 14433 10270 14497
rect 10334 14433 10350 14497
rect 10414 14433 10430 14497
rect 10494 14433 10510 14497
rect 10574 14433 10590 14497
rect 10654 14433 10670 14497
rect 10734 14433 10750 14497
rect 10814 14433 10830 14497
rect 10894 14433 10910 14497
rect 10974 14433 10990 14497
rect 11054 14433 11070 14497
rect 11134 14433 11150 14497
rect 11214 14433 11230 14497
rect 11294 14433 11310 14497
rect 11374 14433 11390 14497
rect 11454 14433 11470 14497
rect 11534 14433 11550 14497
rect 11614 14433 11630 14497
rect 11694 14433 11710 14497
rect 11774 14433 11790 14497
rect 11854 14433 11870 14497
rect 11934 14433 11950 14497
rect 12014 14433 12030 14497
rect 12094 14433 12110 14497
rect 12174 14433 12190 14497
rect 12254 14433 12270 14497
rect 12334 14433 12350 14497
rect 12414 14433 12430 14497
rect 12494 14433 12510 14497
rect 12574 14433 12590 14497
rect 12654 14433 12670 14497
rect 12734 14433 12750 14497
rect 12814 14433 12830 14497
rect 12894 14433 12910 14497
rect 12974 14433 12990 14497
rect 13054 14433 13070 14497
rect 13134 14433 13150 14497
rect 13214 14433 13230 14497
rect 13294 14433 13310 14497
rect 13374 14433 13390 14497
rect 13454 14433 13470 14497
rect 13534 14433 13550 14497
rect 13614 14433 13630 14497
rect 13694 14433 13710 14497
rect 13774 14433 13790 14497
rect 13854 14433 13870 14497
rect 13934 14433 13950 14497
rect 14014 14433 14030 14497
rect 14094 14433 14110 14497
rect 14174 14433 14190 14497
rect 14254 14433 14270 14497
rect 14334 14433 14350 14497
rect 14414 14433 14430 14497
rect 14494 14433 14510 14497
rect 14574 14433 14590 14497
rect 14654 14433 14670 14497
rect 14734 14433 14750 14497
rect 14814 14433 14830 14497
rect 14894 14433 15000 14497
rect 10151 14415 15000 14433
rect 10151 14351 10190 14415
rect 10254 14351 10270 14415
rect 10334 14351 10350 14415
rect 10414 14351 10430 14415
rect 10494 14351 10510 14415
rect 10574 14351 10590 14415
rect 10654 14351 10670 14415
rect 10734 14351 10750 14415
rect 10814 14351 10830 14415
rect 10894 14351 10910 14415
rect 10974 14351 10990 14415
rect 11054 14351 11070 14415
rect 11134 14351 11150 14415
rect 11214 14351 11230 14415
rect 11294 14351 11310 14415
rect 11374 14351 11390 14415
rect 11454 14351 11470 14415
rect 11534 14351 11550 14415
rect 11614 14351 11630 14415
rect 11694 14351 11710 14415
rect 11774 14351 11790 14415
rect 11854 14351 11870 14415
rect 11934 14351 11950 14415
rect 12014 14351 12030 14415
rect 12094 14351 12110 14415
rect 12174 14351 12190 14415
rect 12254 14351 12270 14415
rect 12334 14351 12350 14415
rect 12414 14351 12430 14415
rect 12494 14351 12510 14415
rect 12574 14351 12590 14415
rect 12654 14351 12670 14415
rect 12734 14351 12750 14415
rect 12814 14351 12830 14415
rect 12894 14351 12910 14415
rect 12974 14351 12990 14415
rect 13054 14351 13070 14415
rect 13134 14351 13150 14415
rect 13214 14351 13230 14415
rect 13294 14351 13310 14415
rect 13374 14351 13390 14415
rect 13454 14351 13470 14415
rect 13534 14351 13550 14415
rect 13614 14351 13630 14415
rect 13694 14351 13710 14415
rect 13774 14351 13790 14415
rect 13854 14351 13870 14415
rect 13934 14351 13950 14415
rect 14014 14351 14030 14415
rect 14094 14351 14110 14415
rect 14174 14351 14190 14415
rect 14254 14351 14270 14415
rect 14334 14351 14350 14415
rect 14414 14351 14430 14415
rect 14494 14351 14510 14415
rect 14574 14351 14590 14415
rect 14654 14351 14670 14415
rect 14734 14351 14750 14415
rect 14814 14351 14830 14415
rect 14894 14351 15000 14415
rect 10151 14333 15000 14351
rect 10151 14269 10190 14333
rect 10254 14269 10270 14333
rect 10334 14269 10350 14333
rect 10414 14269 10430 14333
rect 10494 14269 10510 14333
rect 10574 14269 10590 14333
rect 10654 14269 10670 14333
rect 10734 14269 10750 14333
rect 10814 14269 10830 14333
rect 10894 14269 10910 14333
rect 10974 14269 10990 14333
rect 11054 14269 11070 14333
rect 11134 14269 11150 14333
rect 11214 14269 11230 14333
rect 11294 14269 11310 14333
rect 11374 14269 11390 14333
rect 11454 14269 11470 14333
rect 11534 14269 11550 14333
rect 11614 14269 11630 14333
rect 11694 14269 11710 14333
rect 11774 14269 11790 14333
rect 11854 14269 11870 14333
rect 11934 14269 11950 14333
rect 12014 14269 12030 14333
rect 12094 14269 12110 14333
rect 12174 14269 12190 14333
rect 12254 14269 12270 14333
rect 12334 14269 12350 14333
rect 12414 14269 12430 14333
rect 12494 14269 12510 14333
rect 12574 14269 12590 14333
rect 12654 14269 12670 14333
rect 12734 14269 12750 14333
rect 12814 14269 12830 14333
rect 12894 14269 12910 14333
rect 12974 14269 12990 14333
rect 13054 14269 13070 14333
rect 13134 14269 13150 14333
rect 13214 14269 13230 14333
rect 13294 14269 13310 14333
rect 13374 14269 13390 14333
rect 13454 14269 13470 14333
rect 13534 14269 13550 14333
rect 13614 14269 13630 14333
rect 13694 14269 13710 14333
rect 13774 14269 13790 14333
rect 13854 14269 13870 14333
rect 13934 14269 13950 14333
rect 14014 14269 14030 14333
rect 14094 14269 14110 14333
rect 14174 14269 14190 14333
rect 14254 14269 14270 14333
rect 14334 14269 14350 14333
rect 14414 14269 14430 14333
rect 14494 14269 14510 14333
rect 14574 14269 14590 14333
rect 14654 14269 14670 14333
rect 14734 14269 14750 14333
rect 14814 14269 14830 14333
rect 14894 14269 15000 14333
rect 10151 14251 15000 14269
rect 10151 14187 10190 14251
rect 10254 14187 10270 14251
rect 10334 14187 10350 14251
rect 10414 14187 10430 14251
rect 10494 14187 10510 14251
rect 10574 14187 10590 14251
rect 10654 14187 10670 14251
rect 10734 14187 10750 14251
rect 10814 14187 10830 14251
rect 10894 14187 10910 14251
rect 10974 14187 10990 14251
rect 11054 14187 11070 14251
rect 11134 14187 11150 14251
rect 11214 14187 11230 14251
rect 11294 14187 11310 14251
rect 11374 14187 11390 14251
rect 11454 14187 11470 14251
rect 11534 14187 11550 14251
rect 11614 14187 11630 14251
rect 11694 14187 11710 14251
rect 11774 14187 11790 14251
rect 11854 14187 11870 14251
rect 11934 14187 11950 14251
rect 12014 14187 12030 14251
rect 12094 14187 12110 14251
rect 12174 14187 12190 14251
rect 12254 14187 12270 14251
rect 12334 14187 12350 14251
rect 12414 14187 12430 14251
rect 12494 14187 12510 14251
rect 12574 14187 12590 14251
rect 12654 14187 12670 14251
rect 12734 14187 12750 14251
rect 12814 14187 12830 14251
rect 12894 14187 12910 14251
rect 12974 14187 12990 14251
rect 13054 14187 13070 14251
rect 13134 14187 13150 14251
rect 13214 14187 13230 14251
rect 13294 14187 13310 14251
rect 13374 14187 13390 14251
rect 13454 14187 13470 14251
rect 13534 14187 13550 14251
rect 13614 14187 13630 14251
rect 13694 14187 13710 14251
rect 13774 14187 13790 14251
rect 13854 14187 13870 14251
rect 13934 14187 13950 14251
rect 14014 14187 14030 14251
rect 14094 14187 14110 14251
rect 14174 14187 14190 14251
rect 14254 14187 14270 14251
rect 14334 14187 14350 14251
rect 14414 14187 14430 14251
rect 14494 14187 14510 14251
rect 14574 14187 14590 14251
rect 14654 14187 14670 14251
rect 14734 14187 14750 14251
rect 14814 14187 14830 14251
rect 14894 14187 15000 14251
rect 10151 14169 15000 14187
rect 10151 14105 10190 14169
rect 10254 14105 10270 14169
rect 10334 14105 10350 14169
rect 10414 14105 10430 14169
rect 10494 14105 10510 14169
rect 10574 14105 10590 14169
rect 10654 14105 10670 14169
rect 10734 14105 10750 14169
rect 10814 14105 10830 14169
rect 10894 14105 10910 14169
rect 10974 14105 10990 14169
rect 11054 14105 11070 14169
rect 11134 14105 11150 14169
rect 11214 14105 11230 14169
rect 11294 14105 11310 14169
rect 11374 14105 11390 14169
rect 11454 14105 11470 14169
rect 11534 14105 11550 14169
rect 11614 14105 11630 14169
rect 11694 14105 11710 14169
rect 11774 14105 11790 14169
rect 11854 14105 11870 14169
rect 11934 14105 11950 14169
rect 12014 14105 12030 14169
rect 12094 14105 12110 14169
rect 12174 14105 12190 14169
rect 12254 14105 12270 14169
rect 12334 14105 12350 14169
rect 12414 14105 12430 14169
rect 12494 14105 12510 14169
rect 12574 14105 12590 14169
rect 12654 14105 12670 14169
rect 12734 14105 12750 14169
rect 12814 14105 12830 14169
rect 12894 14105 12910 14169
rect 12974 14105 12990 14169
rect 13054 14105 13070 14169
rect 13134 14105 13150 14169
rect 13214 14105 13230 14169
rect 13294 14105 13310 14169
rect 13374 14105 13390 14169
rect 13454 14105 13470 14169
rect 13534 14105 13550 14169
rect 13614 14105 13630 14169
rect 13694 14105 13710 14169
rect 13774 14105 13790 14169
rect 13854 14105 13870 14169
rect 13934 14105 13950 14169
rect 14014 14105 14030 14169
rect 14094 14105 14110 14169
rect 14174 14105 14190 14169
rect 14254 14105 14270 14169
rect 14334 14105 14350 14169
rect 14414 14105 14430 14169
rect 14494 14105 14510 14169
rect 14574 14105 14590 14169
rect 14654 14105 14670 14169
rect 14734 14105 14750 14169
rect 14814 14105 14830 14169
rect 14894 14105 15000 14169
rect 10151 14087 15000 14105
rect 10151 14023 10190 14087
rect 10254 14023 10270 14087
rect 10334 14023 10350 14087
rect 10414 14023 10430 14087
rect 10494 14023 10510 14087
rect 10574 14023 10590 14087
rect 10654 14023 10670 14087
rect 10734 14023 10750 14087
rect 10814 14023 10830 14087
rect 10894 14023 10910 14087
rect 10974 14023 10990 14087
rect 11054 14023 11070 14087
rect 11134 14023 11150 14087
rect 11214 14023 11230 14087
rect 11294 14023 11310 14087
rect 11374 14023 11390 14087
rect 11454 14023 11470 14087
rect 11534 14023 11550 14087
rect 11614 14023 11630 14087
rect 11694 14023 11710 14087
rect 11774 14023 11790 14087
rect 11854 14023 11870 14087
rect 11934 14023 11950 14087
rect 12014 14023 12030 14087
rect 12094 14023 12110 14087
rect 12174 14023 12190 14087
rect 12254 14023 12270 14087
rect 12334 14023 12350 14087
rect 12414 14023 12430 14087
rect 12494 14023 12510 14087
rect 12574 14023 12590 14087
rect 12654 14023 12670 14087
rect 12734 14023 12750 14087
rect 12814 14023 12830 14087
rect 12894 14023 12910 14087
rect 12974 14023 12990 14087
rect 13054 14023 13070 14087
rect 13134 14023 13150 14087
rect 13214 14023 13230 14087
rect 13294 14023 13310 14087
rect 13374 14023 13390 14087
rect 13454 14023 13470 14087
rect 13534 14023 13550 14087
rect 13614 14023 13630 14087
rect 13694 14023 13710 14087
rect 13774 14023 13790 14087
rect 13854 14023 13870 14087
rect 13934 14023 13950 14087
rect 14014 14023 14030 14087
rect 14094 14023 14110 14087
rect 14174 14023 14190 14087
rect 14254 14023 14270 14087
rect 14334 14023 14350 14087
rect 14414 14023 14430 14087
rect 14494 14023 14510 14087
rect 14574 14023 14590 14087
rect 14654 14023 14670 14087
rect 14734 14023 14750 14087
rect 14814 14023 14830 14087
rect 14894 14023 15000 14087
rect 10151 14005 15000 14023
rect 10151 13941 10190 14005
rect 10254 13941 10270 14005
rect 10334 13941 10350 14005
rect 10414 13941 10430 14005
rect 10494 13941 10510 14005
rect 10574 13941 10590 14005
rect 10654 13941 10670 14005
rect 10734 13941 10750 14005
rect 10814 13941 10830 14005
rect 10894 13941 10910 14005
rect 10974 13941 10990 14005
rect 11054 13941 11070 14005
rect 11134 13941 11150 14005
rect 11214 13941 11230 14005
rect 11294 13941 11310 14005
rect 11374 13941 11390 14005
rect 11454 13941 11470 14005
rect 11534 13941 11550 14005
rect 11614 13941 11630 14005
rect 11694 13941 11710 14005
rect 11774 13941 11790 14005
rect 11854 13941 11870 14005
rect 11934 13941 11950 14005
rect 12014 13941 12030 14005
rect 12094 13941 12110 14005
rect 12174 13941 12190 14005
rect 12254 13941 12270 14005
rect 12334 13941 12350 14005
rect 12414 13941 12430 14005
rect 12494 13941 12510 14005
rect 12574 13941 12590 14005
rect 12654 13941 12670 14005
rect 12734 13941 12750 14005
rect 12814 13941 12830 14005
rect 12894 13941 12910 14005
rect 12974 13941 12990 14005
rect 13054 13941 13070 14005
rect 13134 13941 13150 14005
rect 13214 13941 13230 14005
rect 13294 13941 13310 14005
rect 13374 13941 13390 14005
rect 13454 13941 13470 14005
rect 13534 13941 13550 14005
rect 13614 13941 13630 14005
rect 13694 13941 13710 14005
rect 13774 13941 13790 14005
rect 13854 13941 13870 14005
rect 13934 13941 13950 14005
rect 14014 13941 14030 14005
rect 14094 13941 14110 14005
rect 14174 13941 14190 14005
rect 14254 13941 14270 14005
rect 14334 13941 14350 14005
rect 14414 13941 14430 14005
rect 14494 13941 14510 14005
rect 14574 13941 14590 14005
rect 14654 13941 14670 14005
rect 14734 13941 14750 14005
rect 14814 13941 14830 14005
rect 14894 13941 15000 14005
rect 10151 13923 15000 13941
rect 10151 13859 10190 13923
rect 10254 13859 10270 13923
rect 10334 13859 10350 13923
rect 10414 13859 10430 13923
rect 10494 13859 10510 13923
rect 10574 13859 10590 13923
rect 10654 13859 10670 13923
rect 10734 13859 10750 13923
rect 10814 13859 10830 13923
rect 10894 13859 10910 13923
rect 10974 13859 10990 13923
rect 11054 13859 11070 13923
rect 11134 13859 11150 13923
rect 11214 13859 11230 13923
rect 11294 13859 11310 13923
rect 11374 13859 11390 13923
rect 11454 13859 11470 13923
rect 11534 13859 11550 13923
rect 11614 13859 11630 13923
rect 11694 13859 11710 13923
rect 11774 13859 11790 13923
rect 11854 13859 11870 13923
rect 11934 13859 11950 13923
rect 12014 13859 12030 13923
rect 12094 13859 12110 13923
rect 12174 13859 12190 13923
rect 12254 13859 12270 13923
rect 12334 13859 12350 13923
rect 12414 13859 12430 13923
rect 12494 13859 12510 13923
rect 12574 13859 12590 13923
rect 12654 13859 12670 13923
rect 12734 13859 12750 13923
rect 12814 13859 12830 13923
rect 12894 13859 12910 13923
rect 12974 13859 12990 13923
rect 13054 13859 13070 13923
rect 13134 13859 13150 13923
rect 13214 13859 13230 13923
rect 13294 13859 13310 13923
rect 13374 13859 13390 13923
rect 13454 13859 13470 13923
rect 13534 13859 13550 13923
rect 13614 13859 13630 13923
rect 13694 13859 13710 13923
rect 13774 13859 13790 13923
rect 13854 13859 13870 13923
rect 13934 13859 13950 13923
rect 14014 13859 14030 13923
rect 14094 13859 14110 13923
rect 14174 13859 14190 13923
rect 14254 13859 14270 13923
rect 14334 13859 14350 13923
rect 14414 13859 14430 13923
rect 14494 13859 14510 13923
rect 14574 13859 14590 13923
rect 14654 13859 14670 13923
rect 14734 13859 14750 13923
rect 14814 13859 14830 13923
rect 14894 13859 15000 13923
rect 10151 13841 15000 13859
rect 10151 13777 10190 13841
rect 10254 13777 10270 13841
rect 10334 13777 10350 13841
rect 10414 13777 10430 13841
rect 10494 13777 10510 13841
rect 10574 13777 10590 13841
rect 10654 13777 10670 13841
rect 10734 13777 10750 13841
rect 10814 13777 10830 13841
rect 10894 13777 10910 13841
rect 10974 13777 10990 13841
rect 11054 13777 11070 13841
rect 11134 13777 11150 13841
rect 11214 13777 11230 13841
rect 11294 13777 11310 13841
rect 11374 13777 11390 13841
rect 11454 13777 11470 13841
rect 11534 13777 11550 13841
rect 11614 13777 11630 13841
rect 11694 13777 11710 13841
rect 11774 13777 11790 13841
rect 11854 13777 11870 13841
rect 11934 13777 11950 13841
rect 12014 13777 12030 13841
rect 12094 13777 12110 13841
rect 12174 13777 12190 13841
rect 12254 13777 12270 13841
rect 12334 13777 12350 13841
rect 12414 13777 12430 13841
rect 12494 13777 12510 13841
rect 12574 13777 12590 13841
rect 12654 13777 12670 13841
rect 12734 13777 12750 13841
rect 12814 13777 12830 13841
rect 12894 13777 12910 13841
rect 12974 13777 12990 13841
rect 13054 13777 13070 13841
rect 13134 13777 13150 13841
rect 13214 13777 13230 13841
rect 13294 13777 13310 13841
rect 13374 13777 13390 13841
rect 13454 13777 13470 13841
rect 13534 13777 13550 13841
rect 13614 13777 13630 13841
rect 13694 13777 13710 13841
rect 13774 13777 13790 13841
rect 13854 13777 13870 13841
rect 13934 13777 13950 13841
rect 14014 13777 14030 13841
rect 14094 13777 14110 13841
rect 14174 13777 14190 13841
rect 14254 13777 14270 13841
rect 14334 13777 14350 13841
rect 14414 13777 14430 13841
rect 14494 13777 14510 13841
rect 14574 13777 14590 13841
rect 14654 13777 14670 13841
rect 14734 13777 14750 13841
rect 14814 13777 14830 13841
rect 14894 13777 15000 13841
rect 10151 13759 15000 13777
rect 10151 13695 10190 13759
rect 10254 13695 10270 13759
rect 10334 13695 10350 13759
rect 10414 13695 10430 13759
rect 10494 13695 10510 13759
rect 10574 13695 10590 13759
rect 10654 13695 10670 13759
rect 10734 13695 10750 13759
rect 10814 13695 10830 13759
rect 10894 13695 10910 13759
rect 10974 13695 10990 13759
rect 11054 13695 11070 13759
rect 11134 13695 11150 13759
rect 11214 13695 11230 13759
rect 11294 13695 11310 13759
rect 11374 13695 11390 13759
rect 11454 13695 11470 13759
rect 11534 13695 11550 13759
rect 11614 13695 11630 13759
rect 11694 13695 11710 13759
rect 11774 13695 11790 13759
rect 11854 13695 11870 13759
rect 11934 13695 11950 13759
rect 12014 13695 12030 13759
rect 12094 13695 12110 13759
rect 12174 13695 12190 13759
rect 12254 13695 12270 13759
rect 12334 13695 12350 13759
rect 12414 13695 12430 13759
rect 12494 13695 12510 13759
rect 12574 13695 12590 13759
rect 12654 13695 12670 13759
rect 12734 13695 12750 13759
rect 12814 13695 12830 13759
rect 12894 13695 12910 13759
rect 12974 13695 12990 13759
rect 13054 13695 13070 13759
rect 13134 13695 13150 13759
rect 13214 13695 13230 13759
rect 13294 13695 13310 13759
rect 13374 13695 13390 13759
rect 13454 13695 13470 13759
rect 13534 13695 13550 13759
rect 13614 13695 13630 13759
rect 13694 13695 13710 13759
rect 13774 13695 13790 13759
rect 13854 13695 13870 13759
rect 13934 13695 13950 13759
rect 14014 13695 14030 13759
rect 14094 13695 14110 13759
rect 14174 13695 14190 13759
rect 14254 13695 14270 13759
rect 14334 13695 14350 13759
rect 14414 13695 14430 13759
rect 14494 13695 14510 13759
rect 14574 13695 14590 13759
rect 14654 13695 14670 13759
rect 14734 13695 14750 13759
rect 14814 13695 14830 13759
rect 14894 13695 15000 13759
rect 10151 13677 15000 13695
rect 10151 13613 10190 13677
rect 10254 13613 10270 13677
rect 10334 13613 10350 13677
rect 10414 13613 10430 13677
rect 10494 13613 10510 13677
rect 10574 13613 10590 13677
rect 10654 13613 10670 13677
rect 10734 13613 10750 13677
rect 10814 13613 10830 13677
rect 10894 13613 10910 13677
rect 10974 13613 10990 13677
rect 11054 13613 11070 13677
rect 11134 13613 11150 13677
rect 11214 13613 11230 13677
rect 11294 13613 11310 13677
rect 11374 13613 11390 13677
rect 11454 13613 11470 13677
rect 11534 13613 11550 13677
rect 11614 13613 11630 13677
rect 11694 13613 11710 13677
rect 11774 13613 11790 13677
rect 11854 13613 11870 13677
rect 11934 13613 11950 13677
rect 12014 13613 12030 13677
rect 12094 13613 12110 13677
rect 12174 13613 12190 13677
rect 12254 13613 12270 13677
rect 12334 13613 12350 13677
rect 12414 13613 12430 13677
rect 12494 13613 12510 13677
rect 12574 13613 12590 13677
rect 12654 13613 12670 13677
rect 12734 13613 12750 13677
rect 12814 13613 12830 13677
rect 12894 13613 12910 13677
rect 12974 13613 12990 13677
rect 13054 13613 13070 13677
rect 13134 13613 13150 13677
rect 13214 13613 13230 13677
rect 13294 13613 13310 13677
rect 13374 13613 13390 13677
rect 13454 13613 13470 13677
rect 13534 13613 13550 13677
rect 13614 13613 13630 13677
rect 13694 13613 13710 13677
rect 13774 13613 13790 13677
rect 13854 13613 13870 13677
rect 13934 13613 13950 13677
rect 14014 13613 14030 13677
rect 14094 13613 14110 13677
rect 14174 13613 14190 13677
rect 14254 13613 14270 13677
rect 14334 13613 14350 13677
rect 14414 13613 14430 13677
rect 14494 13613 14510 13677
rect 14574 13613 14590 13677
rect 14654 13613 14670 13677
rect 14734 13613 14750 13677
rect 14814 13613 14830 13677
rect 14894 13613 15000 13677
rect 10151 13612 15000 13613
rect 0 13607 254 13612
rect 14746 13607 15000 13612
rect 0 13304 4895 13307
rect 0 13240 126 13304
rect 190 13240 207 13304
rect 271 13240 288 13304
rect 352 13240 369 13304
rect 433 13240 450 13304
rect 514 13240 531 13304
rect 595 13240 612 13304
rect 676 13240 693 13304
rect 757 13240 774 13304
rect 838 13240 855 13304
rect 919 13240 936 13304
rect 1000 13240 1017 13304
rect 1081 13240 1098 13304
rect 1162 13240 1179 13304
rect 1243 13240 1260 13304
rect 1324 13240 1341 13304
rect 1405 13240 1422 13304
rect 1486 13240 1503 13304
rect 1567 13240 1584 13304
rect 1648 13240 1665 13304
rect 1729 13240 1746 13304
rect 1810 13240 1827 13304
rect 1891 13240 1908 13304
rect 1972 13240 1989 13304
rect 2053 13240 2070 13304
rect 2134 13240 2151 13304
rect 2215 13240 2232 13304
rect 2296 13240 2313 13304
rect 2377 13240 2394 13304
rect 2458 13240 2475 13304
rect 2539 13240 2556 13304
rect 2620 13240 2637 13304
rect 2701 13240 2718 13304
rect 2782 13240 2799 13304
rect 2863 13240 2880 13304
rect 2944 13240 2961 13304
rect 3025 13240 3042 13304
rect 3106 13240 3123 13304
rect 3187 13240 3204 13304
rect 3268 13240 3285 13304
rect 3349 13240 3366 13304
rect 3430 13240 3447 13304
rect 3511 13240 3528 13304
rect 3592 13240 3609 13304
rect 3673 13240 3690 13304
rect 3754 13240 3771 13304
rect 3835 13240 3852 13304
rect 3916 13240 3933 13304
rect 3997 13240 4014 13304
rect 4078 13240 4095 13304
rect 4159 13240 4176 13304
rect 4240 13240 4257 13304
rect 4321 13240 4338 13304
rect 4402 13240 4420 13304
rect 4484 13240 4502 13304
rect 4566 13240 4584 13304
rect 4648 13240 4666 13304
rect 4730 13240 4748 13304
rect 4812 13240 4830 13304
rect 4894 13240 4895 13304
rect 0 13222 4895 13240
rect 0 13158 126 13222
rect 190 13158 207 13222
rect 271 13158 288 13222
rect 352 13158 369 13222
rect 433 13158 450 13222
rect 514 13158 531 13222
rect 595 13158 612 13222
rect 676 13158 693 13222
rect 757 13158 774 13222
rect 838 13158 855 13222
rect 919 13158 936 13222
rect 1000 13158 1017 13222
rect 1081 13158 1098 13222
rect 1162 13158 1179 13222
rect 1243 13158 1260 13222
rect 1324 13158 1341 13222
rect 1405 13158 1422 13222
rect 1486 13158 1503 13222
rect 1567 13158 1584 13222
rect 1648 13158 1665 13222
rect 1729 13158 1746 13222
rect 1810 13158 1827 13222
rect 1891 13158 1908 13222
rect 1972 13158 1989 13222
rect 2053 13158 2070 13222
rect 2134 13158 2151 13222
rect 2215 13158 2232 13222
rect 2296 13158 2313 13222
rect 2377 13158 2394 13222
rect 2458 13158 2475 13222
rect 2539 13158 2556 13222
rect 2620 13158 2637 13222
rect 2701 13158 2718 13222
rect 2782 13158 2799 13222
rect 2863 13158 2880 13222
rect 2944 13158 2961 13222
rect 3025 13158 3042 13222
rect 3106 13158 3123 13222
rect 3187 13158 3204 13222
rect 3268 13158 3285 13222
rect 3349 13158 3366 13222
rect 3430 13158 3447 13222
rect 3511 13158 3528 13222
rect 3592 13158 3609 13222
rect 3673 13158 3690 13222
rect 3754 13158 3771 13222
rect 3835 13158 3852 13222
rect 3916 13158 3933 13222
rect 3997 13158 4014 13222
rect 4078 13158 4095 13222
rect 4159 13158 4176 13222
rect 4240 13158 4257 13222
rect 4321 13158 4338 13222
rect 4402 13158 4420 13222
rect 4484 13158 4502 13222
rect 4566 13158 4584 13222
rect 4648 13158 4666 13222
rect 4730 13158 4748 13222
rect 4812 13158 4830 13222
rect 4894 13158 4895 13222
rect 0 13140 4895 13158
rect 0 13076 126 13140
rect 190 13076 207 13140
rect 271 13076 288 13140
rect 352 13076 369 13140
rect 433 13076 450 13140
rect 514 13076 531 13140
rect 595 13076 612 13140
rect 676 13076 693 13140
rect 757 13076 774 13140
rect 838 13076 855 13140
rect 919 13076 936 13140
rect 1000 13076 1017 13140
rect 1081 13076 1098 13140
rect 1162 13076 1179 13140
rect 1243 13076 1260 13140
rect 1324 13076 1341 13140
rect 1405 13076 1422 13140
rect 1486 13076 1503 13140
rect 1567 13076 1584 13140
rect 1648 13076 1665 13140
rect 1729 13076 1746 13140
rect 1810 13076 1827 13140
rect 1891 13076 1908 13140
rect 1972 13076 1989 13140
rect 2053 13076 2070 13140
rect 2134 13076 2151 13140
rect 2215 13076 2232 13140
rect 2296 13076 2313 13140
rect 2377 13076 2394 13140
rect 2458 13076 2475 13140
rect 2539 13076 2556 13140
rect 2620 13076 2637 13140
rect 2701 13076 2718 13140
rect 2782 13076 2799 13140
rect 2863 13076 2880 13140
rect 2944 13076 2961 13140
rect 3025 13076 3042 13140
rect 3106 13076 3123 13140
rect 3187 13076 3204 13140
rect 3268 13076 3285 13140
rect 3349 13076 3366 13140
rect 3430 13076 3447 13140
rect 3511 13076 3528 13140
rect 3592 13076 3609 13140
rect 3673 13076 3690 13140
rect 3754 13076 3771 13140
rect 3835 13076 3852 13140
rect 3916 13076 3933 13140
rect 3997 13076 4014 13140
rect 4078 13076 4095 13140
rect 4159 13076 4176 13140
rect 4240 13076 4257 13140
rect 4321 13076 4338 13140
rect 4402 13076 4420 13140
rect 4484 13076 4502 13140
rect 4566 13076 4584 13140
rect 4648 13076 4666 13140
rect 4730 13076 4748 13140
rect 4812 13076 4830 13140
rect 4894 13076 4895 13140
rect 0 13058 4895 13076
rect 0 12994 126 13058
rect 190 12994 207 13058
rect 271 12994 288 13058
rect 352 12994 369 13058
rect 433 12994 450 13058
rect 514 12994 531 13058
rect 595 12994 612 13058
rect 676 12994 693 13058
rect 757 12994 774 13058
rect 838 12994 855 13058
rect 919 12994 936 13058
rect 1000 12994 1017 13058
rect 1081 12994 1098 13058
rect 1162 12994 1179 13058
rect 1243 12994 1260 13058
rect 1324 12994 1341 13058
rect 1405 12994 1422 13058
rect 1486 12994 1503 13058
rect 1567 12994 1584 13058
rect 1648 12994 1665 13058
rect 1729 12994 1746 13058
rect 1810 12994 1827 13058
rect 1891 12994 1908 13058
rect 1972 12994 1989 13058
rect 2053 12994 2070 13058
rect 2134 12994 2151 13058
rect 2215 12994 2232 13058
rect 2296 12994 2313 13058
rect 2377 12994 2394 13058
rect 2458 12994 2475 13058
rect 2539 12994 2556 13058
rect 2620 12994 2637 13058
rect 2701 12994 2718 13058
rect 2782 12994 2799 13058
rect 2863 12994 2880 13058
rect 2944 12994 2961 13058
rect 3025 12994 3042 13058
rect 3106 12994 3123 13058
rect 3187 12994 3204 13058
rect 3268 12994 3285 13058
rect 3349 12994 3366 13058
rect 3430 12994 3447 13058
rect 3511 12994 3528 13058
rect 3592 12994 3609 13058
rect 3673 12994 3690 13058
rect 3754 12994 3771 13058
rect 3835 12994 3852 13058
rect 3916 12994 3933 13058
rect 3997 12994 4014 13058
rect 4078 12994 4095 13058
rect 4159 12994 4176 13058
rect 4240 12994 4257 13058
rect 4321 12994 4338 13058
rect 4402 12994 4420 13058
rect 4484 12994 4502 13058
rect 4566 12994 4584 13058
rect 4648 12994 4666 13058
rect 4730 12994 4748 13058
rect 4812 12994 4830 13058
rect 4894 12994 4895 13058
rect 0 12976 4895 12994
rect 0 12912 126 12976
rect 190 12912 207 12976
rect 271 12912 288 12976
rect 352 12912 369 12976
rect 433 12912 450 12976
rect 514 12912 531 12976
rect 595 12912 612 12976
rect 676 12912 693 12976
rect 757 12912 774 12976
rect 838 12912 855 12976
rect 919 12912 936 12976
rect 1000 12912 1017 12976
rect 1081 12912 1098 12976
rect 1162 12912 1179 12976
rect 1243 12912 1260 12976
rect 1324 12912 1341 12976
rect 1405 12912 1422 12976
rect 1486 12912 1503 12976
rect 1567 12912 1584 12976
rect 1648 12912 1665 12976
rect 1729 12912 1746 12976
rect 1810 12912 1827 12976
rect 1891 12912 1908 12976
rect 1972 12912 1989 12976
rect 2053 12912 2070 12976
rect 2134 12912 2151 12976
rect 2215 12912 2232 12976
rect 2296 12912 2313 12976
rect 2377 12912 2394 12976
rect 2458 12912 2475 12976
rect 2539 12912 2556 12976
rect 2620 12912 2637 12976
rect 2701 12912 2718 12976
rect 2782 12912 2799 12976
rect 2863 12912 2880 12976
rect 2944 12912 2961 12976
rect 3025 12912 3042 12976
rect 3106 12912 3123 12976
rect 3187 12912 3204 12976
rect 3268 12912 3285 12976
rect 3349 12912 3366 12976
rect 3430 12912 3447 12976
rect 3511 12912 3528 12976
rect 3592 12912 3609 12976
rect 3673 12912 3690 12976
rect 3754 12912 3771 12976
rect 3835 12912 3852 12976
rect 3916 12912 3933 12976
rect 3997 12912 4014 12976
rect 4078 12912 4095 12976
rect 4159 12912 4176 12976
rect 4240 12912 4257 12976
rect 4321 12912 4338 12976
rect 4402 12912 4420 12976
rect 4484 12912 4502 12976
rect 4566 12912 4584 12976
rect 4648 12912 4666 12976
rect 4730 12912 4748 12976
rect 4812 12912 4830 12976
rect 4894 12912 4895 12976
rect 0 12894 4895 12912
rect 0 12830 126 12894
rect 190 12830 207 12894
rect 271 12830 288 12894
rect 352 12830 369 12894
rect 433 12830 450 12894
rect 514 12830 531 12894
rect 595 12830 612 12894
rect 676 12830 693 12894
rect 757 12830 774 12894
rect 838 12830 855 12894
rect 919 12830 936 12894
rect 1000 12830 1017 12894
rect 1081 12830 1098 12894
rect 1162 12830 1179 12894
rect 1243 12830 1260 12894
rect 1324 12830 1341 12894
rect 1405 12830 1422 12894
rect 1486 12830 1503 12894
rect 1567 12830 1584 12894
rect 1648 12830 1665 12894
rect 1729 12830 1746 12894
rect 1810 12830 1827 12894
rect 1891 12830 1908 12894
rect 1972 12830 1989 12894
rect 2053 12830 2070 12894
rect 2134 12830 2151 12894
rect 2215 12830 2232 12894
rect 2296 12830 2313 12894
rect 2377 12830 2394 12894
rect 2458 12830 2475 12894
rect 2539 12830 2556 12894
rect 2620 12830 2637 12894
rect 2701 12830 2718 12894
rect 2782 12830 2799 12894
rect 2863 12830 2880 12894
rect 2944 12830 2961 12894
rect 3025 12830 3042 12894
rect 3106 12830 3123 12894
rect 3187 12830 3204 12894
rect 3268 12830 3285 12894
rect 3349 12830 3366 12894
rect 3430 12830 3447 12894
rect 3511 12830 3528 12894
rect 3592 12830 3609 12894
rect 3673 12830 3690 12894
rect 3754 12830 3771 12894
rect 3835 12830 3852 12894
rect 3916 12830 3933 12894
rect 3997 12830 4014 12894
rect 4078 12830 4095 12894
rect 4159 12830 4176 12894
rect 4240 12830 4257 12894
rect 4321 12830 4338 12894
rect 4402 12830 4420 12894
rect 4484 12830 4502 12894
rect 4566 12830 4584 12894
rect 4648 12830 4666 12894
rect 4730 12830 4748 12894
rect 4812 12830 4830 12894
rect 4894 12830 4895 12894
rect 0 12812 4895 12830
rect 0 12748 126 12812
rect 190 12748 207 12812
rect 271 12748 288 12812
rect 352 12748 369 12812
rect 433 12748 450 12812
rect 514 12748 531 12812
rect 595 12748 612 12812
rect 676 12748 693 12812
rect 757 12748 774 12812
rect 838 12748 855 12812
rect 919 12748 936 12812
rect 1000 12748 1017 12812
rect 1081 12748 1098 12812
rect 1162 12748 1179 12812
rect 1243 12748 1260 12812
rect 1324 12748 1341 12812
rect 1405 12748 1422 12812
rect 1486 12748 1503 12812
rect 1567 12748 1584 12812
rect 1648 12748 1665 12812
rect 1729 12748 1746 12812
rect 1810 12748 1827 12812
rect 1891 12748 1908 12812
rect 1972 12748 1989 12812
rect 2053 12748 2070 12812
rect 2134 12748 2151 12812
rect 2215 12748 2232 12812
rect 2296 12748 2313 12812
rect 2377 12748 2394 12812
rect 2458 12748 2475 12812
rect 2539 12748 2556 12812
rect 2620 12748 2637 12812
rect 2701 12748 2718 12812
rect 2782 12748 2799 12812
rect 2863 12748 2880 12812
rect 2944 12748 2961 12812
rect 3025 12748 3042 12812
rect 3106 12748 3123 12812
rect 3187 12748 3204 12812
rect 3268 12748 3285 12812
rect 3349 12748 3366 12812
rect 3430 12748 3447 12812
rect 3511 12748 3528 12812
rect 3592 12748 3609 12812
rect 3673 12748 3690 12812
rect 3754 12748 3771 12812
rect 3835 12748 3852 12812
rect 3916 12748 3933 12812
rect 3997 12748 4014 12812
rect 4078 12748 4095 12812
rect 4159 12748 4176 12812
rect 4240 12748 4257 12812
rect 4321 12748 4338 12812
rect 4402 12748 4420 12812
rect 4484 12748 4502 12812
rect 4566 12748 4584 12812
rect 4648 12748 4666 12812
rect 4730 12748 4748 12812
rect 4812 12748 4830 12812
rect 4894 12748 4895 12812
rect 0 12730 4895 12748
rect 0 12666 126 12730
rect 190 12666 207 12730
rect 271 12666 288 12730
rect 352 12666 369 12730
rect 433 12666 450 12730
rect 514 12666 531 12730
rect 595 12666 612 12730
rect 676 12666 693 12730
rect 757 12666 774 12730
rect 838 12666 855 12730
rect 919 12666 936 12730
rect 1000 12666 1017 12730
rect 1081 12666 1098 12730
rect 1162 12666 1179 12730
rect 1243 12666 1260 12730
rect 1324 12666 1341 12730
rect 1405 12666 1422 12730
rect 1486 12666 1503 12730
rect 1567 12666 1584 12730
rect 1648 12666 1665 12730
rect 1729 12666 1746 12730
rect 1810 12666 1827 12730
rect 1891 12666 1908 12730
rect 1972 12666 1989 12730
rect 2053 12666 2070 12730
rect 2134 12666 2151 12730
rect 2215 12666 2232 12730
rect 2296 12666 2313 12730
rect 2377 12666 2394 12730
rect 2458 12666 2475 12730
rect 2539 12666 2556 12730
rect 2620 12666 2637 12730
rect 2701 12666 2718 12730
rect 2782 12666 2799 12730
rect 2863 12666 2880 12730
rect 2944 12666 2961 12730
rect 3025 12666 3042 12730
rect 3106 12666 3123 12730
rect 3187 12666 3204 12730
rect 3268 12666 3285 12730
rect 3349 12666 3366 12730
rect 3430 12666 3447 12730
rect 3511 12666 3528 12730
rect 3592 12666 3609 12730
rect 3673 12666 3690 12730
rect 3754 12666 3771 12730
rect 3835 12666 3852 12730
rect 3916 12666 3933 12730
rect 3997 12666 4014 12730
rect 4078 12666 4095 12730
rect 4159 12666 4176 12730
rect 4240 12666 4257 12730
rect 4321 12666 4338 12730
rect 4402 12666 4420 12730
rect 4484 12666 4502 12730
rect 4566 12666 4584 12730
rect 4648 12666 4666 12730
rect 4730 12666 4748 12730
rect 4812 12666 4830 12730
rect 4894 12666 4895 12730
rect 0 12648 4895 12666
rect 0 12584 126 12648
rect 190 12584 207 12648
rect 271 12584 288 12648
rect 352 12584 369 12648
rect 433 12584 450 12648
rect 514 12584 531 12648
rect 595 12584 612 12648
rect 676 12584 693 12648
rect 757 12584 774 12648
rect 838 12584 855 12648
rect 919 12584 936 12648
rect 1000 12584 1017 12648
rect 1081 12584 1098 12648
rect 1162 12584 1179 12648
rect 1243 12584 1260 12648
rect 1324 12584 1341 12648
rect 1405 12584 1422 12648
rect 1486 12584 1503 12648
rect 1567 12584 1584 12648
rect 1648 12584 1665 12648
rect 1729 12584 1746 12648
rect 1810 12584 1827 12648
rect 1891 12584 1908 12648
rect 1972 12584 1989 12648
rect 2053 12584 2070 12648
rect 2134 12584 2151 12648
rect 2215 12584 2232 12648
rect 2296 12584 2313 12648
rect 2377 12584 2394 12648
rect 2458 12584 2475 12648
rect 2539 12584 2556 12648
rect 2620 12584 2637 12648
rect 2701 12584 2718 12648
rect 2782 12584 2799 12648
rect 2863 12584 2880 12648
rect 2944 12584 2961 12648
rect 3025 12584 3042 12648
rect 3106 12584 3123 12648
rect 3187 12584 3204 12648
rect 3268 12584 3285 12648
rect 3349 12584 3366 12648
rect 3430 12584 3447 12648
rect 3511 12584 3528 12648
rect 3592 12584 3609 12648
rect 3673 12584 3690 12648
rect 3754 12584 3771 12648
rect 3835 12584 3852 12648
rect 3916 12584 3933 12648
rect 3997 12584 4014 12648
rect 4078 12584 4095 12648
rect 4159 12584 4176 12648
rect 4240 12584 4257 12648
rect 4321 12584 4338 12648
rect 4402 12584 4420 12648
rect 4484 12584 4502 12648
rect 4566 12584 4584 12648
rect 4648 12584 4666 12648
rect 4730 12584 4748 12648
rect 4812 12584 4830 12648
rect 4894 12584 4895 12648
rect 0 12566 4895 12584
rect 0 12502 126 12566
rect 190 12502 207 12566
rect 271 12502 288 12566
rect 352 12502 369 12566
rect 433 12502 450 12566
rect 514 12502 531 12566
rect 595 12502 612 12566
rect 676 12502 693 12566
rect 757 12502 774 12566
rect 838 12502 855 12566
rect 919 12502 936 12566
rect 1000 12502 1017 12566
rect 1081 12502 1098 12566
rect 1162 12502 1179 12566
rect 1243 12502 1260 12566
rect 1324 12502 1341 12566
rect 1405 12502 1422 12566
rect 1486 12502 1503 12566
rect 1567 12502 1584 12566
rect 1648 12502 1665 12566
rect 1729 12502 1746 12566
rect 1810 12502 1827 12566
rect 1891 12502 1908 12566
rect 1972 12502 1989 12566
rect 2053 12502 2070 12566
rect 2134 12502 2151 12566
rect 2215 12502 2232 12566
rect 2296 12502 2313 12566
rect 2377 12502 2394 12566
rect 2458 12502 2475 12566
rect 2539 12502 2556 12566
rect 2620 12502 2637 12566
rect 2701 12502 2718 12566
rect 2782 12502 2799 12566
rect 2863 12502 2880 12566
rect 2944 12502 2961 12566
rect 3025 12502 3042 12566
rect 3106 12502 3123 12566
rect 3187 12502 3204 12566
rect 3268 12502 3285 12566
rect 3349 12502 3366 12566
rect 3430 12502 3447 12566
rect 3511 12502 3528 12566
rect 3592 12502 3609 12566
rect 3673 12502 3690 12566
rect 3754 12502 3771 12566
rect 3835 12502 3852 12566
rect 3916 12502 3933 12566
rect 3997 12502 4014 12566
rect 4078 12502 4095 12566
rect 4159 12502 4176 12566
rect 4240 12502 4257 12566
rect 4321 12502 4338 12566
rect 4402 12502 4420 12566
rect 4484 12502 4502 12566
rect 4566 12502 4584 12566
rect 4648 12502 4666 12566
rect 4730 12502 4748 12566
rect 4812 12502 4830 12566
rect 4894 12502 4895 12566
rect 0 12484 4895 12502
rect 0 12420 126 12484
rect 190 12420 207 12484
rect 271 12420 288 12484
rect 352 12420 369 12484
rect 433 12420 450 12484
rect 514 12420 531 12484
rect 595 12420 612 12484
rect 676 12420 693 12484
rect 757 12420 774 12484
rect 838 12420 855 12484
rect 919 12420 936 12484
rect 1000 12420 1017 12484
rect 1081 12420 1098 12484
rect 1162 12420 1179 12484
rect 1243 12420 1260 12484
rect 1324 12420 1341 12484
rect 1405 12420 1422 12484
rect 1486 12420 1503 12484
rect 1567 12420 1584 12484
rect 1648 12420 1665 12484
rect 1729 12420 1746 12484
rect 1810 12420 1827 12484
rect 1891 12420 1908 12484
rect 1972 12420 1989 12484
rect 2053 12420 2070 12484
rect 2134 12420 2151 12484
rect 2215 12420 2232 12484
rect 2296 12420 2313 12484
rect 2377 12420 2394 12484
rect 2458 12420 2475 12484
rect 2539 12420 2556 12484
rect 2620 12420 2637 12484
rect 2701 12420 2718 12484
rect 2782 12420 2799 12484
rect 2863 12420 2880 12484
rect 2944 12420 2961 12484
rect 3025 12420 3042 12484
rect 3106 12420 3123 12484
rect 3187 12420 3204 12484
rect 3268 12420 3285 12484
rect 3349 12420 3366 12484
rect 3430 12420 3447 12484
rect 3511 12420 3528 12484
rect 3592 12420 3609 12484
rect 3673 12420 3690 12484
rect 3754 12420 3771 12484
rect 3835 12420 3852 12484
rect 3916 12420 3933 12484
rect 3997 12420 4014 12484
rect 4078 12420 4095 12484
rect 4159 12420 4176 12484
rect 4240 12420 4257 12484
rect 4321 12420 4338 12484
rect 4402 12420 4420 12484
rect 4484 12420 4502 12484
rect 4566 12420 4584 12484
rect 4648 12420 4666 12484
rect 4730 12420 4748 12484
rect 4812 12420 4830 12484
rect 4894 12420 4895 12484
rect 0 12417 4895 12420
rect 10156 13304 15000 13307
rect 10156 13240 10157 13304
rect 10221 13240 10238 13304
rect 10302 13240 10319 13304
rect 10383 13240 10400 13304
rect 10464 13240 10481 13304
rect 10545 13240 10562 13304
rect 10626 13240 10643 13304
rect 10707 13240 10724 13304
rect 10788 13240 10805 13304
rect 10869 13240 10886 13304
rect 10950 13240 10967 13304
rect 11031 13240 11048 13304
rect 11112 13240 11129 13304
rect 11193 13240 11210 13304
rect 11274 13240 11291 13304
rect 11355 13240 11372 13304
rect 11436 13240 11453 13304
rect 11517 13240 11534 13304
rect 11598 13240 11615 13304
rect 11679 13240 11696 13304
rect 11760 13240 11777 13304
rect 11841 13240 11858 13304
rect 11922 13240 11939 13304
rect 12003 13240 12020 13304
rect 12084 13240 12101 13304
rect 12165 13240 12182 13304
rect 12246 13240 12263 13304
rect 12327 13240 12344 13304
rect 12408 13240 12425 13304
rect 12489 13240 12506 13304
rect 12570 13240 12587 13304
rect 12651 13240 12668 13304
rect 12732 13240 12749 13304
rect 12813 13240 12830 13304
rect 12894 13240 12911 13304
rect 12975 13240 12992 13304
rect 13056 13240 13073 13304
rect 13137 13240 13154 13304
rect 13218 13240 13235 13304
rect 13299 13240 13316 13304
rect 13380 13240 13397 13304
rect 13461 13240 13478 13304
rect 13542 13240 13559 13304
rect 13623 13240 13640 13304
rect 13704 13240 13721 13304
rect 13785 13240 13802 13304
rect 13866 13240 13883 13304
rect 13947 13240 13964 13304
rect 14028 13240 14045 13304
rect 14109 13240 14126 13304
rect 14190 13240 14207 13304
rect 14271 13240 14288 13304
rect 14352 13240 14369 13304
rect 14433 13240 14451 13304
rect 14515 13240 14533 13304
rect 14597 13240 14615 13304
rect 14679 13240 14697 13304
rect 14761 13240 14779 13304
rect 14843 13240 14861 13304
rect 14925 13240 15000 13304
rect 10156 13222 15000 13240
rect 10156 13158 10157 13222
rect 10221 13158 10238 13222
rect 10302 13158 10319 13222
rect 10383 13158 10400 13222
rect 10464 13158 10481 13222
rect 10545 13158 10562 13222
rect 10626 13158 10643 13222
rect 10707 13158 10724 13222
rect 10788 13158 10805 13222
rect 10869 13158 10886 13222
rect 10950 13158 10967 13222
rect 11031 13158 11048 13222
rect 11112 13158 11129 13222
rect 11193 13158 11210 13222
rect 11274 13158 11291 13222
rect 11355 13158 11372 13222
rect 11436 13158 11453 13222
rect 11517 13158 11534 13222
rect 11598 13158 11615 13222
rect 11679 13158 11696 13222
rect 11760 13158 11777 13222
rect 11841 13158 11858 13222
rect 11922 13158 11939 13222
rect 12003 13158 12020 13222
rect 12084 13158 12101 13222
rect 12165 13158 12182 13222
rect 12246 13158 12263 13222
rect 12327 13158 12344 13222
rect 12408 13158 12425 13222
rect 12489 13158 12506 13222
rect 12570 13158 12587 13222
rect 12651 13158 12668 13222
rect 12732 13158 12749 13222
rect 12813 13158 12830 13222
rect 12894 13158 12911 13222
rect 12975 13158 12992 13222
rect 13056 13158 13073 13222
rect 13137 13158 13154 13222
rect 13218 13158 13235 13222
rect 13299 13158 13316 13222
rect 13380 13158 13397 13222
rect 13461 13158 13478 13222
rect 13542 13158 13559 13222
rect 13623 13158 13640 13222
rect 13704 13158 13721 13222
rect 13785 13158 13802 13222
rect 13866 13158 13883 13222
rect 13947 13158 13964 13222
rect 14028 13158 14045 13222
rect 14109 13158 14126 13222
rect 14190 13158 14207 13222
rect 14271 13158 14288 13222
rect 14352 13158 14369 13222
rect 14433 13158 14451 13222
rect 14515 13158 14533 13222
rect 14597 13158 14615 13222
rect 14679 13158 14697 13222
rect 14761 13158 14779 13222
rect 14843 13158 14861 13222
rect 14925 13158 15000 13222
rect 10156 13140 15000 13158
rect 10156 13076 10157 13140
rect 10221 13076 10238 13140
rect 10302 13076 10319 13140
rect 10383 13076 10400 13140
rect 10464 13076 10481 13140
rect 10545 13076 10562 13140
rect 10626 13076 10643 13140
rect 10707 13076 10724 13140
rect 10788 13076 10805 13140
rect 10869 13076 10886 13140
rect 10950 13076 10967 13140
rect 11031 13076 11048 13140
rect 11112 13076 11129 13140
rect 11193 13076 11210 13140
rect 11274 13076 11291 13140
rect 11355 13076 11372 13140
rect 11436 13076 11453 13140
rect 11517 13076 11534 13140
rect 11598 13076 11615 13140
rect 11679 13076 11696 13140
rect 11760 13076 11777 13140
rect 11841 13076 11858 13140
rect 11922 13076 11939 13140
rect 12003 13076 12020 13140
rect 12084 13076 12101 13140
rect 12165 13076 12182 13140
rect 12246 13076 12263 13140
rect 12327 13076 12344 13140
rect 12408 13076 12425 13140
rect 12489 13076 12506 13140
rect 12570 13076 12587 13140
rect 12651 13076 12668 13140
rect 12732 13076 12749 13140
rect 12813 13076 12830 13140
rect 12894 13076 12911 13140
rect 12975 13076 12992 13140
rect 13056 13076 13073 13140
rect 13137 13076 13154 13140
rect 13218 13076 13235 13140
rect 13299 13076 13316 13140
rect 13380 13076 13397 13140
rect 13461 13076 13478 13140
rect 13542 13076 13559 13140
rect 13623 13076 13640 13140
rect 13704 13076 13721 13140
rect 13785 13076 13802 13140
rect 13866 13076 13883 13140
rect 13947 13076 13964 13140
rect 14028 13076 14045 13140
rect 14109 13076 14126 13140
rect 14190 13076 14207 13140
rect 14271 13076 14288 13140
rect 14352 13076 14369 13140
rect 14433 13076 14451 13140
rect 14515 13076 14533 13140
rect 14597 13076 14615 13140
rect 14679 13076 14697 13140
rect 14761 13076 14779 13140
rect 14843 13076 14861 13140
rect 14925 13076 15000 13140
rect 10156 13058 15000 13076
rect 10156 12994 10157 13058
rect 10221 12994 10238 13058
rect 10302 12994 10319 13058
rect 10383 12994 10400 13058
rect 10464 12994 10481 13058
rect 10545 12994 10562 13058
rect 10626 12994 10643 13058
rect 10707 12994 10724 13058
rect 10788 12994 10805 13058
rect 10869 12994 10886 13058
rect 10950 12994 10967 13058
rect 11031 12994 11048 13058
rect 11112 12994 11129 13058
rect 11193 12994 11210 13058
rect 11274 12994 11291 13058
rect 11355 12994 11372 13058
rect 11436 12994 11453 13058
rect 11517 12994 11534 13058
rect 11598 12994 11615 13058
rect 11679 12994 11696 13058
rect 11760 12994 11777 13058
rect 11841 12994 11858 13058
rect 11922 12994 11939 13058
rect 12003 12994 12020 13058
rect 12084 12994 12101 13058
rect 12165 12994 12182 13058
rect 12246 12994 12263 13058
rect 12327 12994 12344 13058
rect 12408 12994 12425 13058
rect 12489 12994 12506 13058
rect 12570 12994 12587 13058
rect 12651 12994 12668 13058
rect 12732 12994 12749 13058
rect 12813 12994 12830 13058
rect 12894 12994 12911 13058
rect 12975 12994 12992 13058
rect 13056 12994 13073 13058
rect 13137 12994 13154 13058
rect 13218 12994 13235 13058
rect 13299 12994 13316 13058
rect 13380 12994 13397 13058
rect 13461 12994 13478 13058
rect 13542 12994 13559 13058
rect 13623 12994 13640 13058
rect 13704 12994 13721 13058
rect 13785 12994 13802 13058
rect 13866 12994 13883 13058
rect 13947 12994 13964 13058
rect 14028 12994 14045 13058
rect 14109 12994 14126 13058
rect 14190 12994 14207 13058
rect 14271 12994 14288 13058
rect 14352 12994 14369 13058
rect 14433 12994 14451 13058
rect 14515 12994 14533 13058
rect 14597 12994 14615 13058
rect 14679 12994 14697 13058
rect 14761 12994 14779 13058
rect 14843 12994 14861 13058
rect 14925 12994 15000 13058
rect 10156 12976 15000 12994
rect 10156 12912 10157 12976
rect 10221 12912 10238 12976
rect 10302 12912 10319 12976
rect 10383 12912 10400 12976
rect 10464 12912 10481 12976
rect 10545 12912 10562 12976
rect 10626 12912 10643 12976
rect 10707 12912 10724 12976
rect 10788 12912 10805 12976
rect 10869 12912 10886 12976
rect 10950 12912 10967 12976
rect 11031 12912 11048 12976
rect 11112 12912 11129 12976
rect 11193 12912 11210 12976
rect 11274 12912 11291 12976
rect 11355 12912 11372 12976
rect 11436 12912 11453 12976
rect 11517 12912 11534 12976
rect 11598 12912 11615 12976
rect 11679 12912 11696 12976
rect 11760 12912 11777 12976
rect 11841 12912 11858 12976
rect 11922 12912 11939 12976
rect 12003 12912 12020 12976
rect 12084 12912 12101 12976
rect 12165 12912 12182 12976
rect 12246 12912 12263 12976
rect 12327 12912 12344 12976
rect 12408 12912 12425 12976
rect 12489 12912 12506 12976
rect 12570 12912 12587 12976
rect 12651 12912 12668 12976
rect 12732 12912 12749 12976
rect 12813 12912 12830 12976
rect 12894 12912 12911 12976
rect 12975 12912 12992 12976
rect 13056 12912 13073 12976
rect 13137 12912 13154 12976
rect 13218 12912 13235 12976
rect 13299 12912 13316 12976
rect 13380 12912 13397 12976
rect 13461 12912 13478 12976
rect 13542 12912 13559 12976
rect 13623 12912 13640 12976
rect 13704 12912 13721 12976
rect 13785 12912 13802 12976
rect 13866 12912 13883 12976
rect 13947 12912 13964 12976
rect 14028 12912 14045 12976
rect 14109 12912 14126 12976
rect 14190 12912 14207 12976
rect 14271 12912 14288 12976
rect 14352 12912 14369 12976
rect 14433 12912 14451 12976
rect 14515 12912 14533 12976
rect 14597 12912 14615 12976
rect 14679 12912 14697 12976
rect 14761 12912 14779 12976
rect 14843 12912 14861 12976
rect 14925 12912 15000 12976
rect 10156 12894 15000 12912
rect 10156 12830 10157 12894
rect 10221 12830 10238 12894
rect 10302 12830 10319 12894
rect 10383 12830 10400 12894
rect 10464 12830 10481 12894
rect 10545 12830 10562 12894
rect 10626 12830 10643 12894
rect 10707 12830 10724 12894
rect 10788 12830 10805 12894
rect 10869 12830 10886 12894
rect 10950 12830 10967 12894
rect 11031 12830 11048 12894
rect 11112 12830 11129 12894
rect 11193 12830 11210 12894
rect 11274 12830 11291 12894
rect 11355 12830 11372 12894
rect 11436 12830 11453 12894
rect 11517 12830 11534 12894
rect 11598 12830 11615 12894
rect 11679 12830 11696 12894
rect 11760 12830 11777 12894
rect 11841 12830 11858 12894
rect 11922 12830 11939 12894
rect 12003 12830 12020 12894
rect 12084 12830 12101 12894
rect 12165 12830 12182 12894
rect 12246 12830 12263 12894
rect 12327 12830 12344 12894
rect 12408 12830 12425 12894
rect 12489 12830 12506 12894
rect 12570 12830 12587 12894
rect 12651 12830 12668 12894
rect 12732 12830 12749 12894
rect 12813 12830 12830 12894
rect 12894 12830 12911 12894
rect 12975 12830 12992 12894
rect 13056 12830 13073 12894
rect 13137 12830 13154 12894
rect 13218 12830 13235 12894
rect 13299 12830 13316 12894
rect 13380 12830 13397 12894
rect 13461 12830 13478 12894
rect 13542 12830 13559 12894
rect 13623 12830 13640 12894
rect 13704 12830 13721 12894
rect 13785 12830 13802 12894
rect 13866 12830 13883 12894
rect 13947 12830 13964 12894
rect 14028 12830 14045 12894
rect 14109 12830 14126 12894
rect 14190 12830 14207 12894
rect 14271 12830 14288 12894
rect 14352 12830 14369 12894
rect 14433 12830 14451 12894
rect 14515 12830 14533 12894
rect 14597 12830 14615 12894
rect 14679 12830 14697 12894
rect 14761 12830 14779 12894
rect 14843 12830 14861 12894
rect 14925 12830 15000 12894
rect 10156 12812 15000 12830
rect 10156 12748 10157 12812
rect 10221 12748 10238 12812
rect 10302 12748 10319 12812
rect 10383 12748 10400 12812
rect 10464 12748 10481 12812
rect 10545 12748 10562 12812
rect 10626 12748 10643 12812
rect 10707 12748 10724 12812
rect 10788 12748 10805 12812
rect 10869 12748 10886 12812
rect 10950 12748 10967 12812
rect 11031 12748 11048 12812
rect 11112 12748 11129 12812
rect 11193 12748 11210 12812
rect 11274 12748 11291 12812
rect 11355 12748 11372 12812
rect 11436 12748 11453 12812
rect 11517 12748 11534 12812
rect 11598 12748 11615 12812
rect 11679 12748 11696 12812
rect 11760 12748 11777 12812
rect 11841 12748 11858 12812
rect 11922 12748 11939 12812
rect 12003 12748 12020 12812
rect 12084 12748 12101 12812
rect 12165 12748 12182 12812
rect 12246 12748 12263 12812
rect 12327 12748 12344 12812
rect 12408 12748 12425 12812
rect 12489 12748 12506 12812
rect 12570 12748 12587 12812
rect 12651 12748 12668 12812
rect 12732 12748 12749 12812
rect 12813 12748 12830 12812
rect 12894 12748 12911 12812
rect 12975 12748 12992 12812
rect 13056 12748 13073 12812
rect 13137 12748 13154 12812
rect 13218 12748 13235 12812
rect 13299 12748 13316 12812
rect 13380 12748 13397 12812
rect 13461 12748 13478 12812
rect 13542 12748 13559 12812
rect 13623 12748 13640 12812
rect 13704 12748 13721 12812
rect 13785 12748 13802 12812
rect 13866 12748 13883 12812
rect 13947 12748 13964 12812
rect 14028 12748 14045 12812
rect 14109 12748 14126 12812
rect 14190 12748 14207 12812
rect 14271 12748 14288 12812
rect 14352 12748 14369 12812
rect 14433 12748 14451 12812
rect 14515 12748 14533 12812
rect 14597 12748 14615 12812
rect 14679 12748 14697 12812
rect 14761 12748 14779 12812
rect 14843 12748 14861 12812
rect 14925 12748 15000 12812
rect 10156 12730 15000 12748
rect 10156 12666 10157 12730
rect 10221 12666 10238 12730
rect 10302 12666 10319 12730
rect 10383 12666 10400 12730
rect 10464 12666 10481 12730
rect 10545 12666 10562 12730
rect 10626 12666 10643 12730
rect 10707 12666 10724 12730
rect 10788 12666 10805 12730
rect 10869 12666 10886 12730
rect 10950 12666 10967 12730
rect 11031 12666 11048 12730
rect 11112 12666 11129 12730
rect 11193 12666 11210 12730
rect 11274 12666 11291 12730
rect 11355 12666 11372 12730
rect 11436 12666 11453 12730
rect 11517 12666 11534 12730
rect 11598 12666 11615 12730
rect 11679 12666 11696 12730
rect 11760 12666 11777 12730
rect 11841 12666 11858 12730
rect 11922 12666 11939 12730
rect 12003 12666 12020 12730
rect 12084 12666 12101 12730
rect 12165 12666 12182 12730
rect 12246 12666 12263 12730
rect 12327 12666 12344 12730
rect 12408 12666 12425 12730
rect 12489 12666 12506 12730
rect 12570 12666 12587 12730
rect 12651 12666 12668 12730
rect 12732 12666 12749 12730
rect 12813 12666 12830 12730
rect 12894 12666 12911 12730
rect 12975 12666 12992 12730
rect 13056 12666 13073 12730
rect 13137 12666 13154 12730
rect 13218 12666 13235 12730
rect 13299 12666 13316 12730
rect 13380 12666 13397 12730
rect 13461 12666 13478 12730
rect 13542 12666 13559 12730
rect 13623 12666 13640 12730
rect 13704 12666 13721 12730
rect 13785 12666 13802 12730
rect 13866 12666 13883 12730
rect 13947 12666 13964 12730
rect 14028 12666 14045 12730
rect 14109 12666 14126 12730
rect 14190 12666 14207 12730
rect 14271 12666 14288 12730
rect 14352 12666 14369 12730
rect 14433 12666 14451 12730
rect 14515 12666 14533 12730
rect 14597 12666 14615 12730
rect 14679 12666 14697 12730
rect 14761 12666 14779 12730
rect 14843 12666 14861 12730
rect 14925 12666 15000 12730
rect 10156 12648 15000 12666
rect 10156 12584 10157 12648
rect 10221 12584 10238 12648
rect 10302 12584 10319 12648
rect 10383 12584 10400 12648
rect 10464 12584 10481 12648
rect 10545 12584 10562 12648
rect 10626 12584 10643 12648
rect 10707 12584 10724 12648
rect 10788 12584 10805 12648
rect 10869 12584 10886 12648
rect 10950 12584 10967 12648
rect 11031 12584 11048 12648
rect 11112 12584 11129 12648
rect 11193 12584 11210 12648
rect 11274 12584 11291 12648
rect 11355 12584 11372 12648
rect 11436 12584 11453 12648
rect 11517 12584 11534 12648
rect 11598 12584 11615 12648
rect 11679 12584 11696 12648
rect 11760 12584 11777 12648
rect 11841 12584 11858 12648
rect 11922 12584 11939 12648
rect 12003 12584 12020 12648
rect 12084 12584 12101 12648
rect 12165 12584 12182 12648
rect 12246 12584 12263 12648
rect 12327 12584 12344 12648
rect 12408 12584 12425 12648
rect 12489 12584 12506 12648
rect 12570 12584 12587 12648
rect 12651 12584 12668 12648
rect 12732 12584 12749 12648
rect 12813 12584 12830 12648
rect 12894 12584 12911 12648
rect 12975 12584 12992 12648
rect 13056 12584 13073 12648
rect 13137 12584 13154 12648
rect 13218 12584 13235 12648
rect 13299 12584 13316 12648
rect 13380 12584 13397 12648
rect 13461 12584 13478 12648
rect 13542 12584 13559 12648
rect 13623 12584 13640 12648
rect 13704 12584 13721 12648
rect 13785 12584 13802 12648
rect 13866 12584 13883 12648
rect 13947 12584 13964 12648
rect 14028 12584 14045 12648
rect 14109 12584 14126 12648
rect 14190 12584 14207 12648
rect 14271 12584 14288 12648
rect 14352 12584 14369 12648
rect 14433 12584 14451 12648
rect 14515 12584 14533 12648
rect 14597 12584 14615 12648
rect 14679 12584 14697 12648
rect 14761 12584 14779 12648
rect 14843 12584 14861 12648
rect 14925 12584 15000 12648
rect 10156 12566 15000 12584
rect 10156 12502 10157 12566
rect 10221 12502 10238 12566
rect 10302 12502 10319 12566
rect 10383 12502 10400 12566
rect 10464 12502 10481 12566
rect 10545 12502 10562 12566
rect 10626 12502 10643 12566
rect 10707 12502 10724 12566
rect 10788 12502 10805 12566
rect 10869 12502 10886 12566
rect 10950 12502 10967 12566
rect 11031 12502 11048 12566
rect 11112 12502 11129 12566
rect 11193 12502 11210 12566
rect 11274 12502 11291 12566
rect 11355 12502 11372 12566
rect 11436 12502 11453 12566
rect 11517 12502 11534 12566
rect 11598 12502 11615 12566
rect 11679 12502 11696 12566
rect 11760 12502 11777 12566
rect 11841 12502 11858 12566
rect 11922 12502 11939 12566
rect 12003 12502 12020 12566
rect 12084 12502 12101 12566
rect 12165 12502 12182 12566
rect 12246 12502 12263 12566
rect 12327 12502 12344 12566
rect 12408 12502 12425 12566
rect 12489 12502 12506 12566
rect 12570 12502 12587 12566
rect 12651 12502 12668 12566
rect 12732 12502 12749 12566
rect 12813 12502 12830 12566
rect 12894 12502 12911 12566
rect 12975 12502 12992 12566
rect 13056 12502 13073 12566
rect 13137 12502 13154 12566
rect 13218 12502 13235 12566
rect 13299 12502 13316 12566
rect 13380 12502 13397 12566
rect 13461 12502 13478 12566
rect 13542 12502 13559 12566
rect 13623 12502 13640 12566
rect 13704 12502 13721 12566
rect 13785 12502 13802 12566
rect 13866 12502 13883 12566
rect 13947 12502 13964 12566
rect 14028 12502 14045 12566
rect 14109 12502 14126 12566
rect 14190 12502 14207 12566
rect 14271 12502 14288 12566
rect 14352 12502 14369 12566
rect 14433 12502 14451 12566
rect 14515 12502 14533 12566
rect 14597 12502 14615 12566
rect 14679 12502 14697 12566
rect 14761 12502 14779 12566
rect 14843 12502 14861 12566
rect 14925 12502 15000 12566
rect 10156 12484 15000 12502
rect 10156 12420 10157 12484
rect 10221 12420 10238 12484
rect 10302 12420 10319 12484
rect 10383 12420 10400 12484
rect 10464 12420 10481 12484
rect 10545 12420 10562 12484
rect 10626 12420 10643 12484
rect 10707 12420 10724 12484
rect 10788 12420 10805 12484
rect 10869 12420 10886 12484
rect 10950 12420 10967 12484
rect 11031 12420 11048 12484
rect 11112 12420 11129 12484
rect 11193 12420 11210 12484
rect 11274 12420 11291 12484
rect 11355 12420 11372 12484
rect 11436 12420 11453 12484
rect 11517 12420 11534 12484
rect 11598 12420 11615 12484
rect 11679 12420 11696 12484
rect 11760 12420 11777 12484
rect 11841 12420 11858 12484
rect 11922 12420 11939 12484
rect 12003 12420 12020 12484
rect 12084 12420 12101 12484
rect 12165 12420 12182 12484
rect 12246 12420 12263 12484
rect 12327 12420 12344 12484
rect 12408 12420 12425 12484
rect 12489 12420 12506 12484
rect 12570 12420 12587 12484
rect 12651 12420 12668 12484
rect 12732 12420 12749 12484
rect 12813 12420 12830 12484
rect 12894 12420 12911 12484
rect 12975 12420 12992 12484
rect 13056 12420 13073 12484
rect 13137 12420 13154 12484
rect 13218 12420 13235 12484
rect 13299 12420 13316 12484
rect 13380 12420 13397 12484
rect 13461 12420 13478 12484
rect 13542 12420 13559 12484
rect 13623 12420 13640 12484
rect 13704 12420 13721 12484
rect 13785 12420 13802 12484
rect 13866 12420 13883 12484
rect 13947 12420 13964 12484
rect 14028 12420 14045 12484
rect 14109 12420 14126 12484
rect 14190 12420 14207 12484
rect 14271 12420 14288 12484
rect 14352 12420 14369 12484
rect 14433 12420 14451 12484
rect 14515 12420 14533 12484
rect 14597 12420 14615 12484
rect 14679 12420 14697 12484
rect 14761 12420 14779 12484
rect 14843 12420 14861 12484
rect 14925 12420 15000 12484
rect 10156 12417 15000 12420
rect 0 11247 254 12137
rect 14746 11247 15000 12137
rect 0 10881 254 10947
rect 14746 10881 15000 10947
rect 0 10225 254 10821
rect 14746 10225 15000 10821
rect 0 9929 254 10165
rect 14746 9929 15000 10165
rect 0 9273 254 9869
rect 14746 9273 15000 9869
rect 0 9147 254 9213
rect 14746 9147 15000 9213
rect 0 7917 254 8847
rect 14746 7917 15000 8847
rect 0 6947 254 7637
rect 14746 6947 15000 7637
rect 0 5977 254 6667
rect 14746 5977 15000 6667
rect 0 4767 254 5697
rect 14746 4767 15000 5697
rect 0 4484 4895 4487
rect 0 4420 126 4484
rect 190 4420 207 4484
rect 271 4420 288 4484
rect 352 4420 369 4484
rect 433 4420 450 4484
rect 514 4420 531 4484
rect 595 4420 612 4484
rect 676 4420 693 4484
rect 757 4420 774 4484
rect 838 4420 855 4484
rect 919 4420 936 4484
rect 1000 4420 1017 4484
rect 1081 4420 1098 4484
rect 1162 4420 1179 4484
rect 1243 4420 1260 4484
rect 1324 4420 1341 4484
rect 1405 4420 1422 4484
rect 1486 4420 1503 4484
rect 1567 4420 1584 4484
rect 1648 4420 1665 4484
rect 1729 4420 1746 4484
rect 1810 4420 1827 4484
rect 1891 4420 1908 4484
rect 1972 4420 1989 4484
rect 2053 4420 2070 4484
rect 2134 4420 2151 4484
rect 2215 4420 2232 4484
rect 2296 4420 2313 4484
rect 2377 4420 2394 4484
rect 2458 4420 2475 4484
rect 2539 4420 2556 4484
rect 2620 4420 2637 4484
rect 2701 4420 2718 4484
rect 2782 4420 2799 4484
rect 2863 4420 2880 4484
rect 2944 4420 2961 4484
rect 3025 4420 3042 4484
rect 3106 4420 3123 4484
rect 3187 4420 3204 4484
rect 3268 4420 3285 4484
rect 3349 4420 3366 4484
rect 3430 4420 3447 4484
rect 3511 4420 3528 4484
rect 3592 4420 3609 4484
rect 3673 4420 3690 4484
rect 3754 4420 3771 4484
rect 3835 4420 3852 4484
rect 3916 4420 3933 4484
rect 3997 4420 4014 4484
rect 4078 4420 4095 4484
rect 4159 4420 4176 4484
rect 4240 4420 4257 4484
rect 4321 4420 4338 4484
rect 4402 4420 4420 4484
rect 4484 4420 4502 4484
rect 4566 4420 4584 4484
rect 4648 4420 4666 4484
rect 4730 4420 4748 4484
rect 4812 4420 4830 4484
rect 4894 4420 4895 4484
rect 0 4398 4895 4420
rect 0 4334 126 4398
rect 190 4334 207 4398
rect 271 4334 288 4398
rect 352 4334 369 4398
rect 433 4334 450 4398
rect 514 4334 531 4398
rect 595 4334 612 4398
rect 676 4334 693 4398
rect 757 4334 774 4398
rect 838 4334 855 4398
rect 919 4334 936 4398
rect 1000 4334 1017 4398
rect 1081 4334 1098 4398
rect 1162 4334 1179 4398
rect 1243 4334 1260 4398
rect 1324 4334 1341 4398
rect 1405 4334 1422 4398
rect 1486 4334 1503 4398
rect 1567 4334 1584 4398
rect 1648 4334 1665 4398
rect 1729 4334 1746 4398
rect 1810 4334 1827 4398
rect 1891 4334 1908 4398
rect 1972 4334 1989 4398
rect 2053 4334 2070 4398
rect 2134 4334 2151 4398
rect 2215 4334 2232 4398
rect 2296 4334 2313 4398
rect 2377 4334 2394 4398
rect 2458 4334 2475 4398
rect 2539 4334 2556 4398
rect 2620 4334 2637 4398
rect 2701 4334 2718 4398
rect 2782 4334 2799 4398
rect 2863 4334 2880 4398
rect 2944 4334 2961 4398
rect 3025 4334 3042 4398
rect 3106 4334 3123 4398
rect 3187 4334 3204 4398
rect 3268 4334 3285 4398
rect 3349 4334 3366 4398
rect 3430 4334 3447 4398
rect 3511 4334 3528 4398
rect 3592 4334 3609 4398
rect 3673 4334 3690 4398
rect 3754 4334 3771 4398
rect 3835 4334 3852 4398
rect 3916 4334 3933 4398
rect 3997 4334 4014 4398
rect 4078 4334 4095 4398
rect 4159 4334 4176 4398
rect 4240 4334 4257 4398
rect 4321 4334 4338 4398
rect 4402 4334 4420 4398
rect 4484 4334 4502 4398
rect 4566 4334 4584 4398
rect 4648 4334 4666 4398
rect 4730 4334 4748 4398
rect 4812 4334 4830 4398
rect 4894 4334 4895 4398
rect 0 4312 4895 4334
rect 0 4248 126 4312
rect 190 4248 207 4312
rect 271 4248 288 4312
rect 352 4248 369 4312
rect 433 4248 450 4312
rect 514 4248 531 4312
rect 595 4248 612 4312
rect 676 4248 693 4312
rect 757 4248 774 4312
rect 838 4248 855 4312
rect 919 4248 936 4312
rect 1000 4248 1017 4312
rect 1081 4248 1098 4312
rect 1162 4248 1179 4312
rect 1243 4248 1260 4312
rect 1324 4248 1341 4312
rect 1405 4248 1422 4312
rect 1486 4248 1503 4312
rect 1567 4248 1584 4312
rect 1648 4248 1665 4312
rect 1729 4248 1746 4312
rect 1810 4248 1827 4312
rect 1891 4248 1908 4312
rect 1972 4248 1989 4312
rect 2053 4248 2070 4312
rect 2134 4248 2151 4312
rect 2215 4248 2232 4312
rect 2296 4248 2313 4312
rect 2377 4248 2394 4312
rect 2458 4248 2475 4312
rect 2539 4248 2556 4312
rect 2620 4248 2637 4312
rect 2701 4248 2718 4312
rect 2782 4248 2799 4312
rect 2863 4248 2880 4312
rect 2944 4248 2961 4312
rect 3025 4248 3042 4312
rect 3106 4248 3123 4312
rect 3187 4248 3204 4312
rect 3268 4248 3285 4312
rect 3349 4248 3366 4312
rect 3430 4248 3447 4312
rect 3511 4248 3528 4312
rect 3592 4248 3609 4312
rect 3673 4248 3690 4312
rect 3754 4248 3771 4312
rect 3835 4248 3852 4312
rect 3916 4248 3933 4312
rect 3997 4248 4014 4312
rect 4078 4248 4095 4312
rect 4159 4248 4176 4312
rect 4240 4248 4257 4312
rect 4321 4248 4338 4312
rect 4402 4248 4420 4312
rect 4484 4248 4502 4312
rect 4566 4248 4584 4312
rect 4648 4248 4666 4312
rect 4730 4248 4748 4312
rect 4812 4248 4830 4312
rect 4894 4248 4895 4312
rect 0 4226 4895 4248
rect 0 4162 126 4226
rect 190 4162 207 4226
rect 271 4162 288 4226
rect 352 4162 369 4226
rect 433 4162 450 4226
rect 514 4162 531 4226
rect 595 4162 612 4226
rect 676 4162 693 4226
rect 757 4162 774 4226
rect 838 4162 855 4226
rect 919 4162 936 4226
rect 1000 4162 1017 4226
rect 1081 4162 1098 4226
rect 1162 4162 1179 4226
rect 1243 4162 1260 4226
rect 1324 4162 1341 4226
rect 1405 4162 1422 4226
rect 1486 4162 1503 4226
rect 1567 4162 1584 4226
rect 1648 4162 1665 4226
rect 1729 4162 1746 4226
rect 1810 4162 1827 4226
rect 1891 4162 1908 4226
rect 1972 4162 1989 4226
rect 2053 4162 2070 4226
rect 2134 4162 2151 4226
rect 2215 4162 2232 4226
rect 2296 4162 2313 4226
rect 2377 4162 2394 4226
rect 2458 4162 2475 4226
rect 2539 4162 2556 4226
rect 2620 4162 2637 4226
rect 2701 4162 2718 4226
rect 2782 4162 2799 4226
rect 2863 4162 2880 4226
rect 2944 4162 2961 4226
rect 3025 4162 3042 4226
rect 3106 4162 3123 4226
rect 3187 4162 3204 4226
rect 3268 4162 3285 4226
rect 3349 4162 3366 4226
rect 3430 4162 3447 4226
rect 3511 4162 3528 4226
rect 3592 4162 3609 4226
rect 3673 4162 3690 4226
rect 3754 4162 3771 4226
rect 3835 4162 3852 4226
rect 3916 4162 3933 4226
rect 3997 4162 4014 4226
rect 4078 4162 4095 4226
rect 4159 4162 4176 4226
rect 4240 4162 4257 4226
rect 4321 4162 4338 4226
rect 4402 4162 4420 4226
rect 4484 4162 4502 4226
rect 4566 4162 4584 4226
rect 4648 4162 4666 4226
rect 4730 4162 4748 4226
rect 4812 4162 4830 4226
rect 4894 4162 4895 4226
rect 0 4140 4895 4162
rect 0 4076 126 4140
rect 190 4076 207 4140
rect 271 4076 288 4140
rect 352 4076 369 4140
rect 433 4076 450 4140
rect 514 4076 531 4140
rect 595 4076 612 4140
rect 676 4076 693 4140
rect 757 4076 774 4140
rect 838 4076 855 4140
rect 919 4076 936 4140
rect 1000 4076 1017 4140
rect 1081 4076 1098 4140
rect 1162 4076 1179 4140
rect 1243 4076 1260 4140
rect 1324 4076 1341 4140
rect 1405 4076 1422 4140
rect 1486 4076 1503 4140
rect 1567 4076 1584 4140
rect 1648 4076 1665 4140
rect 1729 4076 1746 4140
rect 1810 4076 1827 4140
rect 1891 4076 1908 4140
rect 1972 4076 1989 4140
rect 2053 4076 2070 4140
rect 2134 4076 2151 4140
rect 2215 4076 2232 4140
rect 2296 4076 2313 4140
rect 2377 4076 2394 4140
rect 2458 4076 2475 4140
rect 2539 4076 2556 4140
rect 2620 4076 2637 4140
rect 2701 4076 2718 4140
rect 2782 4076 2799 4140
rect 2863 4076 2880 4140
rect 2944 4076 2961 4140
rect 3025 4076 3042 4140
rect 3106 4076 3123 4140
rect 3187 4076 3204 4140
rect 3268 4076 3285 4140
rect 3349 4076 3366 4140
rect 3430 4076 3447 4140
rect 3511 4076 3528 4140
rect 3592 4076 3609 4140
rect 3673 4076 3690 4140
rect 3754 4076 3771 4140
rect 3835 4076 3852 4140
rect 3916 4076 3933 4140
rect 3997 4076 4014 4140
rect 4078 4076 4095 4140
rect 4159 4076 4176 4140
rect 4240 4076 4257 4140
rect 4321 4076 4338 4140
rect 4402 4076 4420 4140
rect 4484 4076 4502 4140
rect 4566 4076 4584 4140
rect 4648 4076 4666 4140
rect 4730 4076 4748 4140
rect 4812 4076 4830 4140
rect 4894 4076 4895 4140
rect 0 4054 4895 4076
rect 0 3990 126 4054
rect 190 3990 207 4054
rect 271 3990 288 4054
rect 352 3990 369 4054
rect 433 3990 450 4054
rect 514 3990 531 4054
rect 595 3990 612 4054
rect 676 3990 693 4054
rect 757 3990 774 4054
rect 838 3990 855 4054
rect 919 3990 936 4054
rect 1000 3990 1017 4054
rect 1081 3990 1098 4054
rect 1162 3990 1179 4054
rect 1243 3990 1260 4054
rect 1324 3990 1341 4054
rect 1405 3990 1422 4054
rect 1486 3990 1503 4054
rect 1567 3990 1584 4054
rect 1648 3990 1665 4054
rect 1729 3990 1746 4054
rect 1810 3990 1827 4054
rect 1891 3990 1908 4054
rect 1972 3990 1989 4054
rect 2053 3990 2070 4054
rect 2134 3990 2151 4054
rect 2215 3990 2232 4054
rect 2296 3990 2313 4054
rect 2377 3990 2394 4054
rect 2458 3990 2475 4054
rect 2539 3990 2556 4054
rect 2620 3990 2637 4054
rect 2701 3990 2718 4054
rect 2782 3990 2799 4054
rect 2863 3990 2880 4054
rect 2944 3990 2961 4054
rect 3025 3990 3042 4054
rect 3106 3990 3123 4054
rect 3187 3990 3204 4054
rect 3268 3990 3285 4054
rect 3349 3990 3366 4054
rect 3430 3990 3447 4054
rect 3511 3990 3528 4054
rect 3592 3990 3609 4054
rect 3673 3990 3690 4054
rect 3754 3990 3771 4054
rect 3835 3990 3852 4054
rect 3916 3990 3933 4054
rect 3997 3990 4014 4054
rect 4078 3990 4095 4054
rect 4159 3990 4176 4054
rect 4240 3990 4257 4054
rect 4321 3990 4338 4054
rect 4402 3990 4420 4054
rect 4484 3990 4502 4054
rect 4566 3990 4584 4054
rect 4648 3990 4666 4054
rect 4730 3990 4748 4054
rect 4812 3990 4830 4054
rect 4894 3990 4895 4054
rect 0 3968 4895 3990
rect 0 3904 126 3968
rect 190 3904 207 3968
rect 271 3904 288 3968
rect 352 3904 369 3968
rect 433 3904 450 3968
rect 514 3904 531 3968
rect 595 3904 612 3968
rect 676 3904 693 3968
rect 757 3904 774 3968
rect 838 3904 855 3968
rect 919 3904 936 3968
rect 1000 3904 1017 3968
rect 1081 3904 1098 3968
rect 1162 3904 1179 3968
rect 1243 3904 1260 3968
rect 1324 3904 1341 3968
rect 1405 3904 1422 3968
rect 1486 3904 1503 3968
rect 1567 3904 1584 3968
rect 1648 3904 1665 3968
rect 1729 3904 1746 3968
rect 1810 3904 1827 3968
rect 1891 3904 1908 3968
rect 1972 3904 1989 3968
rect 2053 3904 2070 3968
rect 2134 3904 2151 3968
rect 2215 3904 2232 3968
rect 2296 3904 2313 3968
rect 2377 3904 2394 3968
rect 2458 3904 2475 3968
rect 2539 3904 2556 3968
rect 2620 3904 2637 3968
rect 2701 3904 2718 3968
rect 2782 3904 2799 3968
rect 2863 3904 2880 3968
rect 2944 3904 2961 3968
rect 3025 3904 3042 3968
rect 3106 3904 3123 3968
rect 3187 3904 3204 3968
rect 3268 3904 3285 3968
rect 3349 3904 3366 3968
rect 3430 3904 3447 3968
rect 3511 3904 3528 3968
rect 3592 3904 3609 3968
rect 3673 3904 3690 3968
rect 3754 3904 3771 3968
rect 3835 3904 3852 3968
rect 3916 3904 3933 3968
rect 3997 3904 4014 3968
rect 4078 3904 4095 3968
rect 4159 3904 4176 3968
rect 4240 3904 4257 3968
rect 4321 3904 4338 3968
rect 4402 3904 4420 3968
rect 4484 3904 4502 3968
rect 4566 3904 4584 3968
rect 4648 3904 4666 3968
rect 4730 3904 4748 3968
rect 4812 3904 4830 3968
rect 4894 3904 4895 3968
rect 0 3882 4895 3904
rect 0 3818 126 3882
rect 190 3818 207 3882
rect 271 3818 288 3882
rect 352 3818 369 3882
rect 433 3818 450 3882
rect 514 3818 531 3882
rect 595 3818 612 3882
rect 676 3818 693 3882
rect 757 3818 774 3882
rect 838 3818 855 3882
rect 919 3818 936 3882
rect 1000 3818 1017 3882
rect 1081 3818 1098 3882
rect 1162 3818 1179 3882
rect 1243 3818 1260 3882
rect 1324 3818 1341 3882
rect 1405 3818 1422 3882
rect 1486 3818 1503 3882
rect 1567 3818 1584 3882
rect 1648 3818 1665 3882
rect 1729 3818 1746 3882
rect 1810 3818 1827 3882
rect 1891 3818 1908 3882
rect 1972 3818 1989 3882
rect 2053 3818 2070 3882
rect 2134 3818 2151 3882
rect 2215 3818 2232 3882
rect 2296 3818 2313 3882
rect 2377 3818 2394 3882
rect 2458 3818 2475 3882
rect 2539 3818 2556 3882
rect 2620 3818 2637 3882
rect 2701 3818 2718 3882
rect 2782 3818 2799 3882
rect 2863 3818 2880 3882
rect 2944 3818 2961 3882
rect 3025 3818 3042 3882
rect 3106 3818 3123 3882
rect 3187 3818 3204 3882
rect 3268 3818 3285 3882
rect 3349 3818 3366 3882
rect 3430 3818 3447 3882
rect 3511 3818 3528 3882
rect 3592 3818 3609 3882
rect 3673 3818 3690 3882
rect 3754 3818 3771 3882
rect 3835 3818 3852 3882
rect 3916 3818 3933 3882
rect 3997 3818 4014 3882
rect 4078 3818 4095 3882
rect 4159 3818 4176 3882
rect 4240 3818 4257 3882
rect 4321 3818 4338 3882
rect 4402 3818 4420 3882
rect 4484 3818 4502 3882
rect 4566 3818 4584 3882
rect 4648 3818 4666 3882
rect 4730 3818 4748 3882
rect 4812 3818 4830 3882
rect 4894 3818 4895 3882
rect 0 3796 4895 3818
rect 0 3732 126 3796
rect 190 3732 207 3796
rect 271 3732 288 3796
rect 352 3732 369 3796
rect 433 3732 450 3796
rect 514 3732 531 3796
rect 595 3732 612 3796
rect 676 3732 693 3796
rect 757 3732 774 3796
rect 838 3732 855 3796
rect 919 3732 936 3796
rect 1000 3732 1017 3796
rect 1081 3732 1098 3796
rect 1162 3732 1179 3796
rect 1243 3732 1260 3796
rect 1324 3732 1341 3796
rect 1405 3732 1422 3796
rect 1486 3732 1503 3796
rect 1567 3732 1584 3796
rect 1648 3732 1665 3796
rect 1729 3732 1746 3796
rect 1810 3732 1827 3796
rect 1891 3732 1908 3796
rect 1972 3732 1989 3796
rect 2053 3732 2070 3796
rect 2134 3732 2151 3796
rect 2215 3732 2232 3796
rect 2296 3732 2313 3796
rect 2377 3732 2394 3796
rect 2458 3732 2475 3796
rect 2539 3732 2556 3796
rect 2620 3732 2637 3796
rect 2701 3732 2718 3796
rect 2782 3732 2799 3796
rect 2863 3732 2880 3796
rect 2944 3732 2961 3796
rect 3025 3732 3042 3796
rect 3106 3732 3123 3796
rect 3187 3732 3204 3796
rect 3268 3732 3285 3796
rect 3349 3732 3366 3796
rect 3430 3732 3447 3796
rect 3511 3732 3528 3796
rect 3592 3732 3609 3796
rect 3673 3732 3690 3796
rect 3754 3732 3771 3796
rect 3835 3732 3852 3796
rect 3916 3732 3933 3796
rect 3997 3732 4014 3796
rect 4078 3732 4095 3796
rect 4159 3732 4176 3796
rect 4240 3732 4257 3796
rect 4321 3732 4338 3796
rect 4402 3732 4420 3796
rect 4484 3732 4502 3796
rect 4566 3732 4584 3796
rect 4648 3732 4666 3796
rect 4730 3732 4748 3796
rect 4812 3732 4830 3796
rect 4894 3732 4895 3796
rect 0 3710 4895 3732
rect 0 3646 126 3710
rect 190 3646 207 3710
rect 271 3646 288 3710
rect 352 3646 369 3710
rect 433 3646 450 3710
rect 514 3646 531 3710
rect 595 3646 612 3710
rect 676 3646 693 3710
rect 757 3646 774 3710
rect 838 3646 855 3710
rect 919 3646 936 3710
rect 1000 3646 1017 3710
rect 1081 3646 1098 3710
rect 1162 3646 1179 3710
rect 1243 3646 1260 3710
rect 1324 3646 1341 3710
rect 1405 3646 1422 3710
rect 1486 3646 1503 3710
rect 1567 3646 1584 3710
rect 1648 3646 1665 3710
rect 1729 3646 1746 3710
rect 1810 3646 1827 3710
rect 1891 3646 1908 3710
rect 1972 3646 1989 3710
rect 2053 3646 2070 3710
rect 2134 3646 2151 3710
rect 2215 3646 2232 3710
rect 2296 3646 2313 3710
rect 2377 3646 2394 3710
rect 2458 3646 2475 3710
rect 2539 3646 2556 3710
rect 2620 3646 2637 3710
rect 2701 3646 2718 3710
rect 2782 3646 2799 3710
rect 2863 3646 2880 3710
rect 2944 3646 2961 3710
rect 3025 3646 3042 3710
rect 3106 3646 3123 3710
rect 3187 3646 3204 3710
rect 3268 3646 3285 3710
rect 3349 3646 3366 3710
rect 3430 3646 3447 3710
rect 3511 3646 3528 3710
rect 3592 3646 3609 3710
rect 3673 3646 3690 3710
rect 3754 3646 3771 3710
rect 3835 3646 3852 3710
rect 3916 3646 3933 3710
rect 3997 3646 4014 3710
rect 4078 3646 4095 3710
rect 4159 3646 4176 3710
rect 4240 3646 4257 3710
rect 4321 3646 4338 3710
rect 4402 3646 4420 3710
rect 4484 3646 4502 3710
rect 4566 3646 4584 3710
rect 4648 3646 4666 3710
rect 4730 3646 4748 3710
rect 4812 3646 4830 3710
rect 4894 3646 4895 3710
rect 0 3624 4895 3646
rect 0 3560 126 3624
rect 190 3560 207 3624
rect 271 3560 288 3624
rect 352 3560 369 3624
rect 433 3560 450 3624
rect 514 3560 531 3624
rect 595 3560 612 3624
rect 676 3560 693 3624
rect 757 3560 774 3624
rect 838 3560 855 3624
rect 919 3560 936 3624
rect 1000 3560 1017 3624
rect 1081 3560 1098 3624
rect 1162 3560 1179 3624
rect 1243 3560 1260 3624
rect 1324 3560 1341 3624
rect 1405 3560 1422 3624
rect 1486 3560 1503 3624
rect 1567 3560 1584 3624
rect 1648 3560 1665 3624
rect 1729 3560 1746 3624
rect 1810 3560 1827 3624
rect 1891 3560 1908 3624
rect 1972 3560 1989 3624
rect 2053 3560 2070 3624
rect 2134 3560 2151 3624
rect 2215 3560 2232 3624
rect 2296 3560 2313 3624
rect 2377 3560 2394 3624
rect 2458 3560 2475 3624
rect 2539 3560 2556 3624
rect 2620 3560 2637 3624
rect 2701 3560 2718 3624
rect 2782 3560 2799 3624
rect 2863 3560 2880 3624
rect 2944 3560 2961 3624
rect 3025 3560 3042 3624
rect 3106 3560 3123 3624
rect 3187 3560 3204 3624
rect 3268 3560 3285 3624
rect 3349 3560 3366 3624
rect 3430 3560 3447 3624
rect 3511 3560 3528 3624
rect 3592 3560 3609 3624
rect 3673 3560 3690 3624
rect 3754 3560 3771 3624
rect 3835 3560 3852 3624
rect 3916 3560 3933 3624
rect 3997 3560 4014 3624
rect 4078 3560 4095 3624
rect 4159 3560 4176 3624
rect 4240 3560 4257 3624
rect 4321 3560 4338 3624
rect 4402 3560 4420 3624
rect 4484 3560 4502 3624
rect 4566 3560 4584 3624
rect 4648 3560 4666 3624
rect 4730 3560 4748 3624
rect 4812 3560 4830 3624
rect 4894 3560 4895 3624
rect 0 3557 4895 3560
rect 10156 4484 15000 4487
rect 10156 4420 10157 4484
rect 10221 4420 10238 4484
rect 10302 4420 10319 4484
rect 10383 4420 10400 4484
rect 10464 4420 10481 4484
rect 10545 4420 10562 4484
rect 10626 4420 10643 4484
rect 10707 4420 10724 4484
rect 10788 4420 10805 4484
rect 10869 4420 10886 4484
rect 10950 4420 10967 4484
rect 11031 4420 11048 4484
rect 11112 4420 11129 4484
rect 11193 4420 11210 4484
rect 11274 4420 11291 4484
rect 11355 4420 11372 4484
rect 11436 4420 11453 4484
rect 11517 4420 11534 4484
rect 11598 4420 11615 4484
rect 11679 4420 11696 4484
rect 11760 4420 11777 4484
rect 11841 4420 11858 4484
rect 11922 4420 11939 4484
rect 12003 4420 12020 4484
rect 12084 4420 12101 4484
rect 12165 4420 12182 4484
rect 12246 4420 12263 4484
rect 12327 4420 12344 4484
rect 12408 4420 12425 4484
rect 12489 4420 12506 4484
rect 12570 4420 12587 4484
rect 12651 4420 12668 4484
rect 12732 4420 12749 4484
rect 12813 4420 12830 4484
rect 12894 4420 12911 4484
rect 12975 4420 12992 4484
rect 13056 4420 13073 4484
rect 13137 4420 13154 4484
rect 13218 4420 13235 4484
rect 13299 4420 13316 4484
rect 13380 4420 13397 4484
rect 13461 4420 13478 4484
rect 13542 4420 13559 4484
rect 13623 4420 13640 4484
rect 13704 4420 13721 4484
rect 13785 4420 13802 4484
rect 13866 4420 13883 4484
rect 13947 4420 13964 4484
rect 14028 4420 14045 4484
rect 14109 4420 14126 4484
rect 14190 4420 14207 4484
rect 14271 4420 14288 4484
rect 14352 4420 14369 4484
rect 14433 4420 14451 4484
rect 14515 4420 14533 4484
rect 14597 4420 14615 4484
rect 14679 4420 14697 4484
rect 14761 4420 14779 4484
rect 14843 4420 14861 4484
rect 14925 4420 15000 4484
rect 10156 4398 15000 4420
rect 10156 4334 10157 4398
rect 10221 4334 10238 4398
rect 10302 4334 10319 4398
rect 10383 4334 10400 4398
rect 10464 4334 10481 4398
rect 10545 4334 10562 4398
rect 10626 4334 10643 4398
rect 10707 4334 10724 4398
rect 10788 4334 10805 4398
rect 10869 4334 10886 4398
rect 10950 4334 10967 4398
rect 11031 4334 11048 4398
rect 11112 4334 11129 4398
rect 11193 4334 11210 4398
rect 11274 4334 11291 4398
rect 11355 4334 11372 4398
rect 11436 4334 11453 4398
rect 11517 4334 11534 4398
rect 11598 4334 11615 4398
rect 11679 4334 11696 4398
rect 11760 4334 11777 4398
rect 11841 4334 11858 4398
rect 11922 4334 11939 4398
rect 12003 4334 12020 4398
rect 12084 4334 12101 4398
rect 12165 4334 12182 4398
rect 12246 4334 12263 4398
rect 12327 4334 12344 4398
rect 12408 4334 12425 4398
rect 12489 4334 12506 4398
rect 12570 4334 12587 4398
rect 12651 4334 12668 4398
rect 12732 4334 12749 4398
rect 12813 4334 12830 4398
rect 12894 4334 12911 4398
rect 12975 4334 12992 4398
rect 13056 4334 13073 4398
rect 13137 4334 13154 4398
rect 13218 4334 13235 4398
rect 13299 4334 13316 4398
rect 13380 4334 13397 4398
rect 13461 4334 13478 4398
rect 13542 4334 13559 4398
rect 13623 4334 13640 4398
rect 13704 4334 13721 4398
rect 13785 4334 13802 4398
rect 13866 4334 13883 4398
rect 13947 4334 13964 4398
rect 14028 4334 14045 4398
rect 14109 4334 14126 4398
rect 14190 4334 14207 4398
rect 14271 4334 14288 4398
rect 14352 4334 14369 4398
rect 14433 4334 14451 4398
rect 14515 4334 14533 4398
rect 14597 4334 14615 4398
rect 14679 4334 14697 4398
rect 14761 4334 14779 4398
rect 14843 4334 14861 4398
rect 14925 4334 15000 4398
rect 10156 4312 15000 4334
rect 10156 4248 10157 4312
rect 10221 4248 10238 4312
rect 10302 4248 10319 4312
rect 10383 4248 10400 4312
rect 10464 4248 10481 4312
rect 10545 4248 10562 4312
rect 10626 4248 10643 4312
rect 10707 4248 10724 4312
rect 10788 4248 10805 4312
rect 10869 4248 10886 4312
rect 10950 4248 10967 4312
rect 11031 4248 11048 4312
rect 11112 4248 11129 4312
rect 11193 4248 11210 4312
rect 11274 4248 11291 4312
rect 11355 4248 11372 4312
rect 11436 4248 11453 4312
rect 11517 4248 11534 4312
rect 11598 4248 11615 4312
rect 11679 4248 11696 4312
rect 11760 4248 11777 4312
rect 11841 4248 11858 4312
rect 11922 4248 11939 4312
rect 12003 4248 12020 4312
rect 12084 4248 12101 4312
rect 12165 4248 12182 4312
rect 12246 4248 12263 4312
rect 12327 4248 12344 4312
rect 12408 4248 12425 4312
rect 12489 4248 12506 4312
rect 12570 4248 12587 4312
rect 12651 4248 12668 4312
rect 12732 4248 12749 4312
rect 12813 4248 12830 4312
rect 12894 4248 12911 4312
rect 12975 4248 12992 4312
rect 13056 4248 13073 4312
rect 13137 4248 13154 4312
rect 13218 4248 13235 4312
rect 13299 4248 13316 4312
rect 13380 4248 13397 4312
rect 13461 4248 13478 4312
rect 13542 4248 13559 4312
rect 13623 4248 13640 4312
rect 13704 4248 13721 4312
rect 13785 4248 13802 4312
rect 13866 4248 13883 4312
rect 13947 4248 13964 4312
rect 14028 4248 14045 4312
rect 14109 4248 14126 4312
rect 14190 4248 14207 4312
rect 14271 4248 14288 4312
rect 14352 4248 14369 4312
rect 14433 4248 14451 4312
rect 14515 4248 14533 4312
rect 14597 4248 14615 4312
rect 14679 4248 14697 4312
rect 14761 4248 14779 4312
rect 14843 4248 14861 4312
rect 14925 4248 15000 4312
rect 10156 4226 15000 4248
rect 10156 4162 10157 4226
rect 10221 4162 10238 4226
rect 10302 4162 10319 4226
rect 10383 4162 10400 4226
rect 10464 4162 10481 4226
rect 10545 4162 10562 4226
rect 10626 4162 10643 4226
rect 10707 4162 10724 4226
rect 10788 4162 10805 4226
rect 10869 4162 10886 4226
rect 10950 4162 10967 4226
rect 11031 4162 11048 4226
rect 11112 4162 11129 4226
rect 11193 4162 11210 4226
rect 11274 4162 11291 4226
rect 11355 4162 11372 4226
rect 11436 4162 11453 4226
rect 11517 4162 11534 4226
rect 11598 4162 11615 4226
rect 11679 4162 11696 4226
rect 11760 4162 11777 4226
rect 11841 4162 11858 4226
rect 11922 4162 11939 4226
rect 12003 4162 12020 4226
rect 12084 4162 12101 4226
rect 12165 4162 12182 4226
rect 12246 4162 12263 4226
rect 12327 4162 12344 4226
rect 12408 4162 12425 4226
rect 12489 4162 12506 4226
rect 12570 4162 12587 4226
rect 12651 4162 12668 4226
rect 12732 4162 12749 4226
rect 12813 4162 12830 4226
rect 12894 4162 12911 4226
rect 12975 4162 12992 4226
rect 13056 4162 13073 4226
rect 13137 4162 13154 4226
rect 13218 4162 13235 4226
rect 13299 4162 13316 4226
rect 13380 4162 13397 4226
rect 13461 4162 13478 4226
rect 13542 4162 13559 4226
rect 13623 4162 13640 4226
rect 13704 4162 13721 4226
rect 13785 4162 13802 4226
rect 13866 4162 13883 4226
rect 13947 4162 13964 4226
rect 14028 4162 14045 4226
rect 14109 4162 14126 4226
rect 14190 4162 14207 4226
rect 14271 4162 14288 4226
rect 14352 4162 14369 4226
rect 14433 4162 14451 4226
rect 14515 4162 14533 4226
rect 14597 4162 14615 4226
rect 14679 4162 14697 4226
rect 14761 4162 14779 4226
rect 14843 4162 14861 4226
rect 14925 4162 15000 4226
rect 10156 4140 15000 4162
rect 10156 4076 10157 4140
rect 10221 4076 10238 4140
rect 10302 4076 10319 4140
rect 10383 4076 10400 4140
rect 10464 4076 10481 4140
rect 10545 4076 10562 4140
rect 10626 4076 10643 4140
rect 10707 4076 10724 4140
rect 10788 4076 10805 4140
rect 10869 4076 10886 4140
rect 10950 4076 10967 4140
rect 11031 4076 11048 4140
rect 11112 4076 11129 4140
rect 11193 4076 11210 4140
rect 11274 4076 11291 4140
rect 11355 4076 11372 4140
rect 11436 4076 11453 4140
rect 11517 4076 11534 4140
rect 11598 4076 11615 4140
rect 11679 4076 11696 4140
rect 11760 4076 11777 4140
rect 11841 4076 11858 4140
rect 11922 4076 11939 4140
rect 12003 4076 12020 4140
rect 12084 4076 12101 4140
rect 12165 4076 12182 4140
rect 12246 4076 12263 4140
rect 12327 4076 12344 4140
rect 12408 4076 12425 4140
rect 12489 4076 12506 4140
rect 12570 4076 12587 4140
rect 12651 4076 12668 4140
rect 12732 4076 12749 4140
rect 12813 4076 12830 4140
rect 12894 4076 12911 4140
rect 12975 4076 12992 4140
rect 13056 4076 13073 4140
rect 13137 4076 13154 4140
rect 13218 4076 13235 4140
rect 13299 4076 13316 4140
rect 13380 4076 13397 4140
rect 13461 4076 13478 4140
rect 13542 4076 13559 4140
rect 13623 4076 13640 4140
rect 13704 4076 13721 4140
rect 13785 4076 13802 4140
rect 13866 4076 13883 4140
rect 13947 4076 13964 4140
rect 14028 4076 14045 4140
rect 14109 4076 14126 4140
rect 14190 4076 14207 4140
rect 14271 4076 14288 4140
rect 14352 4076 14369 4140
rect 14433 4076 14451 4140
rect 14515 4076 14533 4140
rect 14597 4076 14615 4140
rect 14679 4076 14697 4140
rect 14761 4076 14779 4140
rect 14843 4076 14861 4140
rect 14925 4076 15000 4140
rect 10156 4054 15000 4076
rect 10156 3990 10157 4054
rect 10221 3990 10238 4054
rect 10302 3990 10319 4054
rect 10383 3990 10400 4054
rect 10464 3990 10481 4054
rect 10545 3990 10562 4054
rect 10626 3990 10643 4054
rect 10707 3990 10724 4054
rect 10788 3990 10805 4054
rect 10869 3990 10886 4054
rect 10950 3990 10967 4054
rect 11031 3990 11048 4054
rect 11112 3990 11129 4054
rect 11193 3990 11210 4054
rect 11274 3990 11291 4054
rect 11355 3990 11372 4054
rect 11436 3990 11453 4054
rect 11517 3990 11534 4054
rect 11598 3990 11615 4054
rect 11679 3990 11696 4054
rect 11760 3990 11777 4054
rect 11841 3990 11858 4054
rect 11922 3990 11939 4054
rect 12003 3990 12020 4054
rect 12084 3990 12101 4054
rect 12165 3990 12182 4054
rect 12246 3990 12263 4054
rect 12327 3990 12344 4054
rect 12408 3990 12425 4054
rect 12489 3990 12506 4054
rect 12570 3990 12587 4054
rect 12651 3990 12668 4054
rect 12732 3990 12749 4054
rect 12813 3990 12830 4054
rect 12894 3990 12911 4054
rect 12975 3990 12992 4054
rect 13056 3990 13073 4054
rect 13137 3990 13154 4054
rect 13218 3990 13235 4054
rect 13299 3990 13316 4054
rect 13380 3990 13397 4054
rect 13461 3990 13478 4054
rect 13542 3990 13559 4054
rect 13623 3990 13640 4054
rect 13704 3990 13721 4054
rect 13785 3990 13802 4054
rect 13866 3990 13883 4054
rect 13947 3990 13964 4054
rect 14028 3990 14045 4054
rect 14109 3990 14126 4054
rect 14190 3990 14207 4054
rect 14271 3990 14288 4054
rect 14352 3990 14369 4054
rect 14433 3990 14451 4054
rect 14515 3990 14533 4054
rect 14597 3990 14615 4054
rect 14679 3990 14697 4054
rect 14761 3990 14779 4054
rect 14843 3990 14861 4054
rect 14925 3990 15000 4054
rect 10156 3968 15000 3990
rect 10156 3904 10157 3968
rect 10221 3904 10238 3968
rect 10302 3904 10319 3968
rect 10383 3904 10400 3968
rect 10464 3904 10481 3968
rect 10545 3904 10562 3968
rect 10626 3904 10643 3968
rect 10707 3904 10724 3968
rect 10788 3904 10805 3968
rect 10869 3904 10886 3968
rect 10950 3904 10967 3968
rect 11031 3904 11048 3968
rect 11112 3904 11129 3968
rect 11193 3904 11210 3968
rect 11274 3904 11291 3968
rect 11355 3904 11372 3968
rect 11436 3904 11453 3968
rect 11517 3904 11534 3968
rect 11598 3904 11615 3968
rect 11679 3904 11696 3968
rect 11760 3904 11777 3968
rect 11841 3904 11858 3968
rect 11922 3904 11939 3968
rect 12003 3904 12020 3968
rect 12084 3904 12101 3968
rect 12165 3904 12182 3968
rect 12246 3904 12263 3968
rect 12327 3904 12344 3968
rect 12408 3904 12425 3968
rect 12489 3904 12506 3968
rect 12570 3904 12587 3968
rect 12651 3904 12668 3968
rect 12732 3904 12749 3968
rect 12813 3904 12830 3968
rect 12894 3904 12911 3968
rect 12975 3904 12992 3968
rect 13056 3904 13073 3968
rect 13137 3904 13154 3968
rect 13218 3904 13235 3968
rect 13299 3904 13316 3968
rect 13380 3904 13397 3968
rect 13461 3904 13478 3968
rect 13542 3904 13559 3968
rect 13623 3904 13640 3968
rect 13704 3904 13721 3968
rect 13785 3904 13802 3968
rect 13866 3904 13883 3968
rect 13947 3904 13964 3968
rect 14028 3904 14045 3968
rect 14109 3904 14126 3968
rect 14190 3904 14207 3968
rect 14271 3904 14288 3968
rect 14352 3904 14369 3968
rect 14433 3904 14451 3968
rect 14515 3904 14533 3968
rect 14597 3904 14615 3968
rect 14679 3904 14697 3968
rect 14761 3904 14779 3968
rect 14843 3904 14861 3968
rect 14925 3904 15000 3968
rect 10156 3882 15000 3904
rect 10156 3818 10157 3882
rect 10221 3818 10238 3882
rect 10302 3818 10319 3882
rect 10383 3818 10400 3882
rect 10464 3818 10481 3882
rect 10545 3818 10562 3882
rect 10626 3818 10643 3882
rect 10707 3818 10724 3882
rect 10788 3818 10805 3882
rect 10869 3818 10886 3882
rect 10950 3818 10967 3882
rect 11031 3818 11048 3882
rect 11112 3818 11129 3882
rect 11193 3818 11210 3882
rect 11274 3818 11291 3882
rect 11355 3818 11372 3882
rect 11436 3818 11453 3882
rect 11517 3818 11534 3882
rect 11598 3818 11615 3882
rect 11679 3818 11696 3882
rect 11760 3818 11777 3882
rect 11841 3818 11858 3882
rect 11922 3818 11939 3882
rect 12003 3818 12020 3882
rect 12084 3818 12101 3882
rect 12165 3818 12182 3882
rect 12246 3818 12263 3882
rect 12327 3818 12344 3882
rect 12408 3818 12425 3882
rect 12489 3818 12506 3882
rect 12570 3818 12587 3882
rect 12651 3818 12668 3882
rect 12732 3818 12749 3882
rect 12813 3818 12830 3882
rect 12894 3818 12911 3882
rect 12975 3818 12992 3882
rect 13056 3818 13073 3882
rect 13137 3818 13154 3882
rect 13218 3818 13235 3882
rect 13299 3818 13316 3882
rect 13380 3818 13397 3882
rect 13461 3818 13478 3882
rect 13542 3818 13559 3882
rect 13623 3818 13640 3882
rect 13704 3818 13721 3882
rect 13785 3818 13802 3882
rect 13866 3818 13883 3882
rect 13947 3818 13964 3882
rect 14028 3818 14045 3882
rect 14109 3818 14126 3882
rect 14190 3818 14207 3882
rect 14271 3818 14288 3882
rect 14352 3818 14369 3882
rect 14433 3818 14451 3882
rect 14515 3818 14533 3882
rect 14597 3818 14615 3882
rect 14679 3818 14697 3882
rect 14761 3818 14779 3882
rect 14843 3818 14861 3882
rect 14925 3818 15000 3882
rect 10156 3796 15000 3818
rect 10156 3732 10157 3796
rect 10221 3732 10238 3796
rect 10302 3732 10319 3796
rect 10383 3732 10400 3796
rect 10464 3732 10481 3796
rect 10545 3732 10562 3796
rect 10626 3732 10643 3796
rect 10707 3732 10724 3796
rect 10788 3732 10805 3796
rect 10869 3732 10886 3796
rect 10950 3732 10967 3796
rect 11031 3732 11048 3796
rect 11112 3732 11129 3796
rect 11193 3732 11210 3796
rect 11274 3732 11291 3796
rect 11355 3732 11372 3796
rect 11436 3732 11453 3796
rect 11517 3732 11534 3796
rect 11598 3732 11615 3796
rect 11679 3732 11696 3796
rect 11760 3732 11777 3796
rect 11841 3732 11858 3796
rect 11922 3732 11939 3796
rect 12003 3732 12020 3796
rect 12084 3732 12101 3796
rect 12165 3732 12182 3796
rect 12246 3732 12263 3796
rect 12327 3732 12344 3796
rect 12408 3732 12425 3796
rect 12489 3732 12506 3796
rect 12570 3732 12587 3796
rect 12651 3732 12668 3796
rect 12732 3732 12749 3796
rect 12813 3732 12830 3796
rect 12894 3732 12911 3796
rect 12975 3732 12992 3796
rect 13056 3732 13073 3796
rect 13137 3732 13154 3796
rect 13218 3732 13235 3796
rect 13299 3732 13316 3796
rect 13380 3732 13397 3796
rect 13461 3732 13478 3796
rect 13542 3732 13559 3796
rect 13623 3732 13640 3796
rect 13704 3732 13721 3796
rect 13785 3732 13802 3796
rect 13866 3732 13883 3796
rect 13947 3732 13964 3796
rect 14028 3732 14045 3796
rect 14109 3732 14126 3796
rect 14190 3732 14207 3796
rect 14271 3732 14288 3796
rect 14352 3732 14369 3796
rect 14433 3732 14451 3796
rect 14515 3732 14533 3796
rect 14597 3732 14615 3796
rect 14679 3732 14697 3796
rect 14761 3732 14779 3796
rect 14843 3732 14861 3796
rect 14925 3732 15000 3796
rect 10156 3710 15000 3732
rect 10156 3646 10157 3710
rect 10221 3646 10238 3710
rect 10302 3646 10319 3710
rect 10383 3646 10400 3710
rect 10464 3646 10481 3710
rect 10545 3646 10562 3710
rect 10626 3646 10643 3710
rect 10707 3646 10724 3710
rect 10788 3646 10805 3710
rect 10869 3646 10886 3710
rect 10950 3646 10967 3710
rect 11031 3646 11048 3710
rect 11112 3646 11129 3710
rect 11193 3646 11210 3710
rect 11274 3646 11291 3710
rect 11355 3646 11372 3710
rect 11436 3646 11453 3710
rect 11517 3646 11534 3710
rect 11598 3646 11615 3710
rect 11679 3646 11696 3710
rect 11760 3646 11777 3710
rect 11841 3646 11858 3710
rect 11922 3646 11939 3710
rect 12003 3646 12020 3710
rect 12084 3646 12101 3710
rect 12165 3646 12182 3710
rect 12246 3646 12263 3710
rect 12327 3646 12344 3710
rect 12408 3646 12425 3710
rect 12489 3646 12506 3710
rect 12570 3646 12587 3710
rect 12651 3646 12668 3710
rect 12732 3646 12749 3710
rect 12813 3646 12830 3710
rect 12894 3646 12911 3710
rect 12975 3646 12992 3710
rect 13056 3646 13073 3710
rect 13137 3646 13154 3710
rect 13218 3646 13235 3710
rect 13299 3646 13316 3710
rect 13380 3646 13397 3710
rect 13461 3646 13478 3710
rect 13542 3646 13559 3710
rect 13623 3646 13640 3710
rect 13704 3646 13721 3710
rect 13785 3646 13802 3710
rect 13866 3646 13883 3710
rect 13947 3646 13964 3710
rect 14028 3646 14045 3710
rect 14109 3646 14126 3710
rect 14190 3646 14207 3710
rect 14271 3646 14288 3710
rect 14352 3646 14369 3710
rect 14433 3646 14451 3710
rect 14515 3646 14533 3710
rect 14597 3646 14615 3710
rect 14679 3646 14697 3710
rect 14761 3646 14779 3710
rect 14843 3646 14861 3710
rect 14925 3646 15000 3710
rect 10156 3624 15000 3646
rect 10156 3560 10157 3624
rect 10221 3560 10238 3624
rect 10302 3560 10319 3624
rect 10383 3560 10400 3624
rect 10464 3560 10481 3624
rect 10545 3560 10562 3624
rect 10626 3560 10643 3624
rect 10707 3560 10724 3624
rect 10788 3560 10805 3624
rect 10869 3560 10886 3624
rect 10950 3560 10967 3624
rect 11031 3560 11048 3624
rect 11112 3560 11129 3624
rect 11193 3560 11210 3624
rect 11274 3560 11291 3624
rect 11355 3560 11372 3624
rect 11436 3560 11453 3624
rect 11517 3560 11534 3624
rect 11598 3560 11615 3624
rect 11679 3560 11696 3624
rect 11760 3560 11777 3624
rect 11841 3560 11858 3624
rect 11922 3560 11939 3624
rect 12003 3560 12020 3624
rect 12084 3560 12101 3624
rect 12165 3560 12182 3624
rect 12246 3560 12263 3624
rect 12327 3560 12344 3624
rect 12408 3560 12425 3624
rect 12489 3560 12506 3624
rect 12570 3560 12587 3624
rect 12651 3560 12668 3624
rect 12732 3560 12749 3624
rect 12813 3560 12830 3624
rect 12894 3560 12911 3624
rect 12975 3560 12992 3624
rect 13056 3560 13073 3624
rect 13137 3560 13154 3624
rect 13218 3560 13235 3624
rect 13299 3560 13316 3624
rect 13380 3560 13397 3624
rect 13461 3560 13478 3624
rect 13542 3560 13559 3624
rect 13623 3560 13640 3624
rect 13704 3560 13721 3624
rect 13785 3560 13802 3624
rect 13866 3560 13883 3624
rect 13947 3560 13964 3624
rect 14028 3560 14045 3624
rect 14109 3560 14126 3624
rect 14190 3560 14207 3624
rect 14271 3560 14288 3624
rect 14352 3560 14369 3624
rect 14433 3560 14451 3624
rect 14515 3560 14533 3624
rect 14597 3560 14615 3624
rect 14679 3560 14697 3624
rect 14761 3560 14779 3624
rect 14843 3560 14861 3624
rect 14925 3560 15000 3624
rect 10156 3557 15000 3560
rect 0 2587 193 3277
rect 14807 2587 15000 3277
rect 0 1377 254 2307
rect 14746 1377 15000 2307
rect 0 7 254 1097
rect 14746 7 15000 1097
<< metal5 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18597
rect 14746 13607 15000 18597
rect 0 12437 254 13287
rect 14746 12437 15000 13287
rect 0 11267 254 12117
rect 14746 11267 15000 12117
rect 0 9147 254 10947
rect 14746 9147 15000 10947
rect 0 7937 254 8827
rect 14746 7937 15000 8827
rect 0 6968 254 7617
rect 14746 6968 15000 7617
rect 0 5997 254 6647
rect 14746 5997 15000 6647
rect 0 4787 254 5677
rect 14746 4787 15000 5677
rect 0 3577 254 4467
rect 14746 3577 15000 4467
rect 0 2607 193 3257
rect 14807 2607 15000 3257
rect 0 1397 254 2287
rect 14746 1397 15000 2287
rect 0 27 254 1077
rect 14746 27 15000 1077
use sky130_fd_io__com_bus_hookup  sky130_fd_io__com_bus_hookup_0
timestamp 1619862920
transform 1 0 0 0 1 149
box 0 -142 15000 39451
<< labels >>
flabel metal5 s 14746 12437 15000 13287 3 FreeSans 520 180 0 0 VDDIO_Q
port 1 nsew power bidirectional
flabel metal5 s 14807 2607 15000 3257 3 FreeSans 520 180 0 0 VDDA
port 2 nsew power bidirectional
flabel metal5 s 0 12437 254 13287 3 FreeSans 520 0 0 0 VDDIO_Q
port 1 nsew power bidirectional
flabel metal5 s 14746 9147 15000 10947 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal5 s 14746 6968 15000 7617 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal5 s 0 1397 254 2287 3 FreeSans 520 0 0 0 VCCD
port 4 nsew power bidirectional
flabel metal5 s 0 9147 254 10947 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal5 s 0 6968 254 7617 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal5 s 0 27 254 1077 3 FreeSans 520 0 0 0 VCCHIB
port 5 nsew power bidirectional
flabel metal5 s 14746 7937 15000 8827 3 FreeSans 520 180 0 0 VSSD
port 6 nsew ground bidirectional
flabel metal5 s 0 2607 193 3257 3 FreeSans 520 0 0 0 VDDA
port 2 nsew power bidirectional
flabel metal5 s 14746 13607 15000 18597 3 FreeSans 520 180 0 0 VDDIO
port 7 nsew power bidirectional
flabel metal5 s 14746 3577 15000 4467 3 FreeSans 520 180 0 0 VDDIO
port 7 nsew power bidirectional
flabel metal5 s 0 13607 254 18597 3 FreeSans 520 0 0 0 VDDIO
port 7 nsew power bidirectional
flabel metal5 s 0 3577 254 4467 3 FreeSans 520 0 0 0 VDDIO
port 7 nsew power bidirectional
flabel metal5 s 14746 1397 15000 2287 3 FreeSans 520 180 0 0 VCCD
port 4 nsew power bidirectional
flabel metal5 s 14746 27 15000 1077 3 FreeSans 520 180 0 0 VCCHIB
port 5 nsew power bidirectional
flabel metal5 s 0 5997 254 6647 3 FreeSans 520 0 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal5 s 14746 5997 15000 6647 3 FreeSans 520 180 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal5 s 0 11267 254 12117 3 FreeSans 520 0 0 0 VSSIO_Q
port 9 nsew ground bidirectional
flabel metal5 s 14746 11267 15000 12117 3 FreeSans 520 180 0 0 VSSIO_Q
port 9 nsew ground bidirectional
flabel metal5 s 0 4787 254 5677 3 FreeSans 520 0 0 0 VSSIO
port 10 nsew ground bidirectional
flabel metal5 s 0 34757 254 39600 3 FreeSans 520 0 0 0 VSSIO
port 10 nsew ground bidirectional
flabel metal5 s 14746 4787 15000 5677 3 FreeSans 520 180 0 0 VSSIO
port 10 nsew ground bidirectional
flabel metal5 s 14746 34757 15000 39600 3 FreeSans 520 180 0 0 VSSIO
port 10 nsew ground bidirectional
flabel metal5 s 0 7937 254 8827 3 FreeSans 520 0 0 0 VSSD
port 6 nsew ground bidirectional
flabel metal4 s 0 12417 254 13307 3 FreeSans 520 0 0 0 VDDIO_Q
port 1 nsew power bidirectional
flabel metal4 s 14746 6947 15000 7637 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 14746 9147 15000 9213 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 14746 10881 15000 10947 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 14746 9929 15000 10165 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 0 9147 254 9213 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 0 9929 254 10165 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 0 10881 254 10947 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 0 6947 254 7637 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 14746 7917 15000 8847 3 FreeSans 520 180 0 0 VSSD
port 6 nsew ground bidirectional
flabel metal4 s 0 2587 193 3277 3 FreeSans 520 0 0 0 VDDA
port 2 nsew power bidirectional
flabel metal4 s 14746 3557 15000 4487 3 FreeSans 520 180 0 0 VDDIO
port 7 nsew power bidirectional
flabel metal4 s 14746 13607 15000 18600 3 FreeSans 520 180 0 0 VDDIO
port 7 nsew power bidirectional
flabel metal4 s 0 3557 254 4487 3 FreeSans 520 0 0 0 VDDIO
port 7 nsew power bidirectional
flabel metal4 s 0 13607 254 18600 3 FreeSans 520 0 0 0 VDDIO
port 7 nsew power bidirectional
flabel metal4 s 14746 12417 15000 13307 3 FreeSans 520 180 0 0 VDDIO_Q
port 1 nsew power bidirectional
flabel metal4 s 14746 10225 15000 10821 3 FreeSans 520 180 0 0 AMUXBUS_A
port 11 nsew signal bidirectional
flabel metal4 s 0 10225 254 10821 3 FreeSans 520 0 0 0 AMUXBUS_A
port 11 nsew signal bidirectional
flabel metal4 s 14746 9273 15000 9869 3 FreeSans 520 180 0 0 AMUXBUS_B
port 12 nsew signal bidirectional
flabel metal4 s 0 9273 254 9869 3 FreeSans 520 0 0 0 AMUXBUS_B
port 12 nsew signal bidirectional
flabel metal4 s 14746 1377 15000 2307 3 FreeSans 520 180 0 0 VCCD
port 4 nsew power bidirectional
flabel metal4 s 0 1377 254 2307 3 FreeSans 520 0 0 0 VCCD
port 4 nsew power bidirectional
flabel metal4 s 14746 7 15000 1097 3 FreeSans 520 180 0 0 VCCHIB
port 5 nsew power bidirectional
flabel metal4 s 0 7 254 1097 3 FreeSans 520 0 0 0 VCCHIB
port 5 nsew power bidirectional
flabel metal4 s 14807 2587 15000 3277 3 FreeSans 520 180 0 0 VDDA
port 2 nsew power bidirectional
flabel metal4 s 0 5977 254 6667 3 FreeSans 520 0 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal4 s 14746 5977 15000 6667 3 FreeSans 520 180 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal4 s 0 11247 254 12137 3 FreeSans 520 0 0 0 VSSIO_Q
port 9 nsew ground bidirectional
flabel metal4 s 14746 11247 15000 12137 3 FreeSans 520 180 0 0 VSSIO_Q
port 9 nsew ground bidirectional
flabel metal4 s 0 4767 254 5697 3 FreeSans 520 0 0 0 VSSIO
port 10 nsew ground bidirectional
flabel metal4 s 0 34757 254 39600 3 FreeSans 520 0 0 0 VSSIO
port 10 nsew ground bidirectional
flabel metal4 s 14746 4767 15000 5697 3 FreeSans 520 180 0 0 VSSIO
port 10 nsew ground bidirectional
flabel metal4 s 14746 34757 15000 39600 3 FreeSans 520 180 0 0 VSSIO
port 10 nsew ground bidirectional
flabel metal4 s 0 7917 254 8847 3 FreeSans 520 0 0 0 VSSD
port 6 nsew ground bidirectional
rlabel metal4 s 126 3646 190 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 126 3646 190 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 126 3732 190 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 126 3732 190 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 126 3818 190 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 126 3818 190 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 126 3904 190 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 126 3904 190 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 126 3990 190 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 126 3990 190 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 126 4076 190 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 126 4076 190 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 126 4162 190 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 126 4162 190 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 126 4248 190 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 126 4248 190 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 126 4334 190 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 126 4334 190 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 126 4420 190 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 126 4420 190 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 16559 199 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16559 199 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 16641 199 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16641 199 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 16723 199 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16723 199 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 16805 199 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16805 199 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 16887 199 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16887 199 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 16969 199 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16969 199 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 17051 199 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17051 199 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 17133 199 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17133 199 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 17215 199 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17215 199 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 17297 199 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17297 199 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 17379 199 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17379 199 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 17461 199 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17461 199 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 17543 199 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17543 199 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 17625 199 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17625 199 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 17707 199 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17707 199 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 17789 199 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17789 199 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 17871 199 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17871 199 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 17953 199 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17953 199 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 18035 199 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18035 199 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 18117 199 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18117 199 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 18199 199 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18199 199 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 18281 199 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18281 199 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 18363 199 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18363 199 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 18445 199 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18445 199 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 135 18527 199 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18527 199 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 13613 221 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 13613 221 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 13695 221 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 13695 221 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 13777 221 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 13777 221 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 13859 221 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 13859 221 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 13941 221 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 13941 221 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 14023 221 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14023 221 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 14105 221 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14105 221 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 14187 221 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14187 221 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 14269 221 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14269 221 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 14351 221 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14351 221 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 14433 221 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14433 221 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 14515 221 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14515 221 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 14597 221 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14597 221 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 14678 221 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14678 221 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 14759 221 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14759 221 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 14840 221 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14840 221 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 14921 221 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14921 221 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 15002 221 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15002 221 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 15083 221 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15083 221 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 15164 221 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15164 221 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 15245 221 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15245 221 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 15326 221 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15326 221 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 15407 221 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15407 221 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 15488 221 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15488 221 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 15569 221 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15569 221 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 15650 221 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15650 221 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 15731 221 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15731 221 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 15812 221 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15812 221 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 15893 221 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15893 221 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 15974 221 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15974 221 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 16055 221 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16055 221 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 16136 221 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16136 221 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 16217 221 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16217 221 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 16298 221 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16298 221 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 16379 221 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16379 221 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 157 16460 221 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16460 221 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 207 3560 271 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 207 3560 271 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 207 3646 271 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 207 3646 271 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 207 3732 271 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 207 3732 271 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 207 3818 271 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 207 3818 271 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 207 3904 271 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 207 3904 271 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 207 3990 271 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 207 3990 271 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 207 4076 271 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 207 4076 271 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 207 4162 271 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 207 4162 271 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 207 4248 271 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 207 4248 271 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 207 4334 271 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 207 4334 271 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 207 4420 271 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 207 4420 271 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 16559 281 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16559 281 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 16641 281 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16641 281 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 16723 281 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16723 281 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 16805 281 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16805 281 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 16887 281 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16887 281 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 16969 281 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16969 281 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 17051 281 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17051 281 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 17133 281 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17133 281 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 17215 281 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17215 281 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 17297 281 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17297 281 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 17379 281 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17379 281 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 17461 281 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17461 281 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 17543 281 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17543 281 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 17625 281 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17625 281 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 17707 281 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17707 281 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 17789 281 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17789 281 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 17871 281 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17871 281 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 17953 281 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17953 281 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 18035 281 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18035 281 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 18117 281 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18117 281 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 18199 281 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18199 281 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 18281 281 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18281 281 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 18363 281 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18363 281 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 18445 281 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18445 281 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 217 18527 281 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18527 281 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 13613 301 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 13613 301 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 13695 301 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 13695 301 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 13777 301 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 13777 301 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 13859 301 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 13859 301 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 13941 301 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 13941 301 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 14023 301 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14023 301 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 14105 301 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14105 301 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 14187 301 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14187 301 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 14269 301 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14269 301 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 14351 301 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14351 301 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 14433 301 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14433 301 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 14515 301 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14515 301 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 14597 301 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14597 301 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 14678 301 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14678 301 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 14759 301 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14759 301 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 14840 301 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14840 301 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 14921 301 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14921 301 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 15002 301 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15002 301 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 15083 301 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15083 301 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 15164 301 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15164 301 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 15245 301 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15245 301 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 15326 301 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15326 301 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 15407 301 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15407 301 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 15488 301 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15488 301 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 15569 301 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15569 301 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 15650 301 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15650 301 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 15731 301 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15731 301 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 15812 301 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15812 301 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 15893 301 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15893 301 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 15974 301 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15974 301 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 16055 301 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16055 301 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 16136 301 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16136 301 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 16217 301 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16217 301 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 16298 301 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16298 301 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 16379 301 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16379 301 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 237 16460 301 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16460 301 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 288 3560 352 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 288 3560 352 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 288 3646 352 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 288 3646 352 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 288 3732 352 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 288 3732 352 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 288 3818 352 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 288 3818 352 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 288 3904 352 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 288 3904 352 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 288 3990 352 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 288 3990 352 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 288 4076 352 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 288 4076 352 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 288 4162 352 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 288 4162 352 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 288 4248 352 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 288 4248 352 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 288 4334 352 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 288 4334 352 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 288 4420 352 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 288 4420 352 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 16559 363 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16559 363 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 16641 363 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16641 363 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 16723 363 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16723 363 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 16805 363 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16805 363 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 16887 363 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16887 363 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 16969 363 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16969 363 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17051 363 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17051 363 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17133 363 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17133 363 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17215 363 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17215 363 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17297 363 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17297 363 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17379 363 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17379 363 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17461 363 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17461 363 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17543 363 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17543 363 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17625 363 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17625 363 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17707 363 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17707 363 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17789 363 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17789 363 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17871 363 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17871 363 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17953 363 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17953 363 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 18035 363 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18035 363 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 18117 363 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18117 363 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 18199 363 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18199 363 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 18281 363 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18281 363 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 18363 363 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18363 363 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 18445 363 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18445 363 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 18527 363 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18527 363 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 13613 381 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 13613 381 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 13695 381 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 13695 381 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 13777 381 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 13777 381 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 13859 381 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 13859 381 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 13941 381 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 13941 381 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14023 381 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14023 381 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14105 381 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14105 381 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14187 381 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14187 381 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14269 381 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14269 381 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14351 381 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14351 381 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14433 381 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14433 381 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14515 381 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14515 381 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14597 381 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14597 381 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14678 381 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14678 381 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14759 381 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14759 381 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14840 381 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14840 381 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14921 381 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14921 381 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15002 381 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15002 381 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15083 381 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15083 381 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15164 381 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15164 381 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15245 381 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15245 381 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15326 381 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15326 381 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15407 381 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15407 381 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15488 381 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15488 381 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15569 381 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15569 381 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15650 381 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15650 381 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15731 381 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15731 381 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15812 381 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15812 381 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15893 381 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15893 381 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15974 381 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15974 381 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 16055 381 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16055 381 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 16136 381 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16136 381 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 16217 381 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16217 381 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 16298 381 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16298 381 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 16379 381 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16379 381 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 16460 381 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16460 381 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 369 3560 433 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 369 3560 433 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 369 3646 433 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 369 3646 433 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 369 3732 433 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 369 3732 433 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 369 3818 433 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 369 3818 433 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 369 3904 433 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 369 3904 433 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 369 3990 433 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 369 3990 433 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 369 4076 433 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 369 4076 433 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 369 4162 433 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 369 4162 433 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 369 4248 433 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 369 4248 433 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 369 4334 433 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 369 4334 433 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 369 4420 433 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 369 4420 433 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 16559 445 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16559 445 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 16641 445 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16641 445 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 16723 445 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16723 445 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 16805 445 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16805 445 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 16887 445 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16887 445 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 16969 445 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16969 445 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17051 445 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17051 445 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17133 445 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17133 445 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17215 445 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17215 445 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17297 445 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17297 445 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17379 445 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17379 445 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17461 445 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17461 445 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17543 445 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17543 445 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17625 445 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17625 445 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17707 445 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17707 445 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17789 445 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17789 445 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17871 445 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17871 445 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17953 445 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17953 445 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 18035 445 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18035 445 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 18117 445 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18117 445 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 18199 445 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18199 445 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 18281 445 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18281 445 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 18363 445 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18363 445 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 18445 445 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18445 445 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 18527 445 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18527 445 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 13613 461 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 13613 461 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 13695 461 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 13695 461 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 13777 461 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 13777 461 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 13859 461 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 13859 461 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 13941 461 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 13941 461 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14023 461 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14023 461 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14105 461 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14105 461 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14187 461 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14187 461 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14269 461 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14269 461 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14351 461 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14351 461 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14433 461 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14433 461 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14515 461 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14515 461 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14597 461 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14597 461 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14678 461 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14678 461 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14759 461 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14759 461 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14840 461 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14840 461 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14921 461 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14921 461 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15002 461 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15002 461 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15083 461 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15083 461 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15164 461 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15164 461 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15245 461 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15245 461 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15326 461 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15326 461 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15407 461 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15407 461 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15488 461 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15488 461 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15569 461 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15569 461 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15650 461 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15650 461 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15731 461 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15731 461 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15812 461 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15812 461 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15893 461 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15893 461 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15974 461 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15974 461 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 16055 461 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16055 461 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 16136 461 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16136 461 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 16217 461 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16217 461 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 16298 461 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16298 461 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 16379 461 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16379 461 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 16460 461 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16460 461 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 16559 2085 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16559 2085 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 16641 2085 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16641 2085 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 16723 2085 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16723 2085 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 16805 2085 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16805 2085 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 16887 2085 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16887 2085 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 16969 2085 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16969 2085 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17051 2085 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17051 2085 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17133 2085 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17133 2085 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17215 2085 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17215 2085 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17297 2085 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17297 2085 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17379 2085 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17379 2085 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17461 2085 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17461 2085 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17543 2085 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17543 2085 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17625 2085 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17625 2085 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17707 2085 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17707 2085 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17789 2085 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17789 2085 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17871 2085 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17871 2085 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17953 2085 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17953 2085 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 18035 2085 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18035 2085 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 18117 2085 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18117 2085 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 18199 2085 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18199 2085 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 18281 2085 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18281 2085 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 18363 2085 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18363 2085 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 18445 2085 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18445 2085 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 18527 2085 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18527 2085 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2070 3560 2134 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2070 3560 2134 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2070 3646 2134 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2070 3646 2134 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2070 3732 2134 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2070 3732 2134 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2070 3818 2134 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2070 3818 2134 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2070 3904 2134 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2070 3904 2134 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2070 3990 2134 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2070 3990 2134 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2070 4076 2134 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2070 4076 2134 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2070 4162 2134 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2070 4162 2134 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2070 4248 2134 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2070 4248 2134 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2070 4334 2134 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2070 4334 2134 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2070 4420 2134 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2070 4420 2134 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 13613 2141 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 13613 2141 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 13695 2141 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 13695 2141 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 13777 2141 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 13777 2141 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 13859 2141 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 13859 2141 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 13941 2141 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 13941 2141 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14023 2141 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14023 2141 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14105 2141 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14105 2141 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14187 2141 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14187 2141 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14269 2141 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14269 2141 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14351 2141 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14351 2141 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14433 2141 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14433 2141 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14515 2141 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14515 2141 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14597 2141 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14597 2141 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14678 2141 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14678 2141 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14759 2141 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14759 2141 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14840 2141 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14840 2141 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14921 2141 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14921 2141 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15002 2141 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15002 2141 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15083 2141 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15083 2141 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15164 2141 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15164 2141 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15245 2141 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15245 2141 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15326 2141 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15326 2141 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15407 2141 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15407 2141 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15488 2141 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15488 2141 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15569 2141 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15569 2141 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15650 2141 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15650 2141 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15731 2141 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15731 2141 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15812 2141 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15812 2141 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15893 2141 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15893 2141 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15974 2141 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15974 2141 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 16055 2141 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16055 2141 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 16136 2141 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16136 2141 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 16217 2141 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16217 2141 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 16298 2141 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16298 2141 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 16379 2141 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16379 2141 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 16460 2141 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16460 2141 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 16559 2167 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16559 2167 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 16641 2167 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16641 2167 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 16723 2167 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16723 2167 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 16805 2167 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16805 2167 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 16887 2167 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16887 2167 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 16969 2167 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16969 2167 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17051 2167 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17051 2167 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17133 2167 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17133 2167 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17215 2167 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17215 2167 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17297 2167 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17297 2167 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17379 2167 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17379 2167 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17461 2167 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17461 2167 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17543 2167 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17543 2167 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17625 2167 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17625 2167 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17707 2167 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17707 2167 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17789 2167 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17789 2167 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17871 2167 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17871 2167 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17953 2167 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17953 2167 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 18035 2167 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18035 2167 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 18117 2167 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18117 2167 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 18199 2167 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18199 2167 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 18281 2167 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18281 2167 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 18363 2167 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18363 2167 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 18445 2167 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18445 2167 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 18527 2167 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18527 2167 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2151 3560 2215 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2151 3560 2215 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2151 3646 2215 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2151 3646 2215 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2151 3732 2215 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2151 3732 2215 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2151 3818 2215 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2151 3818 2215 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2151 3904 2215 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2151 3904 2215 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2151 3990 2215 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2151 3990 2215 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2151 4076 2215 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2151 4076 2215 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2151 4162 2215 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2151 4162 2215 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2151 4248 2215 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2151 4248 2215 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2151 4334 2215 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2151 4334 2215 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2151 4420 2215 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2151 4420 2215 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 13613 2221 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 13613 2221 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 13695 2221 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 13695 2221 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 13777 2221 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 13777 2221 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 13859 2221 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 13859 2221 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 13941 2221 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 13941 2221 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14023 2221 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14023 2221 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14105 2221 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14105 2221 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14187 2221 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14187 2221 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14269 2221 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14269 2221 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14351 2221 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14351 2221 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14433 2221 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14433 2221 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14515 2221 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14515 2221 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14597 2221 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14597 2221 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14678 2221 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14678 2221 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14759 2221 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14759 2221 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14840 2221 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14840 2221 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14921 2221 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14921 2221 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15002 2221 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15002 2221 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15083 2221 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15083 2221 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15164 2221 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15164 2221 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15245 2221 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15245 2221 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15326 2221 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15326 2221 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15407 2221 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15407 2221 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15488 2221 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15488 2221 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15569 2221 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15569 2221 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15650 2221 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15650 2221 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15731 2221 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15731 2221 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15812 2221 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15812 2221 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15893 2221 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15893 2221 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15974 2221 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15974 2221 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 16055 2221 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16055 2221 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 16136 2221 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16136 2221 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 16217 2221 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16217 2221 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 16298 2221 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16298 2221 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 16379 2221 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16379 2221 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 16460 2221 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16460 2221 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 16559 2249 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16559 2249 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 16641 2249 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16641 2249 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 16723 2249 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16723 2249 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 16805 2249 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16805 2249 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 16887 2249 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16887 2249 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 16969 2249 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16969 2249 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17051 2249 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17051 2249 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17133 2249 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17133 2249 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17215 2249 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17215 2249 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17297 2249 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17297 2249 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17379 2249 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17379 2249 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17461 2249 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17461 2249 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17543 2249 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17543 2249 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17625 2249 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17625 2249 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17707 2249 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17707 2249 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17789 2249 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17789 2249 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17871 2249 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17871 2249 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17953 2249 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17953 2249 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 18035 2249 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18035 2249 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 18117 2249 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18117 2249 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 18199 2249 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18199 2249 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 18281 2249 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18281 2249 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 18363 2249 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18363 2249 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 18445 2249 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18445 2249 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 18527 2249 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18527 2249 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2232 3560 2296 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2232 3560 2296 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2232 3646 2296 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2232 3646 2296 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2232 3732 2296 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2232 3732 2296 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2232 3818 2296 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2232 3818 2296 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2232 3904 2296 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2232 3904 2296 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2232 3990 2296 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2232 3990 2296 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2232 4076 2296 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2232 4076 2296 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2232 4162 2296 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2232 4162 2296 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2232 4248 2296 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2232 4248 2296 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2232 4334 2296 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2232 4334 2296 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2232 4420 2296 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2232 4420 2296 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 13613 2301 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 13613 2301 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 13695 2301 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 13695 2301 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 13777 2301 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 13777 2301 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 13859 2301 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 13859 2301 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 13941 2301 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 13941 2301 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14023 2301 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14023 2301 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14105 2301 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14105 2301 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14187 2301 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14187 2301 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14269 2301 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14269 2301 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14351 2301 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14351 2301 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14433 2301 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14433 2301 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14515 2301 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14515 2301 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14597 2301 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14597 2301 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14678 2301 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14678 2301 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14759 2301 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14759 2301 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14840 2301 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14840 2301 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14921 2301 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14921 2301 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15002 2301 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15002 2301 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15083 2301 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15083 2301 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15164 2301 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15164 2301 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15245 2301 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15245 2301 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15326 2301 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15326 2301 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15407 2301 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15407 2301 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15488 2301 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15488 2301 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15569 2301 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15569 2301 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15650 2301 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15650 2301 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15731 2301 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15731 2301 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15812 2301 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15812 2301 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15893 2301 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15893 2301 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15974 2301 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15974 2301 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 16055 2301 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16055 2301 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 16136 2301 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16136 2301 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 16217 2301 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16217 2301 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 16298 2301 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16298 2301 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 16379 2301 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16379 2301 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 16460 2301 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16460 2301 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 16559 2331 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16559 2331 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 16641 2331 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16641 2331 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 16723 2331 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16723 2331 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 16805 2331 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16805 2331 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 16887 2331 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16887 2331 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 16969 2331 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16969 2331 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17051 2331 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17051 2331 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17133 2331 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17133 2331 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17215 2331 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17215 2331 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17297 2331 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17297 2331 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17379 2331 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17379 2331 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17461 2331 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17461 2331 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17543 2331 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17543 2331 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17625 2331 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17625 2331 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17707 2331 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17707 2331 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17789 2331 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17789 2331 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17871 2331 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17871 2331 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17953 2331 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17953 2331 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 18035 2331 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18035 2331 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 18117 2331 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18117 2331 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 18199 2331 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18199 2331 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 18281 2331 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18281 2331 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 18363 2331 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18363 2331 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 18445 2331 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18445 2331 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 18527 2331 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18527 2331 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2313 3560 2377 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2313 3560 2377 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2313 3646 2377 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2313 3646 2377 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2313 3732 2377 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2313 3732 2377 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2313 3818 2377 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2313 3818 2377 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2313 3904 2377 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2313 3904 2377 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2313 3990 2377 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2313 3990 2377 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2313 4076 2377 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2313 4076 2377 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2313 4162 2377 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2313 4162 2377 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2313 4248 2377 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2313 4248 2377 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2313 4334 2377 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2313 4334 2377 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2313 4420 2377 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2313 4420 2377 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 13613 2381 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 13613 2381 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 13695 2381 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 13695 2381 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 13777 2381 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 13777 2381 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 13859 2381 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 13859 2381 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 13941 2381 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 13941 2381 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14023 2381 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14023 2381 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14105 2381 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14105 2381 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14187 2381 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14187 2381 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14269 2381 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14269 2381 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14351 2381 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14351 2381 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14433 2381 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14433 2381 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14515 2381 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14515 2381 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14597 2381 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14597 2381 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14678 2381 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14678 2381 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14759 2381 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14759 2381 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14840 2381 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14840 2381 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14921 2381 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14921 2381 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15002 2381 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15002 2381 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15083 2381 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15083 2381 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15164 2381 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15164 2381 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15245 2381 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15245 2381 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15326 2381 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15326 2381 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15407 2381 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15407 2381 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15488 2381 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15488 2381 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15569 2381 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15569 2381 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15650 2381 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15650 2381 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15731 2381 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15731 2381 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15812 2381 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15812 2381 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15893 2381 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15893 2381 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15974 2381 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15974 2381 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 16055 2381 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16055 2381 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 16136 2381 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16136 2381 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 16217 2381 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16217 2381 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 16298 2381 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16298 2381 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 16379 2381 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16379 2381 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 16460 2381 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16460 2381 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 16559 2413 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16559 2413 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 16641 2413 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16641 2413 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 16723 2413 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16723 2413 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 16805 2413 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16805 2413 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 16887 2413 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16887 2413 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 16969 2413 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16969 2413 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17051 2413 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17051 2413 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17133 2413 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17133 2413 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17215 2413 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17215 2413 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17297 2413 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17297 2413 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17379 2413 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17379 2413 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17461 2413 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17461 2413 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17543 2413 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17543 2413 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17625 2413 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17625 2413 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17707 2413 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17707 2413 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17789 2413 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17789 2413 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17871 2413 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17871 2413 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17953 2413 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17953 2413 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 18035 2413 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18035 2413 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 18117 2413 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18117 2413 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 18199 2413 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18199 2413 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 18281 2413 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18281 2413 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 18363 2413 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18363 2413 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 18445 2413 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18445 2413 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 18527 2413 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18527 2413 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2394 3560 2458 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2394 3560 2458 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2394 3646 2458 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2394 3646 2458 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2394 3732 2458 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2394 3732 2458 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2394 3818 2458 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2394 3818 2458 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2394 3904 2458 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2394 3904 2458 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2394 3990 2458 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2394 3990 2458 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2394 4076 2458 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2394 4076 2458 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2394 4162 2458 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2394 4162 2458 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2394 4248 2458 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2394 4248 2458 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2394 4334 2458 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2394 4334 2458 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2394 4420 2458 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2394 4420 2458 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 13613 2461 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 13613 2461 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 13695 2461 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 13695 2461 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 13777 2461 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 13777 2461 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 13859 2461 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 13859 2461 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 13941 2461 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 13941 2461 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14023 2461 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14023 2461 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14105 2461 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14105 2461 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14187 2461 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14187 2461 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14269 2461 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14269 2461 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14351 2461 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14351 2461 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14433 2461 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14433 2461 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14515 2461 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14515 2461 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14597 2461 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14597 2461 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14678 2461 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14678 2461 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14759 2461 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14759 2461 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14840 2461 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14840 2461 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14921 2461 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14921 2461 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15002 2461 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15002 2461 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15083 2461 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15083 2461 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15164 2461 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15164 2461 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15245 2461 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15245 2461 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15326 2461 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15326 2461 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15407 2461 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15407 2461 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15488 2461 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15488 2461 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15569 2461 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15569 2461 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15650 2461 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15650 2461 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15731 2461 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15731 2461 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15812 2461 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15812 2461 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15893 2461 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15893 2461 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15974 2461 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15974 2461 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 16055 2461 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16055 2461 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 16136 2461 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16136 2461 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 16217 2461 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16217 2461 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 16298 2461 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16298 2461 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 16379 2461 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16379 2461 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 16460 2461 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16460 2461 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 16559 2495 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16559 2495 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 16641 2495 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16641 2495 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 16723 2495 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16723 2495 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 16805 2495 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16805 2495 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 16887 2495 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16887 2495 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 16969 2495 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16969 2495 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17051 2495 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17051 2495 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17133 2495 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17133 2495 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17215 2495 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17215 2495 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17297 2495 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17297 2495 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17379 2495 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17379 2495 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17461 2495 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17461 2495 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17543 2495 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17543 2495 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17625 2495 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17625 2495 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17707 2495 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17707 2495 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17789 2495 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17789 2495 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17871 2495 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17871 2495 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17953 2495 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17953 2495 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 18035 2495 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18035 2495 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 18117 2495 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18117 2495 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 18199 2495 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18199 2495 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 18281 2495 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18281 2495 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 18363 2495 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18363 2495 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 18445 2495 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18445 2495 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 18527 2495 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18527 2495 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2475 3560 2539 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2475 3560 2539 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2475 3646 2539 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2475 3646 2539 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2475 3732 2539 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2475 3732 2539 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2475 3818 2539 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2475 3818 2539 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2475 3904 2539 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2475 3904 2539 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2475 3990 2539 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2475 3990 2539 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2475 4076 2539 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2475 4076 2539 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2475 4162 2539 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2475 4162 2539 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2475 4248 2539 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2475 4248 2539 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2475 4334 2539 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2475 4334 2539 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2475 4420 2539 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2475 4420 2539 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 13613 2541 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 13613 2541 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 13695 2541 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 13695 2541 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 13777 2541 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 13777 2541 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 13859 2541 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 13859 2541 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 13941 2541 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 13941 2541 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14023 2541 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14023 2541 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14105 2541 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14105 2541 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14187 2541 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14187 2541 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14269 2541 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14269 2541 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14351 2541 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14351 2541 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14433 2541 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14433 2541 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14515 2541 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14515 2541 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14597 2541 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14597 2541 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14678 2541 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14678 2541 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14759 2541 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14759 2541 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14840 2541 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14840 2541 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14921 2541 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14921 2541 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15002 2541 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15002 2541 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15083 2541 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15083 2541 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15164 2541 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15164 2541 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15245 2541 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15245 2541 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15326 2541 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15326 2541 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15407 2541 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15407 2541 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15488 2541 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15488 2541 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15569 2541 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15569 2541 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15650 2541 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15650 2541 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15731 2541 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15731 2541 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15812 2541 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15812 2541 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15893 2541 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15893 2541 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15974 2541 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15974 2541 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 16055 2541 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16055 2541 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 16136 2541 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16136 2541 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 16217 2541 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16217 2541 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 16298 2541 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16298 2541 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 16379 2541 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16379 2541 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 16460 2541 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16460 2541 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 16559 2577 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16559 2577 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 16641 2577 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16641 2577 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 16723 2577 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16723 2577 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 16805 2577 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16805 2577 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 16887 2577 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16887 2577 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 16969 2577 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16969 2577 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17051 2577 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17051 2577 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17133 2577 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17133 2577 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17215 2577 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17215 2577 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17297 2577 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17297 2577 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17379 2577 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17379 2577 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17461 2577 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17461 2577 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17543 2577 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17543 2577 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17625 2577 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17625 2577 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17707 2577 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17707 2577 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17789 2577 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17789 2577 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17871 2577 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17871 2577 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17953 2577 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17953 2577 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 18035 2577 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18035 2577 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 18117 2577 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18117 2577 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 18199 2577 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18199 2577 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 18281 2577 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18281 2577 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 18363 2577 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18363 2577 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 18445 2577 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18445 2577 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 18527 2577 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18527 2577 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2556 3560 2620 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2556 3560 2620 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2556 3646 2620 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2556 3646 2620 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2556 3732 2620 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2556 3732 2620 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2556 3818 2620 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2556 3818 2620 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2556 3904 2620 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2556 3904 2620 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2556 3990 2620 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2556 3990 2620 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2556 4076 2620 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2556 4076 2620 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2556 4162 2620 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2556 4162 2620 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2556 4248 2620 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2556 4248 2620 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2556 4334 2620 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2556 4334 2620 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2556 4420 2620 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2556 4420 2620 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 13613 2621 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 13613 2621 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 13695 2621 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 13695 2621 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 13777 2621 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 13777 2621 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 13859 2621 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 13859 2621 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 13941 2621 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 13941 2621 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14023 2621 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14023 2621 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14105 2621 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14105 2621 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14187 2621 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14187 2621 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14269 2621 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14269 2621 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14351 2621 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14351 2621 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14433 2621 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14433 2621 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14515 2621 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14515 2621 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14597 2621 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14597 2621 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14678 2621 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14678 2621 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14759 2621 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14759 2621 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14840 2621 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14840 2621 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14921 2621 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14921 2621 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15002 2621 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15002 2621 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15083 2621 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15083 2621 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15164 2621 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15164 2621 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15245 2621 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15245 2621 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15326 2621 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15326 2621 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15407 2621 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15407 2621 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15488 2621 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15488 2621 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15569 2621 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15569 2621 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15650 2621 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15650 2621 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15731 2621 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15731 2621 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15812 2621 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15812 2621 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15893 2621 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15893 2621 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15974 2621 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15974 2621 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 16055 2621 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16055 2621 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 16136 2621 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16136 2621 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 16217 2621 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16217 2621 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 16298 2621 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16298 2621 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 16379 2621 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16379 2621 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 16460 2621 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16460 2621 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 16559 2658 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16559 2658 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 16641 2658 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16641 2658 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 16723 2658 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16723 2658 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 16805 2658 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16805 2658 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 16887 2658 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16887 2658 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 16969 2658 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16969 2658 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17051 2658 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17051 2658 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17133 2658 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17133 2658 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17215 2658 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17215 2658 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17297 2658 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17297 2658 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17379 2658 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17379 2658 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17461 2658 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17461 2658 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17543 2658 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17543 2658 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17625 2658 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17625 2658 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17707 2658 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17707 2658 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17789 2658 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17789 2658 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17871 2658 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17871 2658 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17953 2658 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17953 2658 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 18035 2658 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18035 2658 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 18117 2658 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18117 2658 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 18199 2658 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18199 2658 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 18281 2658 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18281 2658 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 18363 2658 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18363 2658 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 18445 2658 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18445 2658 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 18527 2658 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18527 2658 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 3560 2701 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 3560 2701 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 3646 2701 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 3646 2701 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 3732 2701 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 3732 2701 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 3818 2701 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 3818 2701 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 3904 2701 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 3904 2701 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 3990 2701 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 3990 2701 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 4076 2701 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 4076 2701 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 4162 2701 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 4162 2701 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 4248 2701 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 4248 2701 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 4334 2701 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 4334 2701 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 4420 2701 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 4420 2701 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 13613 2701 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 13613 2701 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 13695 2701 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 13695 2701 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 13777 2701 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 13777 2701 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 13859 2701 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 13859 2701 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 13941 2701 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 13941 2701 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14023 2701 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14023 2701 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14105 2701 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14105 2701 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14187 2701 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14187 2701 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14269 2701 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14269 2701 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14351 2701 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14351 2701 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14433 2701 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14433 2701 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14515 2701 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14515 2701 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14597 2701 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14597 2701 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14678 2701 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14678 2701 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14759 2701 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14759 2701 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14840 2701 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14840 2701 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14921 2701 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14921 2701 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15002 2701 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15002 2701 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15083 2701 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15083 2701 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15164 2701 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15164 2701 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15245 2701 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15245 2701 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15326 2701 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15326 2701 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15407 2701 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15407 2701 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15488 2701 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15488 2701 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15569 2701 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15569 2701 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15650 2701 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15650 2701 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15731 2701 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15731 2701 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15812 2701 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15812 2701 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15893 2701 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15893 2701 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15974 2701 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15974 2701 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 16055 2701 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16055 2701 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 16136 2701 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16136 2701 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 16217 2701 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16217 2701 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 16298 2701 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16298 2701 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 16379 2701 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16379 2701 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 16460 2701 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16460 2701 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 16559 2739 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16559 2739 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 16641 2739 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16641 2739 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 16723 2739 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16723 2739 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 16805 2739 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16805 2739 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 16887 2739 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16887 2739 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 16969 2739 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16969 2739 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17051 2739 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17051 2739 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17133 2739 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17133 2739 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17215 2739 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17215 2739 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17297 2739 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17297 2739 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17379 2739 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17379 2739 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17461 2739 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17461 2739 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17543 2739 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17543 2739 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17625 2739 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17625 2739 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17707 2739 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17707 2739 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17789 2739 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17789 2739 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17871 2739 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17871 2739 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17953 2739 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17953 2739 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 18035 2739 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18035 2739 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 18117 2739 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18117 2739 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 18199 2739 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18199 2739 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 18281 2739 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18281 2739 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 18363 2739 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18363 2739 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 18445 2739 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18445 2739 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 18527 2739 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18527 2739 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 13613 2781 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 13613 2781 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 13695 2781 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 13695 2781 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 13777 2781 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 13777 2781 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 13859 2781 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 13859 2781 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 13941 2781 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 13941 2781 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14023 2781 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14023 2781 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14105 2781 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14105 2781 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14187 2781 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14187 2781 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14269 2781 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14269 2781 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14351 2781 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14351 2781 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14433 2781 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14433 2781 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14515 2781 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14515 2781 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14597 2781 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14597 2781 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14678 2781 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14678 2781 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14759 2781 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14759 2781 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14840 2781 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14840 2781 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14921 2781 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14921 2781 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15002 2781 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15002 2781 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15083 2781 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15083 2781 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15164 2781 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15164 2781 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15245 2781 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15245 2781 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15326 2781 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15326 2781 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15407 2781 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15407 2781 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15488 2781 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15488 2781 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15569 2781 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15569 2781 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15650 2781 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15650 2781 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15731 2781 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15731 2781 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15812 2781 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15812 2781 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15893 2781 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15893 2781 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15974 2781 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15974 2781 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 16055 2781 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16055 2781 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 16136 2781 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16136 2781 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 16217 2781 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16217 2781 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 16298 2781 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16298 2781 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 16379 2781 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16379 2781 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 16460 2781 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16460 2781 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2718 3560 2782 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2718 3560 2782 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2718 3646 2782 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2718 3646 2782 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2718 3732 2782 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2718 3732 2782 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2718 3818 2782 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2718 3818 2782 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2718 3904 2782 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2718 3904 2782 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2718 3990 2782 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2718 3990 2782 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2718 4076 2782 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2718 4076 2782 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2718 4162 2782 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2718 4162 2782 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2718 4248 2782 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2718 4248 2782 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2718 4334 2782 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2718 4334 2782 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2718 4420 2782 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2718 4420 2782 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 16559 2820 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16559 2820 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 16641 2820 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16641 2820 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 16723 2820 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16723 2820 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 16805 2820 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16805 2820 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 16887 2820 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16887 2820 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 16969 2820 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16969 2820 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17051 2820 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17051 2820 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17133 2820 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17133 2820 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17215 2820 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17215 2820 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17297 2820 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17297 2820 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17379 2820 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17379 2820 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17461 2820 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17461 2820 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17543 2820 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17543 2820 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17625 2820 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17625 2820 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17707 2820 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17707 2820 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17789 2820 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17789 2820 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17871 2820 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17871 2820 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17953 2820 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17953 2820 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 18035 2820 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18035 2820 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 18117 2820 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18117 2820 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 18199 2820 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18199 2820 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 18281 2820 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18281 2820 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 18363 2820 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18363 2820 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 18445 2820 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18445 2820 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 18527 2820 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18527 2820 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 13613 2861 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 13613 2861 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 13695 2861 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 13695 2861 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 13777 2861 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 13777 2861 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 13859 2861 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 13859 2861 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 13941 2861 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 13941 2861 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14023 2861 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14023 2861 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14105 2861 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14105 2861 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14187 2861 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14187 2861 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14269 2861 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14269 2861 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14351 2861 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14351 2861 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14433 2861 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14433 2861 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14515 2861 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14515 2861 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14597 2861 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14597 2861 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14678 2861 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14678 2861 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14759 2861 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14759 2861 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14840 2861 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14840 2861 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14921 2861 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14921 2861 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15002 2861 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15002 2861 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15083 2861 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15083 2861 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15164 2861 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15164 2861 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15245 2861 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15245 2861 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15326 2861 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15326 2861 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15407 2861 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15407 2861 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15488 2861 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15488 2861 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15569 2861 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15569 2861 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15650 2861 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15650 2861 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15731 2861 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15731 2861 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15812 2861 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15812 2861 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15893 2861 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15893 2861 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15974 2861 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15974 2861 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 16055 2861 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16055 2861 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 16136 2861 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16136 2861 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 16217 2861 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16217 2861 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 16298 2861 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16298 2861 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 16379 2861 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16379 2861 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 16460 2861 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16460 2861 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2799 3560 2863 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2799 3560 2863 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2799 3646 2863 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2799 3646 2863 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2799 3732 2863 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2799 3732 2863 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2799 3818 2863 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2799 3818 2863 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2799 3904 2863 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2799 3904 2863 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2799 3990 2863 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2799 3990 2863 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2799 4076 2863 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2799 4076 2863 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2799 4162 2863 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2799 4162 2863 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2799 4248 2863 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2799 4248 2863 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2799 4334 2863 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2799 4334 2863 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2799 4420 2863 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2799 4420 2863 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2852 18191 2916 18255 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2852 18191 2916 18255 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2852 18277 2916 18341 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2852 18277 2916 18341 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2856 17670 2920 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 17670 2920 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2856 17755 2920 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 17755 2920 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2856 17841 2920 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 17841 2920 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2856 17927 2920 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 17927 2920 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2856 18013 2920 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 18013 2920 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2856 18099 2920 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 18099 2920 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 13613 2941 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 13613 2941 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 13695 2941 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 13695 2941 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 13777 2941 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 13777 2941 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 13859 2941 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 13859 2941 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 13941 2941 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 13941 2941 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14023 2941 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14023 2941 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14105 2941 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14105 2941 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14187 2941 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14187 2941 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14269 2941 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14269 2941 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14351 2941 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14351 2941 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14433 2941 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14433 2941 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14515 2941 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14515 2941 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14597 2941 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14597 2941 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14678 2941 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14678 2941 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14759 2941 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14759 2941 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14840 2941 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14840 2941 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14921 2941 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14921 2941 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15002 2941 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15002 2941 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15083 2941 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15083 2941 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15164 2941 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15164 2941 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15245 2941 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15245 2941 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15326 2941 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15326 2941 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15407 2941 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15407 2941 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15488 2941 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15488 2941 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15569 2941 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15569 2941 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15650 2941 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15650 2941 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15731 2941 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15731 2941 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15812 2941 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15812 2941 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15893 2941 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15893 2941 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15974 2941 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15974 2941 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 16055 2941 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16055 2941 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 16136 2941 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16136 2941 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 16217 2941 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16217 2941 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 16298 2941 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16298 2941 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 16379 2941 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16379 2941 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 16460 2941 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16460 2941 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2880 3560 2944 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2880 3560 2944 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2880 3646 2944 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2880 3646 2944 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2880 3732 2944 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2880 3732 2944 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2880 3818 2944 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2880 3818 2944 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2880 3904 2944 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2880 3904 2944 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2880 3990 2944 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2880 3990 2944 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2880 4076 2944 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2880 4076 2944 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2880 4162 2944 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2880 4162 2944 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2880 4248 2944 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2880 4248 2944 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2880 4334 2944 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2880 4334 2944 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2880 4420 2944 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2880 4420 2944 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2881 16599 2945 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16599 2945 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2881 16679 2945 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16679 2945 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2881 16759 2945 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16759 2945 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2881 16839 2945 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16839 2945 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2881 16919 2945 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16919 2945 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2881 16999 2945 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16999 2945 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2881 17079 2945 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17079 2945 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2881 17159 2945 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17159 2945 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2881 17239 2945 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17239 2945 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2881 17320 2945 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17320 2945 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2881 17401 2945 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17401 2945 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2881 17482 2945 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17482 2945 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2881 17563 2945 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17563 2945 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2938 17670 3002 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 17670 3002 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2938 17755 3002 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 17755 3002 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2938 17841 3002 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 17841 3002 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2938 17927 3002 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 17927 3002 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2938 18013 3002 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 18013 3002 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2938 18099 3002 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 18099 3002 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 13613 3021 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 13613 3021 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 13695 3021 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 13695 3021 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 13777 3021 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 13777 3021 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 13859 3021 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 13859 3021 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 13941 3021 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 13941 3021 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14023 3021 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14023 3021 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14105 3021 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14105 3021 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14187 3021 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14187 3021 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14269 3021 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14269 3021 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14351 3021 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14351 3021 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14433 3021 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14433 3021 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14515 3021 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14515 3021 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14597 3021 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14597 3021 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14678 3021 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14678 3021 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14759 3021 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14759 3021 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14840 3021 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14840 3021 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14921 3021 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14921 3021 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15002 3021 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15002 3021 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15083 3021 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15083 3021 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15164 3021 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15164 3021 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15245 3021 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15245 3021 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15326 3021 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15326 3021 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15407 3021 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15407 3021 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15488 3021 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15488 3021 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15569 3021 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15569 3021 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15650 3021 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15650 3021 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15731 3021 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15731 3021 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15812 3021 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15812 3021 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15893 3021 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15893 3021 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15974 3021 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15974 3021 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 16055 3021 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16055 3021 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 16136 3021 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16136 3021 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 16217 3021 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16217 3021 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 16298 3021 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16298 3021 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 16379 3021 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16379 3021 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 16460 3021 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16460 3021 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2961 3560 3025 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2961 3560 3025 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2961 3646 3025 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2961 3646 3025 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2961 3732 3025 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2961 3732 3025 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2961 3818 3025 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2961 3818 3025 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2961 3904 3025 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2961 3904 3025 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2961 3990 3025 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2961 3990 3025 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2961 4076 3025 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2961 4076 3025 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2961 4162 3025 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2961 4162 3025 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2961 4248 3025 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2961 4248 3025 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2961 4334 3025 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2961 4334 3025 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2961 4420 3025 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2961 4420 3025 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2963 16599 3027 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16599 3027 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2963 16679 3027 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16679 3027 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2963 16759 3027 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16759 3027 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2963 16839 3027 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16839 3027 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2963 16919 3027 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16919 3027 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2963 16999 3027 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16999 3027 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2963 17079 3027 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17079 3027 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2963 17159 3027 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17159 3027 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2963 17239 3027 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17239 3027 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2963 17320 3027 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17320 3027 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2963 17401 3027 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17401 3027 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2963 17482 3027 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17482 3027 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2963 17563 3027 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17563 3027 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3008 18191 3072 18255 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3008 18191 3072 18255 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3008 18277 3072 18341 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3008 18277 3072 18341 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3020 17670 3084 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 17670 3084 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3020 17755 3084 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 17755 3084 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3020 17841 3084 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 17841 3084 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3020 17927 3084 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 17927 3084 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3020 18013 3084 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 18013 3084 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3020 18099 3084 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 18099 3084 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 13613 3101 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 13613 3101 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 13695 3101 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 13695 3101 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 13777 3101 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 13777 3101 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 13859 3101 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 13859 3101 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 13941 3101 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 13941 3101 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14023 3101 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14023 3101 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14105 3101 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14105 3101 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14187 3101 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14187 3101 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14269 3101 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14269 3101 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14351 3101 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14351 3101 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14433 3101 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14433 3101 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14515 3101 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14515 3101 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14597 3101 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14597 3101 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14678 3101 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14678 3101 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14759 3101 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14759 3101 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14840 3101 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14840 3101 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14921 3101 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14921 3101 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15002 3101 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15002 3101 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15083 3101 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15083 3101 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15164 3101 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15164 3101 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15245 3101 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15245 3101 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15326 3101 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15326 3101 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15407 3101 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15407 3101 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15488 3101 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15488 3101 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15569 3101 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15569 3101 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15650 3101 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15650 3101 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15731 3101 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15731 3101 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15812 3101 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15812 3101 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15893 3101 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15893 3101 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15974 3101 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15974 3101 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 16055 3101 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16055 3101 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 16136 3101 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16136 3101 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 16217 3101 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16217 3101 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 16298 3101 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16298 3101 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 16379 3101 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16379 3101 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 16460 3101 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16460 3101 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3042 3560 3106 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3042 3560 3106 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3042 3646 3106 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3042 3646 3106 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3042 3732 3106 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3042 3732 3106 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3042 3818 3106 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3042 3818 3106 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3042 3904 3106 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3042 3904 3106 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3042 3990 3106 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3042 3990 3106 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3042 4076 3106 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3042 4076 3106 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3042 4162 3106 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3042 4162 3106 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3042 4248 3106 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3042 4248 3106 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3042 4334 3106 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3042 4334 3106 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3042 4420 3106 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3042 4420 3106 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3045 16599 3109 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16599 3109 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3045 16679 3109 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16679 3109 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3045 16759 3109 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16759 3109 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3045 16839 3109 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16839 3109 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3045 16919 3109 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16919 3109 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3045 16999 3109 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16999 3109 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3045 17079 3109 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17079 3109 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3045 17159 3109 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17159 3109 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3045 17239 3109 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17239 3109 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3045 17320 3109 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17320 3109 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3045 17401 3109 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17401 3109 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3045 17482 3109 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17482 3109 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3045 17563 3109 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17563 3109 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3102 17670 3166 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 17670 3166 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3102 17755 3166 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 17755 3166 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3102 17841 3166 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 17841 3166 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3102 17927 3166 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 17927 3166 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3102 18013 3166 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 18013 3166 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3102 18099 3166 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 18099 3166 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 13613 3181 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 13613 3181 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 13695 3181 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 13695 3181 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 13777 3181 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 13777 3181 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 13859 3181 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 13859 3181 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 13941 3181 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 13941 3181 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14023 3181 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14023 3181 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14105 3181 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14105 3181 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14187 3181 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14187 3181 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14269 3181 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14269 3181 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14351 3181 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14351 3181 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14433 3181 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14433 3181 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14515 3181 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14515 3181 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14597 3181 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14597 3181 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14678 3181 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14678 3181 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14759 3181 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14759 3181 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14840 3181 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14840 3181 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14921 3181 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14921 3181 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15002 3181 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15002 3181 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15083 3181 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15083 3181 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15164 3181 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15164 3181 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15245 3181 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15245 3181 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15326 3181 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15326 3181 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15407 3181 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15407 3181 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15488 3181 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15488 3181 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15569 3181 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15569 3181 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15650 3181 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15650 3181 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15731 3181 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15731 3181 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15812 3181 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15812 3181 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15893 3181 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15893 3181 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15974 3181 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15974 3181 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 16055 3181 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16055 3181 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 16136 3181 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16136 3181 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 16217 3181 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16217 3181 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 16298 3181 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16298 3181 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 16379 3181 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16379 3181 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 16460 3181 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16460 3181 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3123 3560 3187 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3123 3560 3187 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3123 3646 3187 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3123 3646 3187 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3123 3732 3187 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3123 3732 3187 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3123 3818 3187 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3123 3818 3187 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3123 3904 3187 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3123 3904 3187 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3123 3990 3187 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3123 3990 3187 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3123 4076 3187 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3123 4076 3187 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3123 4162 3187 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3123 4162 3187 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3123 4248 3187 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3123 4248 3187 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3123 4334 3187 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3123 4334 3187 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3123 4420 3187 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3123 4420 3187 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3127 16599 3191 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16599 3191 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3127 16679 3191 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16679 3191 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3127 16759 3191 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16759 3191 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3127 16839 3191 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16839 3191 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3127 16919 3191 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16919 3191 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3127 16999 3191 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16999 3191 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3127 17079 3191 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17079 3191 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3127 17159 3191 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17159 3191 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3127 17239 3191 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17239 3191 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3127 17320 3191 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17320 3191 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3127 17401 3191 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17401 3191 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3127 17482 3191 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17482 3191 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3127 17563 3191 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17563 3191 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3184 17670 3248 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 17670 3248 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3184 17755 3248 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 17755 3248 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3184 17841 3248 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 17841 3248 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3184 17927 3248 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 17927 3248 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3184 18013 3248 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 18013 3248 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3184 18099 3248 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 18099 3248 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 13613 3261 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 13613 3261 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 13695 3261 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 13695 3261 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 13777 3261 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 13777 3261 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 13859 3261 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 13859 3261 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 13941 3261 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 13941 3261 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14023 3261 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14023 3261 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14105 3261 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14105 3261 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14187 3261 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14187 3261 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14269 3261 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14269 3261 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14351 3261 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14351 3261 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14433 3261 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14433 3261 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14515 3261 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14515 3261 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14597 3261 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14597 3261 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14678 3261 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14678 3261 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14759 3261 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14759 3261 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14840 3261 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14840 3261 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14921 3261 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14921 3261 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15002 3261 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15002 3261 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15083 3261 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15083 3261 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15164 3261 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15164 3261 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15245 3261 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15245 3261 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15326 3261 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15326 3261 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15407 3261 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15407 3261 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15488 3261 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15488 3261 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15569 3261 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15569 3261 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15650 3261 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15650 3261 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15731 3261 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15731 3261 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15812 3261 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15812 3261 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15893 3261 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15893 3261 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15974 3261 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15974 3261 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 16055 3261 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16055 3261 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 16136 3261 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16136 3261 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 16217 3261 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16217 3261 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 16298 3261 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16298 3261 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 16379 3261 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16379 3261 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 16460 3261 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16460 3261 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3204 3560 3268 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3204 3560 3268 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3204 3646 3268 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3204 3646 3268 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3204 3732 3268 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3204 3732 3268 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3204 3818 3268 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3204 3818 3268 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3204 3904 3268 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3204 3904 3268 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3204 3990 3268 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3204 3990 3268 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3204 4076 3268 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3204 4076 3268 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3204 4162 3268 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3204 4162 3268 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3204 4248 3268 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3204 4248 3268 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3204 4334 3268 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3204 4334 3268 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3204 4420 3268 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3204 4420 3268 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3209 16599 3273 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16599 3273 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3209 16679 3273 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16679 3273 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3209 16759 3273 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16759 3273 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3209 16839 3273 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16839 3273 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3209 16919 3273 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16919 3273 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3209 16999 3273 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16999 3273 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3209 17079 3273 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17079 3273 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3209 17159 3273 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17159 3273 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3209 17239 3273 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17239 3273 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3209 17320 3273 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17320 3273 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3209 17401 3273 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17401 3273 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3209 17482 3273 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17482 3273 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3209 17563 3273 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17563 3273 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 13613 3341 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 13613 3341 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 13695 3341 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 13695 3341 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 13777 3341 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 13777 3341 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 13859 3341 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 13859 3341 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 13941 3341 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 13941 3341 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14023 3341 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14023 3341 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14105 3341 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14105 3341 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14187 3341 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14187 3341 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14269 3341 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14269 3341 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14351 3341 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14351 3341 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14433 3341 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14433 3341 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14515 3341 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14515 3341 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14597 3341 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14597 3341 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14678 3341 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14678 3341 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14759 3341 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14759 3341 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14840 3341 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14840 3341 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14921 3341 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14921 3341 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15002 3341 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15002 3341 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15083 3341 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15083 3341 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15164 3341 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15164 3341 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15245 3341 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15245 3341 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15326 3341 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15326 3341 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15407 3341 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15407 3341 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15488 3341 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15488 3341 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15569 3341 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15569 3341 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15650 3341 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15650 3341 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15731 3341 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15731 3341 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15812 3341 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15812 3341 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15893 3341 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15893 3341 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15974 3341 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15974 3341 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 16055 3341 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16055 3341 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 16136 3341 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16136 3341 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 16217 3341 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16217 3341 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 16298 3341 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16298 3341 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 16379 3341 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16379 3341 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 16460 3341 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16460 3341 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3284 17674 3348 17738 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3284 17674 3348 17738 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3284 17757 3348 17821 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3284 17757 3348 17821 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3284 17841 3348 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3284 17841 3348 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3285 3560 3349 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3285 3560 3349 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3285 3646 3349 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3285 3646 3349 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3285 3732 3349 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3285 3732 3349 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3285 3818 3349 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3285 3818 3349 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3285 3904 3349 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3285 3904 3349 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3285 3990 3349 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3285 3990 3349 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3285 4076 3349 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3285 4076 3349 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3285 4162 3349 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3285 4162 3349 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3285 4248 3349 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3285 4248 3349 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3285 4334 3349 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3285 4334 3349 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3285 4420 3349 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3285 4420 3349 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3291 16599 3355 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16599 3355 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3291 16679 3355 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16679 3355 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3291 16759 3355 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16759 3355 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3291 16839 3355 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16839 3355 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3291 16919 3355 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16919 3355 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3291 16999 3355 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16999 3355 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3291 17079 3355 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17079 3355 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3291 17159 3355 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17159 3355 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3291 17239 3355 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17239 3355 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3291 17320 3355 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17320 3355 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3291 17401 3355 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17401 3355 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3291 17482 3355 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17482 3355 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3291 17563 3355 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17563 3355 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 13613 3421 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 13613 3421 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 13695 3421 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 13695 3421 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 13777 3421 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 13777 3421 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 13859 3421 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 13859 3421 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 13941 3421 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 13941 3421 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14023 3421 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14023 3421 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14105 3421 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14105 3421 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14187 3421 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14187 3421 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14269 3421 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14269 3421 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14351 3421 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14351 3421 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14433 3421 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14433 3421 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14515 3421 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14515 3421 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14597 3421 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14597 3421 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14678 3421 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14678 3421 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14759 3421 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14759 3421 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14840 3421 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14840 3421 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14921 3421 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14921 3421 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15002 3421 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15002 3421 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15083 3421 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15083 3421 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15164 3421 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15164 3421 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15245 3421 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15245 3421 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15326 3421 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15326 3421 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15407 3421 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15407 3421 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15488 3421 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15488 3421 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15569 3421 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15569 3421 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15650 3421 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15650 3421 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15731 3421 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15731 3421 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15812 3421 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15812 3421 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15893 3421 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15893 3421 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15974 3421 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15974 3421 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 16055 3421 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16055 3421 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 16136 3421 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16136 3421 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 16217 3421 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16217 3421 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 16298 3421 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16298 3421 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 16379 3421 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16379 3421 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 16460 3421 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16460 3421 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3366 3560 3430 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3366 3560 3430 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3366 3646 3430 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3366 3646 3430 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3366 3732 3430 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3366 3732 3430 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3366 3818 3430 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3366 3818 3430 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3366 3904 3430 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3366 3904 3430 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3366 3990 3430 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3366 3990 3430 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3366 4076 3430 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3366 4076 3430 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3366 4162 3430 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3366 4162 3430 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3366 4248 3430 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3366 4248 3430 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3366 4334 3430 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3366 4334 3430 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3366 4420 3430 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3366 4420 3430 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3373 16599 3437 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16599 3437 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3373 16679 3437 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16679 3437 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3373 16759 3437 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16759 3437 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3373 16839 3437 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16839 3437 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3373 16919 3437 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16919 3437 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3373 16999 3437 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16999 3437 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3373 17079 3437 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17079 3437 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3373 17159 3437 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17159 3437 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3373 17239 3437 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17239 3437 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3373 17320 3437 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17320 3437 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3373 17401 3437 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17401 3437 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3373 17482 3437 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17482 3437 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3373 17563 3437 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17563 3437 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 13613 3501 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 13613 3501 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 13695 3501 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 13695 3501 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 13777 3501 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 13777 3501 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 13859 3501 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 13859 3501 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 13941 3501 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 13941 3501 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14023 3501 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14023 3501 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14105 3501 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14105 3501 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14187 3501 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14187 3501 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14269 3501 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14269 3501 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14351 3501 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14351 3501 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14433 3501 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14433 3501 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14515 3501 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14515 3501 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14597 3501 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14597 3501 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14678 3501 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14678 3501 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14759 3501 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14759 3501 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14840 3501 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14840 3501 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14921 3501 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14921 3501 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15002 3501 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15002 3501 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15083 3501 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15083 3501 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15164 3501 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15164 3501 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15245 3501 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15245 3501 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15326 3501 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15326 3501 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15407 3501 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15407 3501 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15488 3501 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15488 3501 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15569 3501 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15569 3501 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15650 3501 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15650 3501 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15731 3501 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15731 3501 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15812 3501 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15812 3501 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15893 3501 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15893 3501 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15974 3501 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15974 3501 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 16055 3501 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16055 3501 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 16136 3501 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16136 3501 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 16217 3501 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16217 3501 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 16298 3501 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16298 3501 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 16379 3501 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16379 3501 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 16460 3501 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16460 3501 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3440 17674 3504 17738 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3440 17674 3504 17738 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3440 17757 3504 17821 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3440 17757 3504 17821 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3440 17841 3504 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3440 17841 3504 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3447 3560 3511 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3447 3560 3511 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3447 3646 3511 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3447 3646 3511 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3447 3732 3511 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3447 3732 3511 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3447 3818 3511 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3447 3818 3511 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3447 3904 3511 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3447 3904 3511 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3447 3990 3511 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3447 3990 3511 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3447 4076 3511 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3447 4076 3511 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3447 4162 3511 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3447 4162 3511 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3447 4248 3511 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3447 4248 3511 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3447 4334 3511 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3447 4334 3511 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3447 4420 3511 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3447 4420 3511 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3455 16599 3519 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16599 3519 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3455 16679 3519 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16679 3519 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3455 16759 3519 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16759 3519 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3455 16839 3519 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16839 3519 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3455 16919 3519 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16919 3519 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3455 16999 3519 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16999 3519 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3455 17079 3519 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17079 3519 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3455 17159 3519 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17159 3519 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3455 17239 3519 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17239 3519 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3455 17320 3519 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17320 3519 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3455 17401 3519 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17401 3519 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3455 17482 3519 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17482 3519 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3455 17563 3519 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17563 3519 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 13613 3581 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 13613 3581 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 13695 3581 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 13695 3581 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 13777 3581 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 13777 3581 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 13859 3581 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 13859 3581 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 13941 3581 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 13941 3581 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14023 3581 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14023 3581 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14105 3581 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14105 3581 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14187 3581 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14187 3581 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14269 3581 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14269 3581 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14351 3581 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14351 3581 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14433 3581 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14433 3581 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14515 3581 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14515 3581 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14597 3581 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14597 3581 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14678 3581 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14678 3581 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14759 3581 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14759 3581 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14840 3581 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14840 3581 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14921 3581 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14921 3581 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15002 3581 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15002 3581 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15083 3581 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15083 3581 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15164 3581 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15164 3581 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15245 3581 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15245 3581 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15326 3581 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15326 3581 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15407 3581 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15407 3581 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15488 3581 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15488 3581 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15569 3581 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15569 3581 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15650 3581 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15650 3581 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15731 3581 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15731 3581 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15812 3581 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15812 3581 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15893 3581 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15893 3581 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15974 3581 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15974 3581 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 16055 3581 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16055 3581 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 16136 3581 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16136 3581 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 16217 3581 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16217 3581 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 16298 3581 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16298 3581 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 16379 3581 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16379 3581 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 16460 3581 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16460 3581 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3528 3560 3592 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3528 3560 3592 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3528 3646 3592 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3528 3646 3592 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3528 3732 3592 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3528 3732 3592 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3528 3818 3592 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3528 3818 3592 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3528 3904 3592 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3528 3904 3592 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3528 3990 3592 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3528 3990 3592 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3528 4076 3592 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3528 4076 3592 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3528 4162 3592 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3528 4162 3592 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3528 4248 3592 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3528 4248 3592 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3528 4334 3592 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3528 4334 3592 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3528 4420 3592 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3528 4420 3592 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3537 16599 3601 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16599 3601 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3537 16679 3601 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16679 3601 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3537 16759 3601 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16759 3601 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3537 16839 3601 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16839 3601 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3537 16919 3601 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16919 3601 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3537 16999 3601 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16999 3601 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3537 17079 3601 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17079 3601 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3537 17159 3601 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17159 3601 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3537 17239 3601 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17239 3601 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3537 17320 3601 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17320 3601 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3537 17401 3601 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17401 3601 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3537 17482 3601 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17482 3601 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3537 17563 3601 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17563 3601 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 13613 3661 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 13613 3661 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 13695 3661 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 13695 3661 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 13777 3661 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 13777 3661 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 13859 3661 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 13859 3661 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 13941 3661 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 13941 3661 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14023 3661 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14023 3661 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14105 3661 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14105 3661 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14187 3661 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14187 3661 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14269 3661 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14269 3661 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14351 3661 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14351 3661 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14433 3661 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14433 3661 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14515 3661 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14515 3661 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14597 3661 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14597 3661 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14678 3661 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14678 3661 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14759 3661 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14759 3661 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14840 3661 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14840 3661 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14921 3661 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14921 3661 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15002 3661 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15002 3661 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15083 3661 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15083 3661 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15164 3661 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15164 3661 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15245 3661 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15245 3661 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15326 3661 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15326 3661 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15407 3661 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15407 3661 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15488 3661 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15488 3661 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15569 3661 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15569 3661 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15650 3661 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15650 3661 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15731 3661 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15731 3661 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15812 3661 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15812 3661 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15893 3661 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15893 3661 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15974 3661 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15974 3661 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 16055 3661 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16055 3661 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 16136 3661 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16136 3661 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 16217 3661 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16217 3661 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 16298 3661 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16298 3661 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 16379 3661 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16379 3661 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 16460 3661 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16460 3661 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3609 3560 3673 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 3560 3673 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3609 3646 3673 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 3646 3673 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3609 3732 3673 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 3732 3673 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3609 3818 3673 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 3818 3673 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3609 3904 3673 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 3904 3673 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3609 3990 3673 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 3990 3673 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3609 4076 3673 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 4076 3673 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3609 4162 3673 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 4162 3673 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3609 4248 3673 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 4248 3673 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3609 4334 3673 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 4334 3673 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3609 4420 3673 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 4420 3673 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3619 16599 3683 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16599 3683 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3619 16679 3683 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16679 3683 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3619 16759 3683 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16759 3683 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3619 16839 3683 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16839 3683 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3619 16919 3683 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16919 3683 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3619 16999 3683 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16999 3683 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3619 17079 3683 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17079 3683 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3619 17159 3683 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17159 3683 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3619 17239 3683 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17239 3683 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3619 17320 3683 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17320 3683 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3619 17401 3683 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17401 3683 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3619 17482 3683 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17482 3683 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3619 17563 3683 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17563 3683 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 13613 3741 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 13613 3741 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 13695 3741 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 13695 3741 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 13777 3741 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 13777 3741 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 13859 3741 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 13859 3741 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 13941 3741 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 13941 3741 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14023 3741 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14023 3741 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14105 3741 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14105 3741 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14187 3741 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14187 3741 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14269 3741 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14269 3741 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14351 3741 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14351 3741 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14433 3741 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14433 3741 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14515 3741 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14515 3741 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14597 3741 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14597 3741 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14678 3741 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14678 3741 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14759 3741 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14759 3741 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14840 3741 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14840 3741 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14921 3741 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14921 3741 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15002 3741 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15002 3741 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15083 3741 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15083 3741 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15164 3741 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15164 3741 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15245 3741 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15245 3741 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15326 3741 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15326 3741 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15407 3741 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15407 3741 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15488 3741 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15488 3741 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15569 3741 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15569 3741 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15650 3741 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15650 3741 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15731 3741 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15731 3741 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15812 3741 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15812 3741 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15893 3741 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15893 3741 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15974 3741 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15974 3741 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 16055 3741 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16055 3741 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 16136 3741 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16136 3741 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 16217 3741 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16217 3741 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 16298 3741 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16298 3741 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 16379 3741 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16379 3741 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 16460 3741 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16460 3741 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3690 3560 3754 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3690 3560 3754 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3690 3646 3754 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3690 3646 3754 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3690 3732 3754 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3690 3732 3754 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3690 3818 3754 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3690 3818 3754 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3690 3904 3754 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3690 3904 3754 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3690 3990 3754 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3690 3990 3754 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3690 4076 3754 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3690 4076 3754 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3690 4162 3754 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3690 4162 3754 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3690 4248 3754 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3690 4248 3754 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3690 4334 3754 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3690 4334 3754 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3690 4420 3754 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3690 4420 3754 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3701 16599 3765 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16599 3765 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3701 16679 3765 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16679 3765 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3701 16759 3765 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16759 3765 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3701 16839 3765 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16839 3765 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3701 16919 3765 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16919 3765 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3701 16999 3765 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16999 3765 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3701 17079 3765 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17079 3765 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3701 17159 3765 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17159 3765 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3701 17239 3765 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17239 3765 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3701 17320 3765 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17320 3765 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3701 17401 3765 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17401 3765 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3701 17482 3765 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17482 3765 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3701 17563 3765 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17563 3765 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 13613 3821 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 13613 3821 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 13695 3821 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 13695 3821 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 13777 3821 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 13777 3821 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 13859 3821 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 13859 3821 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 13941 3821 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 13941 3821 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14023 3821 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14023 3821 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14105 3821 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14105 3821 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14187 3821 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14187 3821 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14269 3821 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14269 3821 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14351 3821 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14351 3821 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14433 3821 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14433 3821 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14515 3821 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14515 3821 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14597 3821 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14597 3821 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14678 3821 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14678 3821 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14759 3821 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14759 3821 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14840 3821 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14840 3821 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14921 3821 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14921 3821 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15002 3821 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15002 3821 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15083 3821 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15083 3821 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15164 3821 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15164 3821 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15245 3821 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15245 3821 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15326 3821 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15326 3821 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15407 3821 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15407 3821 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15488 3821 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15488 3821 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15569 3821 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15569 3821 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15650 3821 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15650 3821 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15731 3821 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15731 3821 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15812 3821 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15812 3821 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15893 3821 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15893 3821 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15974 3821 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15974 3821 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 16055 3821 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16055 3821 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 16136 3821 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16136 3821 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 16217 3821 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16217 3821 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 16298 3821 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16298 3821 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 16379 3821 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16379 3821 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 16460 3821 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16460 3821 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3771 3560 3835 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3771 3560 3835 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3771 3646 3835 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3771 3646 3835 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3771 3732 3835 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3771 3732 3835 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3771 3818 3835 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3771 3818 3835 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3771 3904 3835 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3771 3904 3835 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3771 3990 3835 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3771 3990 3835 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3771 4076 3835 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3771 4076 3835 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3771 4162 3835 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3771 4162 3835 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3771 4248 3835 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3771 4248 3835 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3771 4334 3835 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3771 4334 3835 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3771 4420 3835 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3771 4420 3835 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3800 17163 3864 17227 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3800 17163 3864 17227 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3800 17250 3864 17314 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3800 17250 3864 17314 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3800 17338 3864 17402 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3800 17338 3864 17402 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 13613 3901 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 13613 3901 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 13695 3901 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 13695 3901 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 13777 3901 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 13777 3901 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 13859 3901 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 13859 3901 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 13941 3901 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 13941 3901 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14023 3901 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14023 3901 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14105 3901 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14105 3901 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14187 3901 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14187 3901 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14269 3901 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14269 3901 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14351 3901 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14351 3901 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14433 3901 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14433 3901 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14515 3901 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14515 3901 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14597 3901 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14597 3901 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14678 3901 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14678 3901 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14759 3901 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14759 3901 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14840 3901 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14840 3901 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14921 3901 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14921 3901 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15002 3901 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15002 3901 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15083 3901 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15083 3901 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15164 3901 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15164 3901 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15245 3901 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15245 3901 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15326 3901 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15326 3901 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15407 3901 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15407 3901 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15488 3901 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15488 3901 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15569 3901 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15569 3901 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15650 3901 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15650 3901 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15731 3901 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15731 3901 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15812 3901 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15812 3901 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15893 3901 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15893 3901 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15974 3901 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15974 3901 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 16055 3901 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16055 3901 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 16136 3901 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16136 3901 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 16217 3901 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16217 3901 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 16298 3901 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16298 3901 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 16379 3901 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16379 3901 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 16460 3901 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16460 3901 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3838 16590 3902 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 16590 3902 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3838 16682 3902 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 16682 3902 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3838 16774 3902 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 16774 3902 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3838 16867 3902 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 16867 3902 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3838 16960 3902 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 16960 3902 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3838 17053 3902 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 17053 3902 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3852 3560 3916 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3852 3560 3916 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3852 3646 3916 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3852 3646 3916 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3852 3732 3916 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3852 3732 3916 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3852 3818 3916 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3852 3818 3916 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3852 3904 3916 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3852 3904 3916 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3852 3990 3916 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3852 3990 3916 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3852 4076 3916 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3852 4076 3916 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3852 4162 3916 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3852 4162 3916 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3852 4248 3916 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3852 4248 3916 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3852 4334 3916 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3852 4334 3916 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3852 4420 3916 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3852 4420 3916 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 13613 3981 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 13613 3981 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 13695 3981 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 13695 3981 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 13777 3981 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 13777 3981 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 13859 3981 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 13859 3981 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 13941 3981 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 13941 3981 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14023 3981 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14023 3981 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14105 3981 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14105 3981 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14187 3981 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14187 3981 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14269 3981 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14269 3981 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14351 3981 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14351 3981 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14433 3981 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14433 3981 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14515 3981 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14515 3981 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14597 3981 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14597 3981 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14678 3981 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14678 3981 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14759 3981 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14759 3981 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14840 3981 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14840 3981 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14921 3981 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14921 3981 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15002 3981 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15002 3981 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15083 3981 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15083 3981 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15164 3981 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15164 3981 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15245 3981 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15245 3981 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15326 3981 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15326 3981 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15407 3981 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15407 3981 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15488 3981 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15488 3981 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15569 3981 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15569 3981 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15650 3981 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15650 3981 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15731 3981 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15731 3981 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15812 3981 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15812 3981 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15893 3981 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15893 3981 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15974 3981 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15974 3981 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 16055 3981 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16055 3981 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 16136 3981 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16136 3981 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 16217 3981 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16217 3981 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 16298 3981 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16298 3981 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 16379 3981 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16379 3981 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 16460 3981 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16460 3981 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3933 3560 3997 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3933 3560 3997 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3933 3646 3997 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3933 3646 3997 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3933 3732 3997 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3933 3732 3997 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3933 3818 3997 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3933 3818 3997 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3933 3904 3997 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3933 3904 3997 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3933 3990 3997 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3933 3990 3997 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3933 4076 3997 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3933 4076 3997 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3933 4162 3997 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3933 4162 3997 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3933 4248 3997 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3933 4248 3997 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3933 4334 3997 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3933 4334 3997 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3933 4420 3997 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3933 4420 3997 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3934 16590 3998 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 16590 3998 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3934 16682 3998 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 16682 3998 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3934 16774 3998 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 16774 3998 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3934 16867 3998 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 16867 3998 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3934 16960 3998 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 16960 3998 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3934 17053 3998 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 17053 3998 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3948 17163 4012 17227 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3948 17163 4012 17227 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3948 17250 4012 17314 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3948 17250 4012 17314 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3948 17338 4012 17402 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3948 17338 4012 17402 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 13613 4061 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 13613 4061 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 13695 4061 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 13695 4061 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 13777 4061 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 13777 4061 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 13859 4061 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 13859 4061 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 13941 4061 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 13941 4061 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14023 4061 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14023 4061 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14105 4061 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14105 4061 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14187 4061 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14187 4061 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14269 4061 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14269 4061 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14351 4061 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14351 4061 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14433 4061 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14433 4061 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14515 4061 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14515 4061 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14597 4061 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14597 4061 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14678 4061 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14678 4061 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14759 4061 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14759 4061 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14840 4061 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14840 4061 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14921 4061 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14921 4061 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15002 4061 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15002 4061 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15083 4061 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15083 4061 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15164 4061 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15164 4061 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15245 4061 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15245 4061 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15326 4061 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15326 4061 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15407 4061 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15407 4061 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15488 4061 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15488 4061 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15569 4061 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15569 4061 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15650 4061 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15650 4061 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15731 4061 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15731 4061 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15812 4061 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15812 4061 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15893 4061 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15893 4061 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15974 4061 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15974 4061 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 16055 4061 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16055 4061 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 16136 4061 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16136 4061 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 16217 4061 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16217 4061 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 16298 4061 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16298 4061 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 16379 4061 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16379 4061 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 16460 4061 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16460 4061 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 450 3560 514 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 450 3560 514 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 450 3646 514 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 450 3646 514 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 450 3732 514 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 450 3732 514 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 450 3818 514 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 450 3818 514 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 450 3904 514 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 450 3904 514 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 450 3990 514 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 450 3990 514 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 450 4076 514 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 450 4076 514 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 450 4162 514 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 450 4162 514 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 450 4248 514 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 450 4248 514 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 450 4334 514 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 450 4334 514 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 450 4420 514 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 450 4420 514 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 16559 527 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16559 527 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 16641 527 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16641 527 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 16723 527 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16723 527 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 16805 527 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16805 527 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 16887 527 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16887 527 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 16969 527 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16969 527 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17051 527 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17051 527 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17133 527 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17133 527 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17215 527 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17215 527 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17297 527 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17297 527 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17379 527 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17379 527 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17461 527 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17461 527 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17543 527 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17543 527 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17625 527 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17625 527 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17707 527 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17707 527 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17789 527 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17789 527 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17871 527 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17871 527 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17953 527 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17953 527 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 18035 527 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18035 527 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 18117 527 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18117 527 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 18199 527 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18199 527 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 18281 527 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18281 527 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 18363 527 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18363 527 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 18445 527 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18445 527 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 18527 527 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18527 527 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 13613 541 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 13613 541 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 13695 541 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 13695 541 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 13777 541 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 13777 541 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 13859 541 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 13859 541 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 13941 541 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 13941 541 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14023 541 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14023 541 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14105 541 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14105 541 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14187 541 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14187 541 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14269 541 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14269 541 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14351 541 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14351 541 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14433 541 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14433 541 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14515 541 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14515 541 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14597 541 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14597 541 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14678 541 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14678 541 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14759 541 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14759 541 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14840 541 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14840 541 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14921 541 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14921 541 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15002 541 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15002 541 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15083 541 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15083 541 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15164 541 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15164 541 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15245 541 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15245 541 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15326 541 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15326 541 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15407 541 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15407 541 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15488 541 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15488 541 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15569 541 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15569 541 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15650 541 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15650 541 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15731 541 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15731 541 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15812 541 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15812 541 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15893 541 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15893 541 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15974 541 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15974 541 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 16055 541 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16055 541 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 16136 541 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16136 541 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 16217 541 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16217 541 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 16298 541 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16298 541 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 16379 541 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16379 541 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 16460 541 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16460 541 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 531 3560 595 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 531 3560 595 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 531 3646 595 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 531 3646 595 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 531 3732 595 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 531 3732 595 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 531 3818 595 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 531 3818 595 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 531 3904 595 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 531 3904 595 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 531 3990 595 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 531 3990 595 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 531 4076 595 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 531 4076 595 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 531 4162 595 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 531 4162 595 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 531 4248 595 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 531 4248 595 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 531 4334 595 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 531 4334 595 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 531 4420 595 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 531 4420 595 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 16559 609 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16559 609 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 16641 609 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16641 609 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 16723 609 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16723 609 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 16805 609 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16805 609 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 16887 609 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16887 609 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 16969 609 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16969 609 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17051 609 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17051 609 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17133 609 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17133 609 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17215 609 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17215 609 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17297 609 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17297 609 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17379 609 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17379 609 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17461 609 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17461 609 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17543 609 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17543 609 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17625 609 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17625 609 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17707 609 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17707 609 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17789 609 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17789 609 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17871 609 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17871 609 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17953 609 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17953 609 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 18035 609 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18035 609 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 18117 609 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18117 609 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 18199 609 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18199 609 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 18281 609 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18281 609 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 18363 609 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18363 609 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 18445 609 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18445 609 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 18527 609 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18527 609 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 13613 621 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 13613 621 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 13695 621 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 13695 621 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 13777 621 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 13777 621 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 13859 621 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 13859 621 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 13941 621 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 13941 621 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14023 621 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14023 621 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14105 621 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14105 621 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14187 621 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14187 621 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14269 621 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14269 621 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14351 621 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14351 621 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14433 621 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14433 621 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14515 621 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14515 621 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14597 621 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14597 621 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14678 621 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14678 621 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14759 621 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14759 621 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14840 621 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14840 621 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14921 621 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14921 621 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15002 621 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15002 621 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15083 621 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15083 621 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15164 621 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15164 621 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15245 621 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15245 621 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15326 621 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15326 621 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15407 621 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15407 621 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15488 621 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15488 621 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15569 621 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15569 621 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15650 621 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15650 621 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15731 621 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15731 621 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15812 621 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15812 621 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15893 621 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15893 621 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15974 621 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15974 621 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 16055 621 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16055 621 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 16136 621 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16136 621 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 16217 621 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16217 621 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 16298 621 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16298 621 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 16379 621 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16379 621 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 16460 621 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16460 621 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4014 3560 4078 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4014 3560 4078 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4014 3646 4078 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4014 3646 4078 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4014 3732 4078 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4014 3732 4078 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4014 3818 4078 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4014 3818 4078 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4014 3904 4078 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4014 3904 4078 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4014 3990 4078 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4014 3990 4078 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4014 4076 4078 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4014 4076 4078 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4014 4162 4078 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4014 4162 4078 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4014 4248 4078 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4014 4248 4078 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4014 4334 4078 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4014 4334 4078 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4014 4420 4078 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4014 4420 4078 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4030 16590 4094 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 16590 4094 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4030 16682 4094 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 16682 4094 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4030 16774 4094 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 16774 4094 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4030 16867 4094 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 16867 4094 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4030 16960 4094 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 16960 4094 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4030 17053 4094 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 17053 4094 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 13613 4141 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 13613 4141 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 13695 4141 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 13695 4141 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 13777 4141 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 13777 4141 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 13859 4141 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 13859 4141 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 13941 4141 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 13941 4141 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14023 4141 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14023 4141 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14105 4141 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14105 4141 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14187 4141 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14187 4141 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14269 4141 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14269 4141 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14351 4141 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14351 4141 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14433 4141 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14433 4141 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14515 4141 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14515 4141 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14597 4141 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14597 4141 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14678 4141 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14678 4141 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14759 4141 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14759 4141 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14840 4141 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14840 4141 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14921 4141 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14921 4141 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15002 4141 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15002 4141 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15083 4141 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15083 4141 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15164 4141 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15164 4141 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15245 4141 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15245 4141 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15326 4141 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15326 4141 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15407 4141 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15407 4141 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15488 4141 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15488 4141 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15569 4141 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15569 4141 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15650 4141 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15650 4141 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15731 4141 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15731 4141 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15812 4141 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15812 4141 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15893 4141 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15893 4141 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15974 4141 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15974 4141 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 16055 4141 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16055 4141 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 16136 4141 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16136 4141 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 16217 4141 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16217 4141 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 16298 4141 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16298 4141 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 16379 4141 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16379 4141 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 16460 4141 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16460 4141 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4095 3560 4159 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4095 3560 4159 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4095 3646 4159 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4095 3646 4159 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4095 3732 4159 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4095 3732 4159 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4095 3818 4159 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4095 3818 4159 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4095 3904 4159 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4095 3904 4159 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4095 3990 4159 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4095 3990 4159 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4095 4076 4159 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4095 4076 4159 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4095 4162 4159 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4095 4162 4159 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4095 4248 4159 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4095 4248 4159 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4095 4334 4159 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4095 4334 4159 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4095 4420 4159 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4095 4420 4159 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4126 16590 4190 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 16590 4190 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4126 16682 4190 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 16682 4190 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4126 16774 4190 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 16774 4190 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4126 16867 4190 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 16867 4190 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4126 16960 4190 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 16960 4190 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4126 17053 4190 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 17053 4190 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 13613 4221 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 13613 4221 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 13695 4221 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 13695 4221 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 13777 4221 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 13777 4221 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 13859 4221 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 13859 4221 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 13941 4221 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 13941 4221 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14023 4221 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14023 4221 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14105 4221 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14105 4221 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14187 4221 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14187 4221 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14269 4221 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14269 4221 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14351 4221 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14351 4221 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14433 4221 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14433 4221 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14515 4221 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14515 4221 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14597 4221 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14597 4221 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14678 4221 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14678 4221 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14759 4221 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14759 4221 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14840 4221 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14840 4221 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14921 4221 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14921 4221 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15002 4221 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15002 4221 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15083 4221 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15083 4221 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15164 4221 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15164 4221 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15245 4221 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15245 4221 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15326 4221 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15326 4221 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15407 4221 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15407 4221 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15488 4221 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15488 4221 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15569 4221 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15569 4221 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15650 4221 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15650 4221 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15731 4221 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15731 4221 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15812 4221 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15812 4221 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15893 4221 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15893 4221 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15974 4221 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15974 4221 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 16055 4221 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16055 4221 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 16136 4221 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16136 4221 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 16217 4221 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16217 4221 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 16298 4221 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16298 4221 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 16379 4221 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16379 4221 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 16460 4221 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16460 4221 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4176 3560 4240 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4176 3560 4240 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4176 3646 4240 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4176 3646 4240 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4176 3732 4240 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4176 3732 4240 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4176 3818 4240 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4176 3818 4240 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4176 3904 4240 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4176 3904 4240 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4176 3990 4240 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4176 3990 4240 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4176 4076 4240 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4176 4076 4240 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4176 4162 4240 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4176 4162 4240 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4176 4248 4240 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4176 4248 4240 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4176 4334 4240 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4176 4334 4240 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4176 4420 4240 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4176 4420 4240 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4222 16590 4286 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 16590 4286 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4222 16682 4286 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 16682 4286 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4222 16774 4286 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 16774 4286 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4222 16867 4286 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 16867 4286 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4222 16960 4286 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 16960 4286 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4222 17053 4286 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 17053 4286 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 13613 4301 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 13613 4301 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 13695 4301 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 13695 4301 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 13777 4301 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 13777 4301 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 13859 4301 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 13859 4301 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 13941 4301 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 13941 4301 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14023 4301 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14023 4301 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14105 4301 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14105 4301 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14187 4301 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14187 4301 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14269 4301 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14269 4301 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14351 4301 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14351 4301 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14433 4301 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14433 4301 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14515 4301 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14515 4301 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14597 4301 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14597 4301 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14678 4301 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14678 4301 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14759 4301 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14759 4301 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14840 4301 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14840 4301 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14921 4301 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14921 4301 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15002 4301 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15002 4301 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15083 4301 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15083 4301 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15164 4301 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15164 4301 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15245 4301 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15245 4301 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15326 4301 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15326 4301 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15407 4301 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15407 4301 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15488 4301 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15488 4301 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15569 4301 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15569 4301 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15650 4301 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15650 4301 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15731 4301 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15731 4301 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15812 4301 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15812 4301 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15893 4301 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15893 4301 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15974 4301 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15974 4301 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 16055 4301 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16055 4301 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 16136 4301 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16136 4301 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 16217 4301 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16217 4301 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 16298 4301 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16298 4301 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 16379 4301 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16379 4301 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 16460 4301 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16460 4301 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4257 3560 4321 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4257 3560 4321 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4257 3646 4321 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4257 3646 4321 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4257 3732 4321 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4257 3732 4321 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4257 3818 4321 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4257 3818 4321 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4257 3904 4321 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4257 3904 4321 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4257 3990 4321 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4257 3990 4321 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4257 4076 4321 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4257 4076 4321 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4257 4162 4321 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4257 4162 4321 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4257 4248 4321 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4257 4248 4321 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4257 4334 4321 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4257 4334 4321 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4257 4420 4321 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4257 4420 4321 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 13613 4381 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 13613 4381 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 13695 4381 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 13695 4381 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 13777 4381 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 13777 4381 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 13859 4381 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 13859 4381 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 13941 4381 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 13941 4381 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14023 4381 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14023 4381 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14105 4381 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14105 4381 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14187 4381 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14187 4381 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14269 4381 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14269 4381 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14351 4381 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14351 4381 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14433 4381 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14433 4381 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14515 4381 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14515 4381 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14597 4381 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14597 4381 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14678 4381 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14678 4381 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14759 4381 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14759 4381 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14840 4381 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14840 4381 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14921 4381 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14921 4381 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15002 4381 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15002 4381 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15083 4381 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15083 4381 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15164 4381 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15164 4381 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15245 4381 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15245 4381 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15326 4381 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15326 4381 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15407 4381 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15407 4381 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15488 4381 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15488 4381 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15569 4381 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15569 4381 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15650 4381 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15650 4381 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15731 4381 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15731 4381 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15812 4381 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15812 4381 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15893 4381 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15893 4381 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15974 4381 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15974 4381 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 16055 4381 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16055 4381 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 16136 4381 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16136 4381 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 16217 4381 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16217 4381 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 16298 4381 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16298 4381 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 16379 4381 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16379 4381 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 16460 4381 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16460 4381 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4331 16572 4395 16636 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4331 16572 4395 16636 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4331 16682 4395 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4331 16682 4395 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4331 16792 4395 16856 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4331 16792 4395 16856 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4338 3560 4402 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4338 3560 4402 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4338 3646 4402 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4338 3646 4402 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4338 3732 4402 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4338 3732 4402 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4338 3818 4402 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4338 3818 4402 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4338 3904 4402 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4338 3904 4402 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4338 3990 4402 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4338 3990 4402 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4338 4076 4402 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4338 4076 4402 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4338 4162 4402 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4338 4162 4402 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4338 4248 4402 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4338 4248 4402 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4338 4334 4402 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4338 4334 4402 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4338 4420 4402 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4338 4420 4402 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 13613 4461 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 13613 4461 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 13695 4461 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 13695 4461 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 13777 4461 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 13777 4461 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 13859 4461 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 13859 4461 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 13941 4461 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 13941 4461 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14023 4461 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14023 4461 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14105 4461 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14105 4461 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14187 4461 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14187 4461 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14269 4461 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14269 4461 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14351 4461 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14351 4461 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14433 4461 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14433 4461 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14515 4461 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14515 4461 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14597 4461 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14597 4461 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14678 4461 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14678 4461 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14759 4461 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14759 4461 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14840 4461 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14840 4461 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14921 4461 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14921 4461 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15002 4461 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15002 4461 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15083 4461 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15083 4461 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15164 4461 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15164 4461 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15245 4461 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15245 4461 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15326 4461 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15326 4461 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15407 4461 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15407 4461 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15488 4461 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15488 4461 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15569 4461 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15569 4461 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15650 4461 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15650 4461 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15731 4461 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15731 4461 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15812 4461 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15812 4461 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15893 4461 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15893 4461 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15974 4461 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15974 4461 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 16055 4461 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16055 4461 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 16136 4461 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16136 4461 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 16217 4461 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16217 4461 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 16298 4461 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16298 4461 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 16379 4461 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16379 4461 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 16460 4461 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16460 4461 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4420 3560 4484 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4420 3560 4484 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4420 3646 4484 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4420 3646 4484 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4420 3732 4484 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4420 3732 4484 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4420 3818 4484 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4420 3818 4484 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4420 3904 4484 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4420 3904 4484 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4420 3990 4484 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4420 3990 4484 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4420 4076 4484 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4420 4076 4484 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4420 4162 4484 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4420 4162 4484 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4420 4248 4484 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4420 4248 4484 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4420 4334 4484 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4420 4334 4484 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4420 4420 4484 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4420 4420 4484 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 13613 4541 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 13613 4541 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 13695 4541 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 13695 4541 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 13777 4541 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 13777 4541 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 13859 4541 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 13859 4541 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 13941 4541 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 13941 4541 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14023 4541 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14023 4541 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14105 4541 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14105 4541 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14187 4541 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14187 4541 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14269 4541 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14269 4541 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14351 4541 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14351 4541 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14433 4541 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14433 4541 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14515 4541 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14515 4541 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14597 4541 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14597 4541 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14678 4541 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14678 4541 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14759 4541 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14759 4541 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14840 4541 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14840 4541 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14921 4541 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14921 4541 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15002 4541 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15002 4541 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15083 4541 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15083 4541 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15164 4541 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15164 4541 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15245 4541 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15245 4541 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15326 4541 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15326 4541 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15407 4541 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15407 4541 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15488 4541 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15488 4541 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15569 4541 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15569 4541 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15650 4541 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15650 4541 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15731 4541 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15731 4541 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15812 4541 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15812 4541 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15893 4541 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15893 4541 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15974 4541 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15974 4541 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 16055 4541 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16055 4541 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 16136 4541 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16136 4541 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 16217 4541 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16217 4541 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 16298 4541 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16298 4541 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 16379 4541 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16379 4541 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 16460 4541 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16460 4541 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4489 16572 4553 16636 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 16572 4553 16636 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4489 16682 4553 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 16682 4553 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4489 16792 4553 16856 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 16792 4553 16856 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4502 3560 4566 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4502 3560 4566 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4502 3646 4566 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4502 3646 4566 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4502 3732 4566 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4502 3732 4566 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4502 3818 4566 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4502 3818 4566 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4502 3904 4566 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4502 3904 4566 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4502 3990 4566 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4502 3990 4566 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4502 4076 4566 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4502 4076 4566 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4502 4162 4566 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4502 4162 4566 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4502 4248 4566 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4502 4248 4566 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4502 4334 4566 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4502 4334 4566 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4502 4420 4566 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4502 4420 4566 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 13613 4621 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 13613 4621 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 13695 4621 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 13695 4621 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 13777 4621 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 13777 4621 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 13859 4621 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 13859 4621 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 13941 4621 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 13941 4621 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14023 4621 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14023 4621 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14105 4621 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14105 4621 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14187 4621 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14187 4621 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14269 4621 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14269 4621 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14351 4621 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14351 4621 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14433 4621 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14433 4621 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14515 4621 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14515 4621 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14597 4621 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14597 4621 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14678 4621 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14678 4621 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14759 4621 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14759 4621 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14840 4621 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14840 4621 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14921 4621 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14921 4621 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15002 4621 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15002 4621 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15083 4621 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15083 4621 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15164 4621 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15164 4621 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15245 4621 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15245 4621 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15326 4621 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15326 4621 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15407 4621 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15407 4621 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15488 4621 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15488 4621 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15569 4621 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15569 4621 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15650 4621 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15650 4621 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15731 4621 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15731 4621 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15812 4621 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15812 4621 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15893 4621 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15893 4621 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15974 4621 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15974 4621 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 16055 4621 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16055 4621 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 16136 4621 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16136 4621 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 16217 4621 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16217 4621 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 16298 4621 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16298 4621 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 16379 4621 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16379 4621 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 16460 4621 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16460 4621 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4584 3560 4648 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4584 3560 4648 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4584 3646 4648 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4584 3646 4648 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4584 3732 4648 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4584 3732 4648 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4584 3818 4648 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4584 3818 4648 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4584 3904 4648 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4584 3904 4648 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4584 3990 4648 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4584 3990 4648 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4584 4076 4648 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4584 4076 4648 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4584 4162 4648 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4584 4162 4648 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4584 4248 4648 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4584 4248 4648 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4584 4334 4648 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4584 4334 4648 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4584 4420 4648 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4584 4420 4648 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 13613 4701 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 13613 4701 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 13695 4701 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 13695 4701 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 13777 4701 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 13777 4701 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 13859 4701 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 13859 4701 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 13941 4701 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 13941 4701 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14023 4701 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14023 4701 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14105 4701 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14105 4701 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14187 4701 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14187 4701 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14269 4701 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14269 4701 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14351 4701 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14351 4701 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14433 4701 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14433 4701 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14515 4701 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14515 4701 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14597 4701 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14597 4701 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14678 4701 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14678 4701 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14759 4701 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14759 4701 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14840 4701 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14840 4701 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14921 4701 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14921 4701 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15002 4701 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15002 4701 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15083 4701 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15083 4701 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15164 4701 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15164 4701 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15245 4701 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15245 4701 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15326 4701 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15326 4701 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15407 4701 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15407 4701 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15488 4701 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15488 4701 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15569 4701 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15569 4701 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15650 4701 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15650 4701 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15731 4701 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15731 4701 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15812 4701 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15812 4701 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15893 4701 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15893 4701 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15974 4701 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15974 4701 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 16055 4701 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16055 4701 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 16136 4701 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16136 4701 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 16217 4701 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16217 4701 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 16298 4701 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16298 4701 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 16379 4701 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16379 4701 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 16460 4701 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16460 4701 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4666 3560 4730 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4666 3560 4730 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4666 3646 4730 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4666 3646 4730 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4666 3732 4730 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4666 3732 4730 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4666 3818 4730 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4666 3818 4730 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4666 3904 4730 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4666 3904 4730 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4666 3990 4730 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4666 3990 4730 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4666 4076 4730 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4666 4076 4730 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4666 4162 4730 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4666 4162 4730 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4666 4248 4730 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4666 4248 4730 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4666 4334 4730 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4666 4334 4730 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4666 4420 4730 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4666 4420 4730 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 13613 4781 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 13613 4781 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 13695 4781 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 13695 4781 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 13777 4781 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 13777 4781 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 13859 4781 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 13859 4781 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 13941 4781 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 13941 4781 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14023 4781 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14023 4781 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14105 4781 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14105 4781 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14187 4781 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14187 4781 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14269 4781 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14269 4781 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14351 4781 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14351 4781 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14433 4781 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14433 4781 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14515 4781 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14515 4781 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14597 4781 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14597 4781 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14678 4781 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14678 4781 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14759 4781 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14759 4781 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14840 4781 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14840 4781 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14921 4781 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14921 4781 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15002 4781 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15002 4781 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15083 4781 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15083 4781 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15164 4781 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15164 4781 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15245 4781 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15245 4781 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15326 4781 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15326 4781 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15407 4781 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15407 4781 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15488 4781 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15488 4781 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15569 4781 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15569 4781 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15650 4781 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15650 4781 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15731 4781 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15731 4781 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15812 4781 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15812 4781 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15893 4781 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15893 4781 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15974 4781 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15974 4781 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 16055 4781 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16055 4781 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 16136 4781 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16136 4781 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 16217 4781 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16217 4781 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 16298 4781 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16298 4781 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 16379 4781 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16379 4781 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 16460 4781 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16460 4781 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4748 3560 4812 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4748 3560 4812 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4748 3646 4812 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4748 3646 4812 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4748 3732 4812 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4748 3732 4812 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4748 3818 4812 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4748 3818 4812 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4748 3904 4812 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4748 3904 4812 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4748 3990 4812 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4748 3990 4812 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4748 4076 4812 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4748 4076 4812 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4748 4162 4812 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4748 4162 4812 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4748 4248 4812 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4748 4248 4812 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4748 4334 4812 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4748 4334 4812 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4748 4420 4812 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4748 4420 4812 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 13613 4861 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 13613 4861 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 13695 4861 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 13695 4861 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 13777 4861 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 13777 4861 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 13859 4861 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 13859 4861 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 13941 4861 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 13941 4861 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14023 4861 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14023 4861 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14105 4861 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14105 4861 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14187 4861 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14187 4861 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14269 4861 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14269 4861 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14351 4861 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14351 4861 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14433 4861 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14433 4861 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14515 4861 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14515 4861 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14597 4861 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14597 4861 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14678 4861 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14678 4861 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14759 4861 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14759 4861 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14840 4861 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14840 4861 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14921 4861 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14921 4861 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15002 4861 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15002 4861 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15083 4861 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15083 4861 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15164 4861 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15164 4861 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15245 4861 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15245 4861 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15326 4861 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15326 4861 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15407 4861 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15407 4861 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15488 4861 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15488 4861 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15569 4861 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15569 4861 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15650 4861 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15650 4861 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15731 4861 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15731 4861 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15812 4861 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15812 4861 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15893 4861 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15893 4861 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15974 4861 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15974 4861 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 16055 4861 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16055 4861 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 16136 4861 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16136 4861 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 16217 4861 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16217 4861 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 16298 4861 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16298 4861 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 16379 4861 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16379 4861 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 16460 4861 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16460 4861 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4830 3560 4894 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4830 3560 4894 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4830 3646 4894 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4830 3646 4894 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4830 3732 4894 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4830 3732 4894 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4830 3818 4894 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4830 3818 4894 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4830 3904 4894 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4830 3904 4894 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4830 3990 4894 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4830 3990 4894 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4830 4076 4894 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4830 4076 4894 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4830 4162 4894 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4830 4162 4894 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4830 4248 4894 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4830 4248 4894 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4830 4334 4894 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4830 4334 4894 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4830 4420 4894 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4830 4420 4894 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 612 3560 676 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 612 3560 676 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 612 3646 676 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 612 3646 676 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 612 3732 676 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 612 3732 676 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 612 3818 676 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 612 3818 676 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 612 3904 676 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 612 3904 676 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 612 3990 676 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 612 3990 676 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 612 4076 676 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 612 4076 676 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 612 4162 676 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 612 4162 676 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 612 4248 676 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 612 4248 676 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 612 4334 676 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 612 4334 676 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 612 4420 676 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 612 4420 676 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 16559 691 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16559 691 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 16641 691 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16641 691 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 16723 691 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16723 691 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 16805 691 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16805 691 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 16887 691 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16887 691 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 16969 691 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16969 691 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17051 691 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17051 691 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17133 691 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17133 691 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17215 691 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17215 691 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17297 691 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17297 691 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17379 691 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17379 691 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17461 691 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17461 691 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17543 691 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17543 691 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17625 691 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17625 691 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17707 691 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17707 691 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17789 691 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17789 691 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17871 691 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17871 691 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17953 691 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17953 691 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 18035 691 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18035 691 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 18117 691 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18117 691 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 18199 691 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18199 691 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 18281 691 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18281 691 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 18363 691 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18363 691 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 18445 691 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18445 691 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 18527 691 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18527 691 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 13613 701 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 13613 701 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 13695 701 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 13695 701 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 13777 701 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 13777 701 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 13859 701 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 13859 701 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 13941 701 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 13941 701 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14023 701 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14023 701 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14105 701 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14105 701 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14187 701 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14187 701 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14269 701 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14269 701 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14351 701 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14351 701 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14433 701 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14433 701 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14515 701 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14515 701 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14597 701 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14597 701 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14678 701 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14678 701 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14759 701 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14759 701 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14840 701 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14840 701 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14921 701 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14921 701 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15002 701 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15002 701 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15083 701 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15083 701 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15164 701 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15164 701 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15245 701 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15245 701 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15326 701 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15326 701 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15407 701 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15407 701 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15488 701 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15488 701 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15569 701 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15569 701 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15650 701 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15650 701 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15731 701 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15731 701 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15812 701 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15812 701 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15893 701 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15893 701 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15974 701 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15974 701 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 16055 701 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16055 701 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 16136 701 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16136 701 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 16217 701 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16217 701 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 16298 701 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16298 701 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 16379 701 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16379 701 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 16460 701 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16460 701 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 693 3560 757 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 693 3560 757 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 693 3646 757 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 693 3646 757 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 693 3732 757 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 693 3732 757 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 693 3818 757 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 693 3818 757 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 693 3904 757 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 693 3904 757 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 693 3990 757 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 693 3990 757 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 693 4076 757 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 693 4076 757 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 693 4162 757 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 693 4162 757 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 693 4248 757 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 693 4248 757 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 693 4334 757 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 693 4334 757 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 693 4420 757 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 693 4420 757 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 16559 773 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16559 773 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 16641 773 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16641 773 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 16723 773 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16723 773 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 16805 773 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16805 773 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 16887 773 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16887 773 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 16969 773 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16969 773 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17051 773 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17051 773 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17133 773 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17133 773 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17215 773 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17215 773 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17297 773 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17297 773 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17379 773 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17379 773 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17461 773 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17461 773 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17543 773 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17543 773 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17625 773 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17625 773 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17707 773 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17707 773 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17789 773 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17789 773 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17871 773 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17871 773 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17953 773 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17953 773 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 18035 773 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18035 773 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 18117 773 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18117 773 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 18199 773 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18199 773 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 18281 773 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18281 773 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 18363 773 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18363 773 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 18445 773 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18445 773 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 18527 773 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18527 773 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 13613 781 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 13613 781 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 13695 781 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 13695 781 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 13777 781 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 13777 781 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 13859 781 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 13859 781 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 13941 781 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 13941 781 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14023 781 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14023 781 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14105 781 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14105 781 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14187 781 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14187 781 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14269 781 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14269 781 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14351 781 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14351 781 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14433 781 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14433 781 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14515 781 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14515 781 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14597 781 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14597 781 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14678 781 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14678 781 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14759 781 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14759 781 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14840 781 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14840 781 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14921 781 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14921 781 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15002 781 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15002 781 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15083 781 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15083 781 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15164 781 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15164 781 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15245 781 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15245 781 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15326 781 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15326 781 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15407 781 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15407 781 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15488 781 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15488 781 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15569 781 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15569 781 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15650 781 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15650 781 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15731 781 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15731 781 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15812 781 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15812 781 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15893 781 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15893 781 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15974 781 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15974 781 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 16055 781 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16055 781 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 16136 781 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16136 781 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 16217 781 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16217 781 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 16298 781 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16298 781 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 16379 781 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16379 781 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 16460 781 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16460 781 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 774 3560 838 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 774 3560 838 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 774 3646 838 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 774 3646 838 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 774 3732 838 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 774 3732 838 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 774 3818 838 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 774 3818 838 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 774 3904 838 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 774 3904 838 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 774 3990 838 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 774 3990 838 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 774 4076 838 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 774 4076 838 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 774 4162 838 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 774 4162 838 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 774 4248 838 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 774 4248 838 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 774 4334 838 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 774 4334 838 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 774 4420 838 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 774 4420 838 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 16559 855 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16559 855 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 16641 855 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16641 855 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 16723 855 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16723 855 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 16805 855 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16805 855 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 16887 855 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16887 855 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 16969 855 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16969 855 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17051 855 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17051 855 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17133 855 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17133 855 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17215 855 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17215 855 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17297 855 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17297 855 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17379 855 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17379 855 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17461 855 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17461 855 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17543 855 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17543 855 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17625 855 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17625 855 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17707 855 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17707 855 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17789 855 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17789 855 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17871 855 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17871 855 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17953 855 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17953 855 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 18035 855 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18035 855 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 18117 855 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18117 855 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 18199 855 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18199 855 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 18281 855 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18281 855 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 18363 855 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18363 855 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 18445 855 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18445 855 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 18527 855 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18527 855 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 13613 861 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 13613 861 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 13695 861 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 13695 861 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 13777 861 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 13777 861 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 13859 861 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 13859 861 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 13941 861 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 13941 861 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14023 861 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14023 861 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14105 861 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14105 861 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14187 861 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14187 861 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14269 861 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14269 861 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14351 861 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14351 861 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14433 861 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14433 861 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14515 861 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14515 861 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14597 861 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14597 861 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14678 861 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14678 861 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14759 861 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14759 861 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14840 861 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14840 861 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14921 861 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14921 861 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15002 861 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15002 861 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15083 861 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15083 861 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15164 861 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15164 861 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15245 861 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15245 861 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15326 861 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15326 861 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15407 861 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15407 861 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15488 861 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15488 861 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15569 861 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15569 861 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15650 861 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15650 861 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15731 861 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15731 861 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15812 861 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15812 861 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15893 861 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15893 861 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15974 861 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15974 861 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 16055 861 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16055 861 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 16136 861 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16136 861 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 16217 861 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16217 861 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 16298 861 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16298 861 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 16379 861 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16379 861 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 16460 861 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16460 861 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 855 3560 919 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 855 3560 919 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 855 3646 919 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 855 3646 919 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 855 3732 919 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 855 3732 919 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 855 3818 919 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 855 3818 919 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 855 3904 919 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 855 3904 919 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 855 3990 919 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 855 3990 919 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 855 4076 919 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 855 4076 919 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 855 4162 919 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 855 4162 919 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 855 4248 919 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 855 4248 919 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 855 4334 919 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 855 4334 919 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 855 4420 919 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 855 4420 919 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 16559 937 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16559 937 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 16641 937 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16641 937 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 16723 937 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16723 937 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 16805 937 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16805 937 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 16887 937 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16887 937 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 16969 937 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16969 937 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17051 937 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17051 937 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17133 937 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17133 937 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17215 937 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17215 937 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17297 937 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17297 937 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17379 937 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17379 937 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17461 937 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17461 937 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17543 937 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17543 937 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17625 937 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17625 937 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17707 937 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17707 937 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17789 937 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17789 937 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17871 937 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17871 937 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17953 937 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17953 937 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 18035 937 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18035 937 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 18117 937 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18117 937 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 18199 937 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18199 937 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 18281 937 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18281 937 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 18363 937 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18363 937 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 18445 937 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18445 937 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 18527 937 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18527 937 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 13613 941 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 13613 941 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 13695 941 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 13695 941 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 13777 941 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 13777 941 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 13859 941 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 13859 941 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 13941 941 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 13941 941 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14023 941 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14023 941 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14105 941 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14105 941 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14187 941 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14187 941 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14269 941 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14269 941 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14351 941 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14351 941 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14433 941 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14433 941 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14515 941 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14515 941 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14597 941 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14597 941 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14678 941 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14678 941 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14759 941 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14759 941 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14840 941 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14840 941 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14921 941 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14921 941 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15002 941 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15002 941 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15083 941 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15083 941 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15164 941 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15164 941 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15245 941 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15245 941 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15326 941 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15326 941 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15407 941 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15407 941 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15488 941 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15488 941 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15569 941 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15569 941 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15650 941 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15650 941 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15731 941 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15731 941 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15812 941 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15812 941 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15893 941 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15893 941 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15974 941 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15974 941 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 16055 941 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16055 941 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 16136 941 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16136 941 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 16217 941 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16217 941 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 16298 941 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16298 941 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 16379 941 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16379 941 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 16460 941 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16460 941 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 936 3560 1000 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 936 3560 1000 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 936 3646 1000 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 936 3646 1000 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 936 3732 1000 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 936 3732 1000 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 936 3818 1000 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 936 3818 1000 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 936 3904 1000 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 936 3904 1000 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 936 3990 1000 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 936 3990 1000 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 936 4076 1000 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 936 4076 1000 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 936 4162 1000 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 936 4162 1000 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 936 4248 1000 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 936 4248 1000 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 936 4334 1000 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 936 4334 1000 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 936 4420 1000 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 936 4420 1000 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 16559 1019 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16559 1019 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 16641 1019 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16641 1019 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 16723 1019 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16723 1019 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 16805 1019 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16805 1019 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 16887 1019 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16887 1019 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 16969 1019 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16969 1019 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17051 1019 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17051 1019 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17133 1019 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17133 1019 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17215 1019 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17215 1019 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17297 1019 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17297 1019 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17379 1019 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17379 1019 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17461 1019 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17461 1019 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17543 1019 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17543 1019 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17625 1019 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17625 1019 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17707 1019 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17707 1019 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17789 1019 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17789 1019 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17871 1019 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17871 1019 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17953 1019 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17953 1019 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 18035 1019 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18035 1019 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 18117 1019 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18117 1019 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 18199 1019 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18199 1019 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 18281 1019 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18281 1019 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 18363 1019 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18363 1019 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 18445 1019 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18445 1019 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 18527 1019 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18527 1019 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 13613 1021 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 13613 1021 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 13695 1021 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 13695 1021 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 13777 1021 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 13777 1021 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 13859 1021 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 13859 1021 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 13941 1021 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 13941 1021 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14023 1021 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14023 1021 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14105 1021 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14105 1021 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14187 1021 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14187 1021 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14269 1021 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14269 1021 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14351 1021 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14351 1021 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14433 1021 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14433 1021 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14515 1021 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14515 1021 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14597 1021 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14597 1021 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14678 1021 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14678 1021 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14759 1021 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14759 1021 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14840 1021 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14840 1021 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14921 1021 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14921 1021 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15002 1021 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15002 1021 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15083 1021 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15083 1021 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15164 1021 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15164 1021 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15245 1021 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15245 1021 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15326 1021 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15326 1021 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15407 1021 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15407 1021 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15488 1021 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15488 1021 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15569 1021 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15569 1021 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15650 1021 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15650 1021 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15731 1021 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15731 1021 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15812 1021 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15812 1021 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15893 1021 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15893 1021 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15974 1021 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15974 1021 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 16055 1021 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16055 1021 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 16136 1021 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16136 1021 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 16217 1021 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16217 1021 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 16298 1021 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16298 1021 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 16379 1021 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16379 1021 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 16460 1021 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16460 1021 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1017 3560 1081 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1017 3560 1081 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1017 3646 1081 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1017 3646 1081 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1017 3732 1081 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1017 3732 1081 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1017 3818 1081 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1017 3818 1081 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1017 3904 1081 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1017 3904 1081 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1017 3990 1081 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1017 3990 1081 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1017 4076 1081 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1017 4076 1081 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1017 4162 1081 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1017 4162 1081 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1017 4248 1081 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1017 4248 1081 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1017 4334 1081 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1017 4334 1081 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1017 4420 1081 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1017 4420 1081 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 13613 1101 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 13613 1101 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 13695 1101 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 13695 1101 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 13777 1101 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 13777 1101 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 13859 1101 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 13859 1101 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 13941 1101 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 13941 1101 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14023 1101 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14023 1101 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14105 1101 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14105 1101 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14187 1101 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14187 1101 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14269 1101 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14269 1101 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14351 1101 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14351 1101 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14433 1101 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14433 1101 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14515 1101 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14515 1101 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14597 1101 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14597 1101 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14678 1101 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14678 1101 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14759 1101 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14759 1101 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14840 1101 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14840 1101 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14921 1101 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14921 1101 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15002 1101 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15002 1101 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15083 1101 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15083 1101 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15164 1101 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15164 1101 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15245 1101 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15245 1101 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15326 1101 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15326 1101 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15407 1101 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15407 1101 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15488 1101 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15488 1101 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15569 1101 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15569 1101 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15650 1101 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15650 1101 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15731 1101 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15731 1101 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15812 1101 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15812 1101 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15893 1101 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15893 1101 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15974 1101 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15974 1101 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16055 1101 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16055 1101 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16136 1101 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16136 1101 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16217 1101 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16217 1101 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16298 1101 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16298 1101 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16379 1101 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16379 1101 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16460 1101 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16460 1101 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16559 1101 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16559 1101 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16641 1101 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16641 1101 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16723 1101 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16723 1101 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16805 1101 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16805 1101 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16887 1101 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16887 1101 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16969 1101 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16969 1101 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17051 1101 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17051 1101 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17133 1101 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17133 1101 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17215 1101 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17215 1101 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17297 1101 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17297 1101 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17379 1101 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17379 1101 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17461 1101 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17461 1101 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17543 1101 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17543 1101 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17625 1101 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17625 1101 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17707 1101 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17707 1101 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17789 1101 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17789 1101 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17871 1101 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17871 1101 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17953 1101 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17953 1101 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 18035 1101 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18035 1101 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 18117 1101 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18117 1101 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 18199 1101 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18199 1101 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 18281 1101 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18281 1101 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 18363 1101 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18363 1101 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 18445 1101 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18445 1101 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 18527 1101 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18527 1101 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1098 3560 1162 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1098 3560 1162 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1098 3646 1162 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1098 3646 1162 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1098 3732 1162 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1098 3732 1162 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1098 3818 1162 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1098 3818 1162 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1098 3904 1162 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1098 3904 1162 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1098 3990 1162 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1098 3990 1162 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1098 4076 1162 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1098 4076 1162 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1098 4162 1162 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1098 4162 1162 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1098 4248 1162 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1098 4248 1162 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1098 4334 1162 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1098 4334 1162 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1098 4420 1162 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1098 4420 1162 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 13613 1181 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 13613 1181 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 13695 1181 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 13695 1181 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 13777 1181 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 13777 1181 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 13859 1181 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 13859 1181 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 13941 1181 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 13941 1181 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14023 1181 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14023 1181 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14105 1181 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14105 1181 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14187 1181 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14187 1181 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14269 1181 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14269 1181 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14351 1181 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14351 1181 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14433 1181 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14433 1181 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14515 1181 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14515 1181 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14597 1181 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14597 1181 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14678 1181 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14678 1181 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14759 1181 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14759 1181 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14840 1181 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14840 1181 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14921 1181 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14921 1181 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15002 1181 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15002 1181 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15083 1181 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15083 1181 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15164 1181 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15164 1181 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15245 1181 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15245 1181 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15326 1181 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15326 1181 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15407 1181 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15407 1181 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15488 1181 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15488 1181 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15569 1181 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15569 1181 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15650 1181 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15650 1181 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15731 1181 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15731 1181 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15812 1181 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15812 1181 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15893 1181 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15893 1181 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15974 1181 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15974 1181 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 16055 1181 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16055 1181 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 16136 1181 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16136 1181 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 16217 1181 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16217 1181 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 16298 1181 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16298 1181 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 16379 1181 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16379 1181 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 16460 1181 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16460 1181 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 16559 1183 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16559 1183 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 16641 1183 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16641 1183 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 16723 1183 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16723 1183 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 16805 1183 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16805 1183 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 16887 1183 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16887 1183 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 16969 1183 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16969 1183 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17051 1183 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17051 1183 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17133 1183 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17133 1183 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17215 1183 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17215 1183 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17297 1183 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17297 1183 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17379 1183 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17379 1183 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17461 1183 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17461 1183 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17543 1183 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17543 1183 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17625 1183 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17625 1183 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17707 1183 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17707 1183 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17789 1183 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17789 1183 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17871 1183 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17871 1183 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17953 1183 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17953 1183 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 18035 1183 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18035 1183 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 18117 1183 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18117 1183 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 18199 1183 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18199 1183 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 18281 1183 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18281 1183 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 18363 1183 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18363 1183 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 18445 1183 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18445 1183 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 18527 1183 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18527 1183 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1179 3560 1243 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1179 3560 1243 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1179 3646 1243 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1179 3646 1243 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1179 3732 1243 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1179 3732 1243 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1179 3818 1243 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1179 3818 1243 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1179 3904 1243 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1179 3904 1243 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1179 3990 1243 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1179 3990 1243 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1179 4076 1243 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1179 4076 1243 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1179 4162 1243 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1179 4162 1243 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1179 4248 1243 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1179 4248 1243 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1179 4334 1243 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1179 4334 1243 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1179 4420 1243 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1179 4420 1243 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 13613 1261 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 13613 1261 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 13695 1261 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 13695 1261 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 13777 1261 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 13777 1261 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 13859 1261 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 13859 1261 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 13941 1261 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 13941 1261 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14023 1261 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14023 1261 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14105 1261 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14105 1261 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14187 1261 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14187 1261 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14269 1261 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14269 1261 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14351 1261 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14351 1261 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14433 1261 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14433 1261 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14515 1261 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14515 1261 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14597 1261 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14597 1261 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14678 1261 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14678 1261 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14759 1261 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14759 1261 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14840 1261 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14840 1261 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14921 1261 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14921 1261 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15002 1261 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15002 1261 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15083 1261 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15083 1261 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15164 1261 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15164 1261 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15245 1261 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15245 1261 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15326 1261 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15326 1261 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15407 1261 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15407 1261 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15488 1261 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15488 1261 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15569 1261 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15569 1261 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15650 1261 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15650 1261 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15731 1261 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15731 1261 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15812 1261 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15812 1261 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15893 1261 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15893 1261 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15974 1261 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15974 1261 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 16055 1261 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16055 1261 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 16136 1261 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16136 1261 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 16217 1261 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16217 1261 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 16298 1261 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16298 1261 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 16379 1261 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16379 1261 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 16460 1261 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16460 1261 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10157 3560 10221 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10157 3560 10221 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10157 3646 10221 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10157 3646 10221 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10157 3732 10221 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10157 3732 10221 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10157 3818 10221 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10157 3818 10221 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10157 3904 10221 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10157 3904 10221 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10157 3990 10221 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10157 3990 10221 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10157 4076 10221 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10157 4076 10221 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10157 4162 10221 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10157 4162 10221 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10157 4248 10221 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10157 4248 10221 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10157 4334 10221 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10157 4334 10221 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10157 4420 10221 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10157 4420 10221 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 13613 10254 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 13613 10254 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 13695 10254 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 13695 10254 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 13777 10254 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 13777 10254 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 13859 10254 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 13859 10254 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 13941 10254 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 13941 10254 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 14023 10254 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 14023 10254 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 14105 10254 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 14105 10254 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 14187 10254 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 14187 10254 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 14269 10254 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 14269 10254 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 14351 10254 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 14351 10254 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 14433 10254 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 14433 10254 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 14515 10254 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 14515 10254 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 14597 10254 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 14597 10254 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 14678 10254 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 14678 10254 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 14759 10254 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 14759 10254 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 14840 10254 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 14840 10254 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 14921 10254 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 14921 10254 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 15002 10254 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 15002 10254 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 15083 10254 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 15083 10254 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 15164 10254 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 15164 10254 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 15245 10254 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 15245 10254 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 15326 10254 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 15326 10254 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 15407 10254 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 15407 10254 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 15488 10254 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 15488 10254 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 15569 10254 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 15569 10254 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 15650 10254 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 15650 10254 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 15731 10254 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 15731 10254 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 15812 10254 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 15812 10254 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 15893 10254 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 15893 10254 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 15974 10254 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 15974 10254 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 16055 10254 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 16055 10254 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 16136 10254 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 16136 10254 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 16217 10254 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 16217 10254 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 16298 10254 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 16298 10254 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 16379 10254 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 16379 10254 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10190 16460 10254 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10190 16460 10254 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10238 3560 10302 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10238 3560 10302 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10238 3646 10302 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10238 3646 10302 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10238 3732 10302 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10238 3732 10302 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10238 3818 10302 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10238 3818 10302 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10238 3904 10302 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10238 3904 10302 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10238 3990 10302 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10238 3990 10302 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10238 4076 10302 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10238 4076 10302 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10238 4162 10302 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10238 4162 10302 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10238 4248 10302 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10238 4248 10302 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10238 4334 10302 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10238 4334 10302 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10238 4420 10302 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10238 4420 10302 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 13613 10334 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 13613 10334 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 13695 10334 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 13695 10334 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 13777 10334 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 13777 10334 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 13859 10334 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 13859 10334 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 13941 10334 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 13941 10334 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 14023 10334 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 14023 10334 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 14105 10334 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 14105 10334 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 14187 10334 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 14187 10334 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 14269 10334 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 14269 10334 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 14351 10334 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 14351 10334 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 14433 10334 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 14433 10334 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 14515 10334 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 14515 10334 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 14597 10334 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 14597 10334 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 14678 10334 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 14678 10334 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 14759 10334 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 14759 10334 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 14840 10334 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 14840 10334 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 14921 10334 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 14921 10334 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 15002 10334 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 15002 10334 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 15083 10334 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 15083 10334 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 15164 10334 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 15164 10334 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 15245 10334 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 15245 10334 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 15326 10334 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 15326 10334 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 15407 10334 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 15407 10334 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 15488 10334 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 15488 10334 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 15569 10334 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 15569 10334 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 15650 10334 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 15650 10334 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 15731 10334 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 15731 10334 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 15812 10334 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 15812 10334 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 15893 10334 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 15893 10334 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 15974 10334 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 15974 10334 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 16055 10334 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 16055 10334 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 16136 10334 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 16136 10334 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 16217 10334 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 16217 10334 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 16298 10334 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 16298 10334 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 16379 10334 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 16379 10334 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10270 16460 10334 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10270 16460 10334 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10319 3560 10383 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10319 3560 10383 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10319 3646 10383 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10319 3646 10383 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10319 3732 10383 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10319 3732 10383 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10319 3818 10383 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10319 3818 10383 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10319 3904 10383 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10319 3904 10383 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10319 3990 10383 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10319 3990 10383 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10319 4076 10383 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10319 4076 10383 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10319 4162 10383 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10319 4162 10383 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10319 4248 10383 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10319 4248 10383 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10319 4334 10383 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10319 4334 10383 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10319 4420 10383 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10319 4420 10383 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 13613 10414 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 13613 10414 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 13695 10414 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 13695 10414 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 13777 10414 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 13777 10414 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 13859 10414 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 13859 10414 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 13941 10414 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 13941 10414 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 14023 10414 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 14023 10414 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 14105 10414 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 14105 10414 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 14187 10414 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 14187 10414 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 14269 10414 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 14269 10414 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 14351 10414 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 14351 10414 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 14433 10414 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 14433 10414 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 14515 10414 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 14515 10414 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 14597 10414 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 14597 10414 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 14678 10414 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 14678 10414 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 14759 10414 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 14759 10414 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 14840 10414 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 14840 10414 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 14921 10414 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 14921 10414 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 15002 10414 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 15002 10414 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 15083 10414 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 15083 10414 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 15164 10414 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 15164 10414 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 15245 10414 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 15245 10414 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 15326 10414 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 15326 10414 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 15407 10414 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 15407 10414 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 15488 10414 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 15488 10414 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 15569 10414 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 15569 10414 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 15650 10414 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 15650 10414 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 15731 10414 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 15731 10414 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 15812 10414 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 15812 10414 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 15893 10414 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 15893 10414 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 15974 10414 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 15974 10414 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 16055 10414 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 16055 10414 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 16136 10414 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 16136 10414 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 16217 10414 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 16217 10414 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 16298 10414 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 16298 10414 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 16379 10414 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 16379 10414 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10350 16460 10414 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10350 16460 10414 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10400 3560 10464 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10400 3560 10464 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10400 3646 10464 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10400 3646 10464 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10400 3732 10464 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10400 3732 10464 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10400 3818 10464 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10400 3818 10464 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10400 3904 10464 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10400 3904 10464 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10400 3990 10464 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10400 3990 10464 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10400 4076 10464 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10400 4076 10464 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10400 4162 10464 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10400 4162 10464 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10400 4248 10464 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10400 4248 10464 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10400 4334 10464 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10400 4334 10464 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10400 4420 10464 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10400 4420 10464 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 13613 10494 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 13613 10494 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 13695 10494 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 13695 10494 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 13777 10494 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 13777 10494 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 13859 10494 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 13859 10494 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 13941 10494 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 13941 10494 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 14023 10494 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 14023 10494 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 14105 10494 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 14105 10494 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 14187 10494 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 14187 10494 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 14269 10494 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 14269 10494 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 14351 10494 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 14351 10494 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 14433 10494 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 14433 10494 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 14515 10494 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 14515 10494 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 14597 10494 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 14597 10494 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 14678 10494 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 14678 10494 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 14759 10494 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 14759 10494 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 14840 10494 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 14840 10494 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 14921 10494 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 14921 10494 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 15002 10494 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 15002 10494 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 15083 10494 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 15083 10494 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 15164 10494 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 15164 10494 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 15245 10494 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 15245 10494 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 15326 10494 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 15326 10494 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 15407 10494 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 15407 10494 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 15488 10494 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 15488 10494 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 15569 10494 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 15569 10494 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 15650 10494 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 15650 10494 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 15731 10494 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 15731 10494 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 15812 10494 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 15812 10494 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 15893 10494 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 15893 10494 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 15974 10494 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 15974 10494 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 16055 10494 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 16055 10494 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 16136 10494 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 16136 10494 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 16217 10494 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 16217 10494 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 16298 10494 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 16298 10494 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 16379 10494 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 16379 10494 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10430 16460 10494 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10430 16460 10494 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10481 3560 10545 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10481 3560 10545 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10481 3646 10545 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10481 3646 10545 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10481 3732 10545 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10481 3732 10545 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10481 3818 10545 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10481 3818 10545 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10481 3904 10545 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10481 3904 10545 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10481 3990 10545 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10481 3990 10545 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10481 4076 10545 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10481 4076 10545 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10481 4162 10545 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10481 4162 10545 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10481 4248 10545 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10481 4248 10545 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10481 4334 10545 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10481 4334 10545 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10481 4420 10545 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10481 4420 10545 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10498 16572 10562 16636 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10498 16572 10562 16636 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10498 16682 10562 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10498 16682 10562 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10498 16792 10562 16856 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10498 16792 10562 16856 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 13613 10574 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 13613 10574 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 13695 10574 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 13695 10574 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 13777 10574 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 13777 10574 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 13859 10574 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 13859 10574 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 13941 10574 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 13941 10574 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 14023 10574 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 14023 10574 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 14105 10574 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 14105 10574 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 14187 10574 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 14187 10574 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 14269 10574 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 14269 10574 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 14351 10574 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 14351 10574 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 14433 10574 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 14433 10574 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 14515 10574 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 14515 10574 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 14597 10574 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 14597 10574 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 14678 10574 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 14678 10574 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 14759 10574 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 14759 10574 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 14840 10574 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 14840 10574 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 14921 10574 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 14921 10574 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 15002 10574 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 15002 10574 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 15083 10574 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 15083 10574 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 15164 10574 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 15164 10574 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 15245 10574 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 15245 10574 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 15326 10574 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 15326 10574 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 15407 10574 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 15407 10574 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 15488 10574 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 15488 10574 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 15569 10574 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 15569 10574 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 15650 10574 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 15650 10574 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 15731 10574 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 15731 10574 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 15812 10574 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 15812 10574 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 15893 10574 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 15893 10574 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 15974 10574 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 15974 10574 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 16055 10574 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 16055 10574 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 16136 10574 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 16136 10574 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 16217 10574 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 16217 10574 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 16298 10574 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 16298 10574 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 16379 10574 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 16379 10574 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10510 16460 10574 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 16460 10574 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10562 3560 10626 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10562 3560 10626 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10562 3646 10626 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10562 3646 10626 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10562 3732 10626 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10562 3732 10626 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10562 3818 10626 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10562 3818 10626 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10562 3904 10626 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10562 3904 10626 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10562 3990 10626 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10562 3990 10626 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10562 4076 10626 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10562 4076 10626 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10562 4162 10626 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10562 4162 10626 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10562 4248 10626 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10562 4248 10626 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10562 4334 10626 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10562 4334 10626 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10562 4420 10626 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10562 4420 10626 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 13613 10654 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 13613 10654 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 13695 10654 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 13695 10654 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 13777 10654 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 13777 10654 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 13859 10654 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 13859 10654 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 13941 10654 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 13941 10654 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 14023 10654 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 14023 10654 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 14105 10654 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 14105 10654 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 14187 10654 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 14187 10654 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 14269 10654 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 14269 10654 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 14351 10654 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 14351 10654 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 14433 10654 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 14433 10654 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 14515 10654 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 14515 10654 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 14597 10654 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 14597 10654 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 14678 10654 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 14678 10654 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 14759 10654 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 14759 10654 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 14840 10654 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 14840 10654 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 14921 10654 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 14921 10654 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 15002 10654 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 15002 10654 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 15083 10654 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 15083 10654 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 15164 10654 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 15164 10654 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 15245 10654 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 15245 10654 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 15326 10654 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 15326 10654 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 15407 10654 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 15407 10654 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 15488 10654 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 15488 10654 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 15569 10654 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 15569 10654 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 15650 10654 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 15650 10654 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 15731 10654 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 15731 10654 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 15812 10654 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 15812 10654 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 15893 10654 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 15893 10654 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 15974 10654 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 15974 10654 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 16055 10654 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 16055 10654 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 16136 10654 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 16136 10654 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 16217 10654 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 16217 10654 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 16298 10654 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 16298 10654 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 16379 10654 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 16379 10654 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10590 16460 10654 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10590 16460 10654 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10643 3560 10707 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10643 3560 10707 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10643 3646 10707 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10643 3646 10707 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10643 3732 10707 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10643 3732 10707 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10643 3818 10707 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10643 3818 10707 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10643 3904 10707 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10643 3904 10707 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10643 3990 10707 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10643 3990 10707 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10643 4076 10707 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10643 4076 10707 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10643 4162 10707 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10643 4162 10707 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10643 4248 10707 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10643 4248 10707 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10643 4334 10707 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10643 4334 10707 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10643 4420 10707 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10643 4420 10707 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10656 16572 10720 16636 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10656 16572 10720 16636 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10656 16682 10720 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10656 16682 10720 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10656 16792 10720 16856 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10656 16792 10720 16856 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 13613 10734 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 13613 10734 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 13695 10734 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 13695 10734 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 13777 10734 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 13777 10734 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 13859 10734 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 13859 10734 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 13941 10734 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 13941 10734 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 14023 10734 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 14023 10734 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 14105 10734 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 14105 10734 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 14187 10734 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 14187 10734 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 14269 10734 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 14269 10734 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 14351 10734 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 14351 10734 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 14433 10734 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 14433 10734 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 14515 10734 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 14515 10734 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 14597 10734 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 14597 10734 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 14678 10734 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 14678 10734 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 14759 10734 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 14759 10734 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 14840 10734 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 14840 10734 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 14921 10734 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 14921 10734 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 15002 10734 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 15002 10734 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 15083 10734 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 15083 10734 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 15164 10734 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 15164 10734 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 15245 10734 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 15245 10734 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 15326 10734 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 15326 10734 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 15407 10734 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 15407 10734 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 15488 10734 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 15488 10734 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 15569 10734 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 15569 10734 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 15650 10734 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 15650 10734 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 15731 10734 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 15731 10734 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 15812 10734 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 15812 10734 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 15893 10734 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 15893 10734 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 15974 10734 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 15974 10734 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 16055 10734 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 16055 10734 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 16136 10734 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 16136 10734 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 16217 10734 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 16217 10734 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 16298 10734 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 16298 10734 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 16379 10734 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 16379 10734 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10670 16460 10734 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10670 16460 10734 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10724 3560 10788 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10724 3560 10788 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10724 3646 10788 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10724 3646 10788 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10724 3732 10788 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10724 3732 10788 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10724 3818 10788 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10724 3818 10788 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10724 3904 10788 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10724 3904 10788 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10724 3990 10788 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10724 3990 10788 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10724 4076 10788 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10724 4076 10788 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10724 4162 10788 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10724 4162 10788 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10724 4248 10788 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10724 4248 10788 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10724 4334 10788 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10724 4334 10788 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10724 4420 10788 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10724 4420 10788 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 13613 10814 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 13613 10814 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 13695 10814 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 13695 10814 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 13777 10814 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 13777 10814 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 13859 10814 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 13859 10814 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 13941 10814 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 13941 10814 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 14023 10814 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 14023 10814 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 14105 10814 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 14105 10814 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 14187 10814 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 14187 10814 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 14269 10814 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 14269 10814 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 14351 10814 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 14351 10814 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 14433 10814 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 14433 10814 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 14515 10814 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 14515 10814 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 14597 10814 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 14597 10814 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 14678 10814 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 14678 10814 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 14759 10814 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 14759 10814 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 14840 10814 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 14840 10814 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 14921 10814 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 14921 10814 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 15002 10814 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 15002 10814 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 15083 10814 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 15083 10814 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 15164 10814 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 15164 10814 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 15245 10814 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 15245 10814 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 15326 10814 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 15326 10814 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 15407 10814 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 15407 10814 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 15488 10814 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 15488 10814 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 15569 10814 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 15569 10814 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 15650 10814 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 15650 10814 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 15731 10814 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 15731 10814 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 15812 10814 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 15812 10814 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 15893 10814 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 15893 10814 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 15974 10814 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 15974 10814 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 16055 10814 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 16055 10814 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 16136 10814 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 16136 10814 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 16217 10814 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 16217 10814 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 16298 10814 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 16298 10814 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 16379 10814 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 16379 10814 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10750 16460 10814 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10750 16460 10814 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10765 16590 10829 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10765 16590 10829 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10765 16682 10829 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10765 16682 10829 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10765 16774 10829 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10765 16774 10829 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10765 16867 10829 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10765 16867 10829 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10765 16960 10829 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10765 16960 10829 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10765 17053 10829 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10765 17053 10829 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10805 3560 10869 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10805 3560 10869 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10805 3646 10869 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10805 3646 10869 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10805 3732 10869 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10805 3732 10869 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10805 3818 10869 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10805 3818 10869 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10805 3904 10869 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10805 3904 10869 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10805 3990 10869 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10805 3990 10869 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10805 4076 10869 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10805 4076 10869 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10805 4162 10869 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10805 4162 10869 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10805 4248 10869 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10805 4248 10869 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10805 4334 10869 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10805 4334 10869 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10805 4420 10869 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10805 4420 10869 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 13613 10894 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 13613 10894 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 13695 10894 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 13695 10894 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 13777 10894 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 13777 10894 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 13859 10894 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 13859 10894 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 13941 10894 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 13941 10894 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 14023 10894 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 14023 10894 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 14105 10894 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 14105 10894 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 14187 10894 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 14187 10894 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 14269 10894 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 14269 10894 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 14351 10894 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 14351 10894 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 14433 10894 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 14433 10894 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 14515 10894 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 14515 10894 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 14597 10894 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 14597 10894 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 14678 10894 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 14678 10894 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 14759 10894 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 14759 10894 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 14840 10894 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 14840 10894 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 14921 10894 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 14921 10894 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 15002 10894 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 15002 10894 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 15083 10894 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 15083 10894 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 15164 10894 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 15164 10894 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 15245 10894 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 15245 10894 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 15326 10894 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 15326 10894 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 15407 10894 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 15407 10894 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 15488 10894 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 15488 10894 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 15569 10894 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 15569 10894 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 15650 10894 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 15650 10894 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 15731 10894 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 15731 10894 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 15812 10894 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 15812 10894 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 15893 10894 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 15893 10894 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 15974 10894 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 15974 10894 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 16055 10894 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 16055 10894 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 16136 10894 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 16136 10894 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 16217 10894 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 16217 10894 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 16298 10894 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 16298 10894 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 16379 10894 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 16379 10894 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10830 16460 10894 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10830 16460 10894 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10861 16590 10925 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10861 16590 10925 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10861 16682 10925 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10861 16682 10925 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10861 16774 10925 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10861 16774 10925 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10861 16867 10925 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10861 16867 10925 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10861 16960 10925 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10861 16960 10925 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10861 17053 10925 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10861 17053 10925 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10886 3560 10950 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10886 3560 10950 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10886 3646 10950 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10886 3646 10950 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10886 3732 10950 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10886 3732 10950 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10886 3818 10950 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10886 3818 10950 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10886 3904 10950 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10886 3904 10950 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10886 3990 10950 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10886 3990 10950 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10886 4076 10950 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10886 4076 10950 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10886 4162 10950 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10886 4162 10950 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10886 4248 10950 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10886 4248 10950 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10886 4334 10950 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10886 4334 10950 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10886 4420 10950 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10886 4420 10950 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 13613 10974 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 13613 10974 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 13695 10974 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 13695 10974 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 13777 10974 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 13777 10974 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 13859 10974 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 13859 10974 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 13941 10974 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 13941 10974 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 14023 10974 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 14023 10974 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 14105 10974 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 14105 10974 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 14187 10974 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 14187 10974 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 14269 10974 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 14269 10974 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 14351 10974 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 14351 10974 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 14433 10974 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 14433 10974 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 14515 10974 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 14515 10974 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 14597 10974 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 14597 10974 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 14678 10974 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 14678 10974 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 14759 10974 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 14759 10974 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 14840 10974 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 14840 10974 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 14921 10974 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 14921 10974 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 15002 10974 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 15002 10974 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 15083 10974 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 15083 10974 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 15164 10974 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 15164 10974 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 15245 10974 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 15245 10974 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 15326 10974 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 15326 10974 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 15407 10974 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 15407 10974 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 15488 10974 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 15488 10974 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 15569 10974 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 15569 10974 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 15650 10974 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 15650 10974 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 15731 10974 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 15731 10974 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 15812 10974 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 15812 10974 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 15893 10974 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 15893 10974 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 15974 10974 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 15974 10974 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 16055 10974 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 16055 10974 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 16136 10974 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 16136 10974 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 16217 10974 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 16217 10974 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 16298 10974 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 16298 10974 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 16379 10974 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 16379 10974 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10910 16460 10974 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10910 16460 10974 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10957 16590 11021 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10957 16590 11021 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10957 16682 11021 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10957 16682 11021 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10957 16774 11021 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10957 16774 11021 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10957 16867 11021 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10957 16867 11021 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10957 16960 11021 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10957 16960 11021 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10957 17053 11021 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10957 17053 11021 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10967 3560 11031 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10967 3560 11031 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10967 3646 11031 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10967 3646 11031 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10967 3732 11031 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10967 3732 11031 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10967 3818 11031 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10967 3818 11031 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10967 3904 11031 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10967 3904 11031 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10967 3990 11031 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10967 3990 11031 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10967 4076 11031 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10967 4076 11031 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10967 4162 11031 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10967 4162 11031 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10967 4248 11031 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10967 4248 11031 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10967 4334 11031 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10967 4334 11031 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10967 4420 11031 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10967 4420 11031 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 13613 11054 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 13613 11054 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 13695 11054 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 13695 11054 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 13777 11054 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 13777 11054 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 13859 11054 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 13859 11054 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 13941 11054 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 13941 11054 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 14023 11054 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 14023 11054 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 14105 11054 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 14105 11054 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 14187 11054 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 14187 11054 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 14269 11054 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 14269 11054 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 14351 11054 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 14351 11054 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 14433 11054 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 14433 11054 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 14515 11054 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 14515 11054 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 14597 11054 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 14597 11054 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 14678 11054 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 14678 11054 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 14759 11054 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 14759 11054 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 14840 11054 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 14840 11054 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 14921 11054 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 14921 11054 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 15002 11054 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 15002 11054 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 15083 11054 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 15083 11054 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 15164 11054 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 15164 11054 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 15245 11054 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 15245 11054 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 15326 11054 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 15326 11054 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 15407 11054 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 15407 11054 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 15488 11054 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 15488 11054 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 15569 11054 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 15569 11054 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 15650 11054 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 15650 11054 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 15731 11054 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 15731 11054 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 15812 11054 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 15812 11054 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 15893 11054 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 15893 11054 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 15974 11054 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 15974 11054 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 16055 11054 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 16055 11054 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 16136 11054 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 16136 11054 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 16217 11054 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 16217 11054 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 16298 11054 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 16298 11054 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 16379 11054 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 16379 11054 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10990 16460 11054 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10990 16460 11054 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11039 17163 11103 17227 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11039 17163 11103 17227 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11039 17250 11103 17314 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11039 17250 11103 17314 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11039 17338 11103 17402 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11039 17338 11103 17402 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11048 3560 11112 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11048 3560 11112 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11048 3646 11112 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11048 3646 11112 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11048 3732 11112 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11048 3732 11112 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11048 3818 11112 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11048 3818 11112 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11048 3904 11112 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11048 3904 11112 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11048 3990 11112 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11048 3990 11112 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11048 4076 11112 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11048 4076 11112 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11048 4162 11112 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11048 4162 11112 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11048 4248 11112 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11048 4248 11112 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11048 4334 11112 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11048 4334 11112 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11048 4420 11112 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11048 4420 11112 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11053 16590 11117 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11053 16590 11117 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11053 16682 11117 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11053 16682 11117 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11053 16774 11117 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11053 16774 11117 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11053 16867 11117 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11053 16867 11117 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11053 16960 11117 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11053 16960 11117 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11053 17053 11117 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11053 17053 11117 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 13613 11134 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 13613 11134 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 13695 11134 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 13695 11134 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 13777 11134 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 13777 11134 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 13859 11134 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 13859 11134 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 13941 11134 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 13941 11134 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 14023 11134 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 14023 11134 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 14105 11134 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 14105 11134 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 14187 11134 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 14187 11134 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 14269 11134 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 14269 11134 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 14351 11134 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 14351 11134 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 14433 11134 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 14433 11134 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 14515 11134 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 14515 11134 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 14597 11134 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 14597 11134 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 14678 11134 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 14678 11134 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 14759 11134 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 14759 11134 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 14840 11134 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 14840 11134 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 14921 11134 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 14921 11134 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 15002 11134 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 15002 11134 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 15083 11134 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 15083 11134 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 15164 11134 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 15164 11134 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 15245 11134 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 15245 11134 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 15326 11134 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 15326 11134 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 15407 11134 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 15407 11134 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 15488 11134 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 15488 11134 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 15569 11134 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 15569 11134 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 15650 11134 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 15650 11134 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 15731 11134 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 15731 11134 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 15812 11134 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 15812 11134 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 15893 11134 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 15893 11134 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 15974 11134 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 15974 11134 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 16055 11134 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 16055 11134 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 16136 11134 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 16136 11134 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 16217 11134 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 16217 11134 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 16298 11134 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 16298 11134 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 16379 11134 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 16379 11134 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11070 16460 11134 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11070 16460 11134 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11129 3560 11193 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11129 3560 11193 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11129 3646 11193 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11129 3646 11193 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11129 3732 11193 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11129 3732 11193 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11129 3818 11193 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11129 3818 11193 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11129 3904 11193 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11129 3904 11193 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11129 3990 11193 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11129 3990 11193 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11129 4076 11193 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11129 4076 11193 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11129 4162 11193 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11129 4162 11193 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11129 4248 11193 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11129 4248 11193 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11129 4334 11193 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11129 4334 11193 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11129 4420 11193 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11129 4420 11193 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11149 16590 11213 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11149 16590 11213 16654 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11149 16682 11213 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11149 16682 11213 16746 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11149 16774 11213 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11149 16774 11213 16838 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11149 16867 11213 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11149 16867 11213 16931 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11149 16960 11213 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11149 16960 11213 17024 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11149 17053 11213 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11149 17053 11213 17117 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 13613 11214 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 13613 11214 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 13695 11214 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 13695 11214 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 13777 11214 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 13777 11214 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 13859 11214 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 13859 11214 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 13941 11214 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 13941 11214 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 14023 11214 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 14023 11214 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 14105 11214 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 14105 11214 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 14187 11214 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 14187 11214 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 14269 11214 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 14269 11214 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 14351 11214 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 14351 11214 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 14433 11214 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 14433 11214 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 14515 11214 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 14515 11214 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 14597 11214 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 14597 11214 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 14678 11214 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 14678 11214 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 14759 11214 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 14759 11214 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 14840 11214 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 14840 11214 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 14921 11214 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 14921 11214 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 15002 11214 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 15002 11214 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 15083 11214 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 15083 11214 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 15164 11214 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 15164 11214 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 15245 11214 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 15245 11214 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 15326 11214 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 15326 11214 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 15407 11214 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 15407 11214 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 15488 11214 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 15488 11214 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 15569 11214 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 15569 11214 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 15650 11214 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 15650 11214 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 15731 11214 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 15731 11214 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 15812 11214 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 15812 11214 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 15893 11214 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 15893 11214 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 15974 11214 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 15974 11214 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 16055 11214 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 16055 11214 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 16136 11214 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 16136 11214 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 16217 11214 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 16217 11214 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 16298 11214 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 16298 11214 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 16379 11214 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 16379 11214 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11150 16460 11214 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11150 16460 11214 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11187 17163 11251 17227 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11187 17163 11251 17227 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11187 17250 11251 17314 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11187 17250 11251 17314 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11187 17338 11251 17402 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11187 17338 11251 17402 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11210 3560 11274 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11210 3560 11274 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11210 3646 11274 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11210 3646 11274 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11210 3732 11274 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11210 3732 11274 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11210 3818 11274 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11210 3818 11274 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11210 3904 11274 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11210 3904 11274 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11210 3990 11274 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11210 3990 11274 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11210 4076 11274 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11210 4076 11274 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11210 4162 11274 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11210 4162 11274 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11210 4248 11274 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11210 4248 11274 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11210 4334 11274 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11210 4334 11274 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11210 4420 11274 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11210 4420 11274 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 13613 11294 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 13613 11294 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 13695 11294 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 13695 11294 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 13777 11294 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 13777 11294 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 13859 11294 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 13859 11294 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 13941 11294 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 13941 11294 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 14023 11294 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 14023 11294 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 14105 11294 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 14105 11294 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 14187 11294 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 14187 11294 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 14269 11294 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 14269 11294 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 14351 11294 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 14351 11294 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 14433 11294 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 14433 11294 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 14515 11294 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 14515 11294 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 14597 11294 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 14597 11294 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 14678 11294 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 14678 11294 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 14759 11294 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 14759 11294 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 14840 11294 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 14840 11294 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 14921 11294 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 14921 11294 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 15002 11294 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 15002 11294 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 15083 11294 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 15083 11294 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 15164 11294 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 15164 11294 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 15245 11294 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 15245 11294 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 15326 11294 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 15326 11294 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 15407 11294 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 15407 11294 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 15488 11294 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 15488 11294 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 15569 11294 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 15569 11294 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 15650 11294 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 15650 11294 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 15731 11294 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 15731 11294 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 15812 11294 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 15812 11294 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 15893 11294 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 15893 11294 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 15974 11294 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 15974 11294 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 16055 11294 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 16055 11294 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 16136 11294 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 16136 11294 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 16217 11294 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 16217 11294 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 16298 11294 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 16298 11294 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 16379 11294 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 16379 11294 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11230 16460 11294 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11230 16460 11294 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11286 16599 11350 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 16599 11350 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11286 16679 11350 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 16679 11350 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11286 16759 11350 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 16759 11350 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11286 16839 11350 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 16839 11350 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11286 16919 11350 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 16919 11350 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11286 16999 11350 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 16999 11350 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11286 17079 11350 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 17079 11350 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11286 17159 11350 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 17159 11350 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11286 17239 11350 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 17239 11350 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11286 17320 11350 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 17320 11350 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11286 17401 11350 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 17401 11350 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11286 17482 11350 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 17482 11350 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11286 17563 11350 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 17563 11350 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11291 3560 11355 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11291 3560 11355 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11291 3646 11355 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11291 3646 11355 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11291 3732 11355 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11291 3732 11355 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11291 3818 11355 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11291 3818 11355 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11291 3904 11355 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11291 3904 11355 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11291 3990 11355 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11291 3990 11355 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11291 4076 11355 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11291 4076 11355 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11291 4162 11355 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11291 4162 11355 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11291 4248 11355 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11291 4248 11355 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11291 4334 11355 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11291 4334 11355 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11291 4420 11355 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11291 4420 11355 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 13613 11374 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 13613 11374 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 13695 11374 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 13695 11374 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 13777 11374 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 13777 11374 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 13859 11374 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 13859 11374 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 13941 11374 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 13941 11374 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 14023 11374 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 14023 11374 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 14105 11374 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 14105 11374 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 14187 11374 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 14187 11374 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 14269 11374 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 14269 11374 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 14351 11374 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 14351 11374 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 14433 11374 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 14433 11374 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 14515 11374 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 14515 11374 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 14597 11374 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 14597 11374 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 14678 11374 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 14678 11374 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 14759 11374 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 14759 11374 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 14840 11374 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 14840 11374 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 14921 11374 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 14921 11374 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 15002 11374 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 15002 11374 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 15083 11374 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 15083 11374 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 15164 11374 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 15164 11374 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 15245 11374 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 15245 11374 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 15326 11374 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 15326 11374 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 15407 11374 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 15407 11374 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 15488 11374 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 15488 11374 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 15569 11374 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 15569 11374 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 15650 11374 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 15650 11374 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 15731 11374 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 15731 11374 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 15812 11374 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 15812 11374 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 15893 11374 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 15893 11374 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 15974 11374 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 15974 11374 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 16055 11374 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 16055 11374 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 16136 11374 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 16136 11374 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 16217 11374 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 16217 11374 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 16298 11374 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 16298 11374 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 16379 11374 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 16379 11374 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11310 16460 11374 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11310 16460 11374 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11368 16599 11432 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 16599 11432 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11368 16679 11432 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 16679 11432 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11368 16759 11432 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 16759 11432 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11368 16839 11432 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 16839 11432 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11368 16919 11432 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 16919 11432 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11368 16999 11432 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 16999 11432 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11368 17079 11432 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 17079 11432 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11368 17159 11432 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 17159 11432 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11368 17239 11432 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 17239 11432 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11368 17320 11432 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 17320 11432 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11368 17401 11432 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 17401 11432 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11368 17482 11432 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 17482 11432 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11368 17563 11432 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 17563 11432 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11372 3560 11436 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11372 3560 11436 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11372 3646 11436 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11372 3646 11436 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11372 3732 11436 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11372 3732 11436 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11372 3818 11436 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11372 3818 11436 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11372 3904 11436 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11372 3904 11436 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11372 3990 11436 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11372 3990 11436 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11372 4076 11436 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11372 4076 11436 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11372 4162 11436 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11372 4162 11436 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11372 4248 11436 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11372 4248 11436 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11372 4334 11436 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11372 4334 11436 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11372 4420 11436 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11372 4420 11436 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 13613 11454 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 13613 11454 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 13695 11454 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 13695 11454 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 13777 11454 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 13777 11454 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 13859 11454 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 13859 11454 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 13941 11454 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 13941 11454 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 14023 11454 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 14023 11454 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 14105 11454 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 14105 11454 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 14187 11454 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 14187 11454 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 14269 11454 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 14269 11454 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 14351 11454 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 14351 11454 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 14433 11454 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 14433 11454 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 14515 11454 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 14515 11454 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 14597 11454 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 14597 11454 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 14678 11454 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 14678 11454 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 14759 11454 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 14759 11454 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 14840 11454 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 14840 11454 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 14921 11454 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 14921 11454 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 15002 11454 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 15002 11454 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 15083 11454 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 15083 11454 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 15164 11454 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 15164 11454 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 15245 11454 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 15245 11454 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 15326 11454 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 15326 11454 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 15407 11454 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 15407 11454 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 15488 11454 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 15488 11454 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 15569 11454 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 15569 11454 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 15650 11454 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 15650 11454 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 15731 11454 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 15731 11454 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 15812 11454 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 15812 11454 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 15893 11454 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 15893 11454 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 15974 11454 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 15974 11454 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 16055 11454 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 16055 11454 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 16136 11454 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 16136 11454 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 16217 11454 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 16217 11454 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 16298 11454 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 16298 11454 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 16379 11454 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 16379 11454 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11390 16460 11454 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11390 16460 11454 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11450 16599 11514 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 16599 11514 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11450 16679 11514 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 16679 11514 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11450 16759 11514 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 16759 11514 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11450 16839 11514 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 16839 11514 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11450 16919 11514 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 16919 11514 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11450 16999 11514 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 16999 11514 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11450 17079 11514 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 17079 11514 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11450 17159 11514 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 17159 11514 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11450 17239 11514 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 17239 11514 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11450 17320 11514 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 17320 11514 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11450 17401 11514 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 17401 11514 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11450 17482 11514 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 17482 11514 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11450 17563 11514 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 17563 11514 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11453 3560 11517 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11453 3560 11517 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11453 3646 11517 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11453 3646 11517 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11453 3732 11517 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11453 3732 11517 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11453 3818 11517 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11453 3818 11517 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11453 3904 11517 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11453 3904 11517 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11453 3990 11517 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11453 3990 11517 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11453 4076 11517 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11453 4076 11517 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11453 4162 11517 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11453 4162 11517 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11453 4248 11517 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11453 4248 11517 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11453 4334 11517 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11453 4334 11517 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11453 4420 11517 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11453 4420 11517 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 13613 11534 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 13613 11534 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 13695 11534 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 13695 11534 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 13777 11534 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 13777 11534 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 13859 11534 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 13859 11534 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 13941 11534 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 13941 11534 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 14023 11534 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 14023 11534 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 14105 11534 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 14105 11534 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 14187 11534 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 14187 11534 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 14269 11534 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 14269 11534 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 14351 11534 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 14351 11534 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 14433 11534 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 14433 11534 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 14515 11534 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 14515 11534 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 14597 11534 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 14597 11534 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 14678 11534 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 14678 11534 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 14759 11534 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 14759 11534 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 14840 11534 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 14840 11534 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 14921 11534 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 14921 11534 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 15002 11534 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 15002 11534 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 15083 11534 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 15083 11534 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 15164 11534 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 15164 11534 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 15245 11534 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 15245 11534 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 15326 11534 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 15326 11534 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 15407 11534 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 15407 11534 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 15488 11534 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 15488 11534 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 15569 11534 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 15569 11534 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 15650 11534 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 15650 11534 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 15731 11534 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 15731 11534 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 15812 11534 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 15812 11534 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 15893 11534 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 15893 11534 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 15974 11534 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 15974 11534 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 16055 11534 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 16055 11534 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 16136 11534 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 16136 11534 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 16217 11534 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 16217 11534 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 16298 11534 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 16298 11534 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 16379 11534 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 16379 11534 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11470 16460 11534 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11470 16460 11534 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11532 16599 11596 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 16599 11596 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11532 16679 11596 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 16679 11596 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11532 16759 11596 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 16759 11596 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11532 16839 11596 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 16839 11596 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11532 16919 11596 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 16919 11596 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11532 16999 11596 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 16999 11596 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11532 17079 11596 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 17079 11596 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11532 17159 11596 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 17159 11596 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11532 17239 11596 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 17239 11596 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11532 17320 11596 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 17320 11596 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11532 17401 11596 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 17401 11596 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11532 17482 11596 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 17482 11596 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11532 17563 11596 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 17563 11596 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11534 3560 11598 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11534 3560 11598 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11534 3646 11598 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11534 3646 11598 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11534 3732 11598 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11534 3732 11598 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11534 3818 11598 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11534 3818 11598 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11534 3904 11598 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11534 3904 11598 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11534 3990 11598 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11534 3990 11598 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11534 4076 11598 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11534 4076 11598 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11534 4162 11598 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11534 4162 11598 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11534 4248 11598 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11534 4248 11598 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11534 4334 11598 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11534 4334 11598 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11534 4420 11598 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11534 4420 11598 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11547 17674 11611 17738 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11547 17674 11611 17738 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11547 17757 11611 17821 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11547 17757 11611 17821 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11547 17841 11611 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11547 17841 11611 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 13613 11614 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 13613 11614 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 13695 11614 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 13695 11614 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 13777 11614 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 13777 11614 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 13859 11614 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 13859 11614 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 13941 11614 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 13941 11614 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 14023 11614 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 14023 11614 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 14105 11614 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 14105 11614 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 14187 11614 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 14187 11614 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 14269 11614 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 14269 11614 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 14351 11614 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 14351 11614 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 14433 11614 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 14433 11614 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 14515 11614 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 14515 11614 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 14597 11614 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 14597 11614 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 14678 11614 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 14678 11614 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 14759 11614 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 14759 11614 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 14840 11614 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 14840 11614 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 14921 11614 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 14921 11614 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 15002 11614 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 15002 11614 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 15083 11614 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 15083 11614 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 15164 11614 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 15164 11614 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 15245 11614 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 15245 11614 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 15326 11614 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 15326 11614 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 15407 11614 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 15407 11614 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 15488 11614 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 15488 11614 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 15569 11614 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 15569 11614 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 15650 11614 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 15650 11614 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 15731 11614 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 15731 11614 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 15812 11614 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 15812 11614 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 15893 11614 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 15893 11614 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 15974 11614 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 15974 11614 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 16055 11614 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 16055 11614 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 16136 11614 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 16136 11614 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 16217 11614 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 16217 11614 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 16298 11614 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 16298 11614 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 16379 11614 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 16379 11614 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11550 16460 11614 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11550 16460 11614 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11614 16599 11678 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 16599 11678 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11614 16679 11678 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 16679 11678 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11614 16759 11678 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 16759 11678 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11614 16839 11678 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 16839 11678 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11614 16919 11678 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 16919 11678 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11614 16999 11678 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 16999 11678 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11614 17079 11678 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 17079 11678 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11614 17159 11678 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 17159 11678 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11614 17239 11678 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 17239 11678 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11614 17320 11678 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 17320 11678 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11614 17401 11678 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 17401 11678 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11614 17482 11678 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 17482 11678 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11614 17563 11678 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 17563 11678 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11615 3560 11679 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11615 3560 11679 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11615 3646 11679 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11615 3646 11679 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11615 3732 11679 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11615 3732 11679 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11615 3818 11679 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11615 3818 11679 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11615 3904 11679 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11615 3904 11679 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11615 3990 11679 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11615 3990 11679 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11615 4076 11679 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11615 4076 11679 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11615 4162 11679 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11615 4162 11679 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11615 4248 11679 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11615 4248 11679 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11615 4334 11679 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11615 4334 11679 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11615 4420 11679 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11615 4420 11679 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 13613 11694 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 13613 11694 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 13695 11694 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 13695 11694 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 13777 11694 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 13777 11694 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 13859 11694 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 13859 11694 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 13941 11694 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 13941 11694 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 14023 11694 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 14023 11694 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 14105 11694 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 14105 11694 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 14187 11694 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 14187 11694 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 14269 11694 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 14269 11694 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 14351 11694 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 14351 11694 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 14433 11694 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 14433 11694 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 14515 11694 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 14515 11694 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 14597 11694 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 14597 11694 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 14678 11694 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 14678 11694 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 14759 11694 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 14759 11694 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 14840 11694 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 14840 11694 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 14921 11694 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 14921 11694 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 15002 11694 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 15002 11694 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 15083 11694 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 15083 11694 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 15164 11694 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 15164 11694 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 15245 11694 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 15245 11694 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 15326 11694 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 15326 11694 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 15407 11694 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 15407 11694 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 15488 11694 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 15488 11694 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 15569 11694 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 15569 11694 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 15650 11694 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 15650 11694 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 15731 11694 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 15731 11694 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 15812 11694 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 15812 11694 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 15893 11694 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 15893 11694 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 15974 11694 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 15974 11694 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 16055 11694 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 16055 11694 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 16136 11694 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 16136 11694 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 16217 11694 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 16217 11694 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 16298 11694 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 16298 11694 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 16379 11694 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 16379 11694 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11630 16460 11694 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11630 16460 11694 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 3560 11760 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 3560 11760 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 3646 11760 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 3646 11760 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 3732 11760 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 3732 11760 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 3818 11760 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 3818 11760 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 3904 11760 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 3904 11760 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 3990 11760 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 3990 11760 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 4076 11760 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 4076 11760 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 4162 11760 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 4162 11760 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 4248 11760 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 4248 11760 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 4334 11760 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 4334 11760 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 4420 11760 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 4420 11760 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 16599 11760 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 16599 11760 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 16679 11760 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 16679 11760 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 16759 11760 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 16759 11760 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 16839 11760 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 16839 11760 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 16919 11760 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 16919 11760 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 16999 11760 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 16999 11760 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 17079 11760 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 17079 11760 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 17159 11760 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 17159 11760 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 17239 11760 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 17239 11760 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 17320 11760 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 17320 11760 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 17401 11760 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 17401 11760 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 17482 11760 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 17482 11760 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11696 17563 11760 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 17563 11760 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11703 17674 11767 17738 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11703 17674 11767 17738 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11703 17757 11767 17821 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11703 17757 11767 17821 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11703 17841 11767 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11703 17841 11767 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 13613 11774 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 13613 11774 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 13695 11774 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 13695 11774 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 13777 11774 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 13777 11774 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 13859 11774 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 13859 11774 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 13941 11774 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 13941 11774 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 14023 11774 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 14023 11774 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 14105 11774 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 14105 11774 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 14187 11774 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 14187 11774 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 14269 11774 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 14269 11774 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 14351 11774 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 14351 11774 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 14433 11774 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 14433 11774 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 14515 11774 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 14515 11774 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 14597 11774 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 14597 11774 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 14678 11774 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 14678 11774 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 14759 11774 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 14759 11774 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 14840 11774 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 14840 11774 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 14921 11774 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 14921 11774 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 15002 11774 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 15002 11774 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 15083 11774 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 15083 11774 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 15164 11774 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 15164 11774 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 15245 11774 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 15245 11774 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 15326 11774 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 15326 11774 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 15407 11774 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 15407 11774 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 15488 11774 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 15488 11774 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 15569 11774 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 15569 11774 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 15650 11774 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 15650 11774 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 15731 11774 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 15731 11774 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 15812 11774 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 15812 11774 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 15893 11774 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 15893 11774 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 15974 11774 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 15974 11774 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 16055 11774 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 16055 11774 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 16136 11774 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 16136 11774 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 16217 11774 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 16217 11774 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 16298 11774 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 16298 11774 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 16379 11774 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 16379 11774 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11710 16460 11774 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11710 16460 11774 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11777 3560 11841 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11777 3560 11841 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11777 3646 11841 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11777 3646 11841 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11777 3732 11841 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11777 3732 11841 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11777 3818 11841 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11777 3818 11841 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11777 3904 11841 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11777 3904 11841 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11777 3990 11841 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11777 3990 11841 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11777 4076 11841 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11777 4076 11841 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11777 4162 11841 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11777 4162 11841 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11777 4248 11841 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11777 4248 11841 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11777 4334 11841 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11777 4334 11841 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11777 4420 11841 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11777 4420 11841 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11778 16599 11842 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 16599 11842 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11778 16679 11842 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 16679 11842 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11778 16759 11842 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 16759 11842 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11778 16839 11842 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 16839 11842 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11778 16919 11842 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 16919 11842 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11778 16999 11842 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 16999 11842 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11778 17079 11842 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 17079 11842 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11778 17159 11842 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 17159 11842 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11778 17239 11842 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 17239 11842 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11778 17320 11842 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 17320 11842 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11778 17401 11842 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 17401 11842 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11778 17482 11842 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 17482 11842 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11778 17563 11842 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 17563 11842 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 13613 11854 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 13613 11854 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 13695 11854 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 13695 11854 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 13777 11854 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 13777 11854 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 13859 11854 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 13859 11854 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 13941 11854 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 13941 11854 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 14023 11854 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 14023 11854 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 14105 11854 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 14105 11854 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 14187 11854 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 14187 11854 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 14269 11854 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 14269 11854 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 14351 11854 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 14351 11854 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 14433 11854 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 14433 11854 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 14515 11854 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 14515 11854 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 14597 11854 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 14597 11854 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 14678 11854 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 14678 11854 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 14759 11854 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 14759 11854 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 14840 11854 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 14840 11854 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 14921 11854 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 14921 11854 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 15002 11854 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 15002 11854 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 15083 11854 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 15083 11854 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 15164 11854 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 15164 11854 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 15245 11854 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 15245 11854 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 15326 11854 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 15326 11854 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 15407 11854 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 15407 11854 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 15488 11854 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 15488 11854 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 15569 11854 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 15569 11854 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 15650 11854 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 15650 11854 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 15731 11854 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 15731 11854 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 15812 11854 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 15812 11854 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 15893 11854 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 15893 11854 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 15974 11854 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 15974 11854 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 16055 11854 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 16055 11854 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 16136 11854 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 16136 11854 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 16217 11854 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 16217 11854 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 16298 11854 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 16298 11854 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 16379 11854 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 16379 11854 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11790 16460 11854 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 16460 11854 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11803 17670 11867 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11803 17670 11867 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11803 17755 11867 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11803 17755 11867 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11803 17841 11867 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11803 17841 11867 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11803 17927 11867 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11803 17927 11867 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11803 18013 11867 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11803 18013 11867 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11803 18099 11867 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11803 18099 11867 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11858 3560 11922 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11858 3560 11922 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11858 3646 11922 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11858 3646 11922 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11858 3732 11922 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11858 3732 11922 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11858 3818 11922 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11858 3818 11922 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11858 3904 11922 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11858 3904 11922 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11858 3990 11922 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11858 3990 11922 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11858 4076 11922 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11858 4076 11922 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11858 4162 11922 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11858 4162 11922 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11858 4248 11922 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11858 4248 11922 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11858 4334 11922 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11858 4334 11922 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11858 4420 11922 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11858 4420 11922 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11860 16599 11924 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 16599 11924 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11860 16679 11924 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 16679 11924 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11860 16759 11924 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 16759 11924 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11860 16839 11924 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 16839 11924 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11860 16919 11924 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 16919 11924 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11860 16999 11924 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 16999 11924 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11860 17079 11924 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 17079 11924 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11860 17159 11924 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 17159 11924 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11860 17239 11924 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 17239 11924 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11860 17320 11924 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 17320 11924 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11860 17401 11924 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 17401 11924 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11860 17482 11924 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 17482 11924 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11860 17563 11924 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 17563 11924 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 13613 11934 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 13613 11934 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 13695 11934 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 13695 11934 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 13777 11934 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 13777 11934 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 13859 11934 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 13859 11934 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 13941 11934 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 13941 11934 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 14023 11934 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 14023 11934 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 14105 11934 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 14105 11934 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 14187 11934 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 14187 11934 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 14269 11934 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 14269 11934 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 14351 11934 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 14351 11934 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 14433 11934 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 14433 11934 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 14515 11934 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 14515 11934 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 14597 11934 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 14597 11934 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 14678 11934 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 14678 11934 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 14759 11934 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 14759 11934 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 14840 11934 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 14840 11934 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 14921 11934 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 14921 11934 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 15002 11934 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 15002 11934 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 15083 11934 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 15083 11934 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 15164 11934 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 15164 11934 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 15245 11934 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 15245 11934 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 15326 11934 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 15326 11934 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 15407 11934 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 15407 11934 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 15488 11934 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 15488 11934 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 15569 11934 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 15569 11934 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 15650 11934 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 15650 11934 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 15731 11934 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 15731 11934 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 15812 11934 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 15812 11934 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 15893 11934 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 15893 11934 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 15974 11934 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 15974 11934 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 16055 11934 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 16055 11934 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 16136 11934 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 16136 11934 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 16217 11934 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 16217 11934 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 16298 11934 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 16298 11934 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 16379 11934 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 16379 11934 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11870 16460 11934 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 16460 11934 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11885 17670 11949 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11885 17670 11949 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11885 17755 11949 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11885 17755 11949 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11885 17841 11949 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11885 17841 11949 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11885 17927 11949 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11885 17927 11949 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11885 18013 11949 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11885 18013 11949 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11885 18099 11949 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11885 18099 11949 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11939 3560 12003 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11939 3560 12003 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11939 3646 12003 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11939 3646 12003 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11939 3732 12003 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11939 3732 12003 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11939 3818 12003 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11939 3818 12003 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11939 3904 12003 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11939 3904 12003 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11939 3990 12003 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11939 3990 12003 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11939 4076 12003 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11939 4076 12003 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11939 4162 12003 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11939 4162 12003 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11939 4248 12003 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11939 4248 12003 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11939 4334 12003 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11939 4334 12003 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11939 4420 12003 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11939 4420 12003 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11942 16599 12006 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 16599 12006 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11942 16679 12006 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 16679 12006 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11942 16759 12006 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 16759 12006 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11942 16839 12006 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 16839 12006 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11942 16919 12006 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 16919 12006 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11942 16999 12006 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 16999 12006 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11942 17079 12006 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 17079 12006 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11942 17159 12006 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 17159 12006 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11942 17239 12006 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 17239 12006 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11942 17320 12006 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 17320 12006 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11942 17401 12006 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 17401 12006 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11942 17482 12006 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 17482 12006 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11942 17563 12006 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 17563 12006 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 13613 12014 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 13613 12014 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 13695 12014 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 13695 12014 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 13777 12014 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 13777 12014 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 13859 12014 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 13859 12014 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 13941 12014 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 13941 12014 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 14023 12014 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 14023 12014 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 14105 12014 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 14105 12014 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 14187 12014 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 14187 12014 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 14269 12014 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 14269 12014 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 14351 12014 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 14351 12014 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 14433 12014 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 14433 12014 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 14515 12014 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 14515 12014 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 14597 12014 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 14597 12014 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 14678 12014 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 14678 12014 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 14759 12014 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 14759 12014 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 14840 12014 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 14840 12014 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 14921 12014 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 14921 12014 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 15002 12014 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 15002 12014 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 15083 12014 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 15083 12014 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 15164 12014 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 15164 12014 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 15245 12014 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 15245 12014 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 15326 12014 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 15326 12014 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 15407 12014 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 15407 12014 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 15488 12014 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 15488 12014 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 15569 12014 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 15569 12014 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 15650 12014 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 15650 12014 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 15731 12014 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 15731 12014 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 15812 12014 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 15812 12014 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 15893 12014 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 15893 12014 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 15974 12014 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 15974 12014 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 16055 12014 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 16055 12014 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 16136 12014 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 16136 12014 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 16217 12014 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 16217 12014 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 16298 12014 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 16298 12014 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 16379 12014 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 16379 12014 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11950 16460 12014 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11950 16460 12014 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11967 17670 12031 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11967 17670 12031 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11967 17755 12031 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11967 17755 12031 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11967 17841 12031 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11967 17841 12031 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11967 17927 12031 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11967 17927 12031 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11967 18013 12031 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11967 18013 12031 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11967 18099 12031 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11967 18099 12031 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11979 18191 12043 18255 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11979 18191 12043 18255 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11979 18277 12043 18341 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11979 18277 12043 18341 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 16559 1265 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16559 1265 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 16641 1265 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16641 1265 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 16723 1265 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16723 1265 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 16805 1265 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16805 1265 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 16887 1265 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16887 1265 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 16969 1265 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16969 1265 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17051 1265 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17051 1265 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17133 1265 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17133 1265 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17215 1265 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17215 1265 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17297 1265 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17297 1265 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17379 1265 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17379 1265 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17461 1265 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17461 1265 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17543 1265 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17543 1265 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17625 1265 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17625 1265 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17707 1265 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17707 1265 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17789 1265 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17789 1265 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17871 1265 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17871 1265 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17953 1265 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17953 1265 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 18035 1265 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18035 1265 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 18117 1265 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18117 1265 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 18199 1265 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18199 1265 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 18281 1265 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18281 1265 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 18363 1265 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18363 1265 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 18445 1265 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18445 1265 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 18527 1265 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18527 1265 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1260 3560 1324 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1260 3560 1324 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1260 3646 1324 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1260 3646 1324 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1260 3732 1324 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1260 3732 1324 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1260 3818 1324 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1260 3818 1324 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1260 3904 1324 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1260 3904 1324 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1260 3990 1324 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1260 3990 1324 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1260 4076 1324 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1260 4076 1324 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1260 4162 1324 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1260 4162 1324 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1260 4248 1324 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1260 4248 1324 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1260 4334 1324 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1260 4334 1324 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1260 4420 1324 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1260 4420 1324 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 13613 1341 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 13613 1341 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 13695 1341 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 13695 1341 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 13777 1341 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 13777 1341 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 13859 1341 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 13859 1341 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 13941 1341 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 13941 1341 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14023 1341 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14023 1341 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14105 1341 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14105 1341 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14187 1341 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14187 1341 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14269 1341 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14269 1341 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14351 1341 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14351 1341 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14433 1341 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14433 1341 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14515 1341 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14515 1341 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14597 1341 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14597 1341 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14678 1341 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14678 1341 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14759 1341 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14759 1341 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14840 1341 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14840 1341 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14921 1341 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14921 1341 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15002 1341 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15002 1341 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15083 1341 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15083 1341 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15164 1341 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15164 1341 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15245 1341 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15245 1341 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15326 1341 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15326 1341 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15407 1341 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15407 1341 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15488 1341 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15488 1341 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15569 1341 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15569 1341 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15650 1341 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15650 1341 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15731 1341 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15731 1341 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15812 1341 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15812 1341 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15893 1341 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15893 1341 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15974 1341 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15974 1341 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 16055 1341 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16055 1341 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 16136 1341 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16136 1341 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 16217 1341 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16217 1341 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 16298 1341 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16298 1341 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 16379 1341 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16379 1341 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 16460 1341 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16460 1341 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 16559 1347 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16559 1347 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 16641 1347 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16641 1347 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 16723 1347 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16723 1347 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 16805 1347 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16805 1347 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 16887 1347 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16887 1347 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 16969 1347 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16969 1347 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17051 1347 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17051 1347 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17133 1347 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17133 1347 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17215 1347 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17215 1347 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17297 1347 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17297 1347 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17379 1347 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17379 1347 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17461 1347 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17461 1347 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17543 1347 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17543 1347 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17625 1347 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17625 1347 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17707 1347 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17707 1347 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17789 1347 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17789 1347 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17871 1347 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17871 1347 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17953 1347 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17953 1347 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 18035 1347 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18035 1347 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 18117 1347 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18117 1347 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 18199 1347 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18199 1347 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 18281 1347 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18281 1347 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 18363 1347 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18363 1347 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 18445 1347 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18445 1347 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 18527 1347 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18527 1347 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1341 3560 1405 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1341 3560 1405 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1341 3646 1405 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1341 3646 1405 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1341 3732 1405 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1341 3732 1405 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1341 3818 1405 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1341 3818 1405 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1341 3904 1405 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1341 3904 1405 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1341 3990 1405 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1341 3990 1405 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1341 4076 1405 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1341 4076 1405 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1341 4162 1405 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1341 4162 1405 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1341 4248 1405 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1341 4248 1405 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1341 4334 1405 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1341 4334 1405 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1341 4420 1405 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1341 4420 1405 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 13613 1421 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 13613 1421 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 13695 1421 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 13695 1421 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 13777 1421 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 13777 1421 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 13859 1421 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 13859 1421 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 13941 1421 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 13941 1421 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14023 1421 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14023 1421 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14105 1421 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14105 1421 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14187 1421 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14187 1421 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14269 1421 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14269 1421 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14351 1421 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14351 1421 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14433 1421 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14433 1421 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14515 1421 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14515 1421 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14597 1421 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14597 1421 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14678 1421 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14678 1421 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14759 1421 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14759 1421 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14840 1421 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14840 1421 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14921 1421 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14921 1421 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15002 1421 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15002 1421 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15083 1421 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15083 1421 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15164 1421 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15164 1421 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15245 1421 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15245 1421 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15326 1421 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15326 1421 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15407 1421 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15407 1421 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15488 1421 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15488 1421 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15569 1421 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15569 1421 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15650 1421 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15650 1421 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15731 1421 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15731 1421 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15812 1421 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15812 1421 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15893 1421 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15893 1421 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15974 1421 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15974 1421 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 16055 1421 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16055 1421 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 16136 1421 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16136 1421 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 16217 1421 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16217 1421 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 16298 1421 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16298 1421 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 16379 1421 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16379 1421 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 16460 1421 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16460 1421 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 16559 1429 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16559 1429 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 16641 1429 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16641 1429 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 16723 1429 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16723 1429 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 16805 1429 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16805 1429 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 16887 1429 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16887 1429 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 16969 1429 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16969 1429 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17051 1429 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17051 1429 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17133 1429 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17133 1429 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17215 1429 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17215 1429 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17297 1429 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17297 1429 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17379 1429 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17379 1429 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17461 1429 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17461 1429 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17543 1429 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17543 1429 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17625 1429 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17625 1429 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17707 1429 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17707 1429 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17789 1429 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17789 1429 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17871 1429 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17871 1429 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17953 1429 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17953 1429 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 18035 1429 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18035 1429 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 18117 1429 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18117 1429 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 18199 1429 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18199 1429 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 18281 1429 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18281 1429 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 18363 1429 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18363 1429 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 18445 1429 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18445 1429 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 18527 1429 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18527 1429 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12020 3560 12084 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12020 3560 12084 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12020 3646 12084 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12020 3646 12084 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12020 3732 12084 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12020 3732 12084 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12020 3818 12084 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12020 3818 12084 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12020 3904 12084 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12020 3904 12084 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12020 3990 12084 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12020 3990 12084 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12020 4076 12084 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12020 4076 12084 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12020 4162 12084 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12020 4162 12084 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12020 4248 12084 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12020 4248 12084 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12020 4334 12084 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12020 4334 12084 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12020 4420 12084 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12020 4420 12084 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12024 16599 12088 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 16599 12088 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12024 16679 12088 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 16679 12088 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12024 16759 12088 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 16759 12088 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12024 16839 12088 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 16839 12088 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12024 16919 12088 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 16919 12088 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12024 16999 12088 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 16999 12088 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12024 17079 12088 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 17079 12088 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12024 17159 12088 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 17159 12088 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12024 17239 12088 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 17239 12088 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12024 17320 12088 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 17320 12088 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12024 17401 12088 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 17401 12088 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12024 17482 12088 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 17482 12088 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12024 17563 12088 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 17563 12088 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 13613 12094 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 13613 12094 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 13695 12094 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 13695 12094 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 13777 12094 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 13777 12094 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 13859 12094 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 13859 12094 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 13941 12094 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 13941 12094 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 14023 12094 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 14023 12094 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 14105 12094 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 14105 12094 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 14187 12094 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 14187 12094 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 14269 12094 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 14269 12094 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 14351 12094 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 14351 12094 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 14433 12094 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 14433 12094 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 14515 12094 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 14515 12094 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 14597 12094 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 14597 12094 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 14678 12094 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 14678 12094 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 14759 12094 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 14759 12094 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 14840 12094 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 14840 12094 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 14921 12094 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 14921 12094 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 15002 12094 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 15002 12094 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 15083 12094 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 15083 12094 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 15164 12094 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 15164 12094 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 15245 12094 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 15245 12094 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 15326 12094 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 15326 12094 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 15407 12094 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 15407 12094 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 15488 12094 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 15488 12094 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 15569 12094 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 15569 12094 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 15650 12094 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 15650 12094 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 15731 12094 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 15731 12094 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 15812 12094 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 15812 12094 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 15893 12094 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 15893 12094 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 15974 12094 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 15974 12094 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 16055 12094 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 16055 12094 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 16136 12094 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 16136 12094 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 16217 12094 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 16217 12094 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 16298 12094 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 16298 12094 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 16379 12094 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 16379 12094 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12030 16460 12094 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12030 16460 12094 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12049 17670 12113 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12049 17670 12113 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12049 17755 12113 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12049 17755 12113 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12049 17841 12113 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12049 17841 12113 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12049 17927 12113 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12049 17927 12113 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12049 18013 12113 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12049 18013 12113 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12049 18099 12113 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12049 18099 12113 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12101 3560 12165 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12101 3560 12165 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12101 3646 12165 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12101 3646 12165 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12101 3732 12165 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12101 3732 12165 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12101 3818 12165 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12101 3818 12165 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12101 3904 12165 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12101 3904 12165 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12101 3990 12165 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12101 3990 12165 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12101 4076 12165 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12101 4076 12165 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12101 4162 12165 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12101 4162 12165 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12101 4248 12165 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12101 4248 12165 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12101 4334 12165 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12101 4334 12165 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12101 4420 12165 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12101 4420 12165 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12106 16599 12170 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 16599 12170 16663 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12106 16679 12170 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 16679 12170 16743 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12106 16759 12170 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 16759 12170 16823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12106 16839 12170 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 16839 12170 16903 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12106 16919 12170 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 16919 12170 16983 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12106 16999 12170 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 16999 12170 17063 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12106 17079 12170 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 17079 12170 17143 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12106 17159 12170 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 17159 12170 17223 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12106 17239 12170 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 17239 12170 17303 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12106 17320 12170 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 17320 12170 17384 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12106 17401 12170 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 17401 12170 17465 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12106 17482 12170 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 17482 12170 17546 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12106 17563 12170 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 17563 12170 17627 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 13613 12174 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 13613 12174 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 13695 12174 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 13695 12174 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 13777 12174 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 13777 12174 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 13859 12174 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 13859 12174 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 13941 12174 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 13941 12174 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 14023 12174 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 14023 12174 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 14105 12174 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 14105 12174 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 14187 12174 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 14187 12174 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 14269 12174 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 14269 12174 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 14351 12174 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 14351 12174 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 14433 12174 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 14433 12174 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 14515 12174 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 14515 12174 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 14597 12174 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 14597 12174 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 14678 12174 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 14678 12174 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 14759 12174 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 14759 12174 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 14840 12174 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 14840 12174 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 14921 12174 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 14921 12174 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 15002 12174 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 15002 12174 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 15083 12174 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 15083 12174 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 15164 12174 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 15164 12174 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 15245 12174 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 15245 12174 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 15326 12174 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 15326 12174 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 15407 12174 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 15407 12174 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 15488 12174 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 15488 12174 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 15569 12174 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 15569 12174 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 15650 12174 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 15650 12174 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 15731 12174 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 15731 12174 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 15812 12174 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 15812 12174 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 15893 12174 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 15893 12174 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 15974 12174 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 15974 12174 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 16055 12174 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 16055 12174 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 16136 12174 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 16136 12174 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 16217 12174 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 16217 12174 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 16298 12174 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 16298 12174 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 16379 12174 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 16379 12174 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12110 16460 12174 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12110 16460 12174 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12131 17670 12195 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12131 17670 12195 17734 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12131 17755 12195 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12131 17755 12195 17819 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12131 17841 12195 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12131 17841 12195 17905 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12131 17927 12195 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12131 17927 12195 17991 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12131 18013 12195 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12131 18013 12195 18077 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12131 18099 12195 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12131 18099 12195 18163 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12135 18191 12199 18255 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12135 18191 12199 18255 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12135 18277 12199 18341 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12135 18277 12199 18341 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12182 3560 12246 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12182 3560 12246 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12182 3646 12246 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12182 3646 12246 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12182 3732 12246 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12182 3732 12246 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12182 3818 12246 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12182 3818 12246 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12182 3904 12246 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12182 3904 12246 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12182 3990 12246 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12182 3990 12246 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12182 4076 12246 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12182 4076 12246 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12182 4162 12246 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12182 4162 12246 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12182 4248 12246 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12182 4248 12246 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12182 4334 12246 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12182 4334 12246 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12182 4420 12246 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12182 4420 12246 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 13613 12254 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 13613 12254 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 13695 12254 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 13695 12254 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 13777 12254 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 13777 12254 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 13859 12254 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 13859 12254 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 13941 12254 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 13941 12254 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 14023 12254 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 14023 12254 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 14105 12254 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 14105 12254 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 14187 12254 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 14187 12254 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 14269 12254 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 14269 12254 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 14351 12254 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 14351 12254 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 14433 12254 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 14433 12254 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 14515 12254 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 14515 12254 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 14597 12254 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 14597 12254 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 14678 12254 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 14678 12254 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 14759 12254 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 14759 12254 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 14840 12254 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 14840 12254 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 14921 12254 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 14921 12254 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 15002 12254 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 15002 12254 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 15083 12254 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 15083 12254 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 15164 12254 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 15164 12254 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 15245 12254 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 15245 12254 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 15326 12254 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 15326 12254 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 15407 12254 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 15407 12254 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 15488 12254 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 15488 12254 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 15569 12254 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 15569 12254 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 15650 12254 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 15650 12254 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 15731 12254 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 15731 12254 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 15812 12254 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 15812 12254 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 15893 12254 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 15893 12254 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 15974 12254 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 15974 12254 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 16055 12254 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 16055 12254 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 16136 12254 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 16136 12254 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 16217 12254 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 16217 12254 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 16298 12254 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 16298 12254 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 16379 12254 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 16379 12254 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12190 16460 12254 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12190 16460 12254 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 16559 12295 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 16559 12295 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 16641 12295 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 16641 12295 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 16723 12295 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 16723 12295 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 16805 12295 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 16805 12295 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 16887 12295 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 16887 12295 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 16969 12295 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 16969 12295 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17051 12295 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17051 12295 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17133 12295 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17133 12295 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17215 12295 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17215 12295 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17297 12295 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17297 12295 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17379 12295 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17379 12295 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17461 12295 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17461 12295 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17543 12295 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17543 12295 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17625 12295 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17625 12295 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17707 12295 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17707 12295 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17789 12295 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17789 12295 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17871 12295 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17871 12295 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17953 12295 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17953 12295 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 18035 12295 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 18035 12295 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 18117 12295 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 18117 12295 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 18199 12295 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 18199 12295 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 18281 12295 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 18281 12295 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 18363 12295 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 18363 12295 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 18445 12295 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 18445 12295 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 18527 12295 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 18527 12295 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12263 3560 12327 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12263 3560 12327 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12263 3646 12327 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12263 3646 12327 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12263 3732 12327 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12263 3732 12327 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12263 3818 12327 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12263 3818 12327 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12263 3904 12327 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12263 3904 12327 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12263 3990 12327 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12263 3990 12327 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12263 4076 12327 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12263 4076 12327 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12263 4162 12327 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12263 4162 12327 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12263 4248 12327 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12263 4248 12327 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12263 4334 12327 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12263 4334 12327 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12263 4420 12327 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12263 4420 12327 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 13613 12334 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 13613 12334 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 13695 12334 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 13695 12334 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 13777 12334 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 13777 12334 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 13859 12334 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 13859 12334 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 13941 12334 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 13941 12334 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 14023 12334 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 14023 12334 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 14105 12334 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 14105 12334 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 14187 12334 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 14187 12334 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 14269 12334 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 14269 12334 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 14351 12334 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 14351 12334 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 14433 12334 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 14433 12334 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 14515 12334 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 14515 12334 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 14597 12334 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 14597 12334 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 14678 12334 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 14678 12334 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 14759 12334 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 14759 12334 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 14840 12334 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 14840 12334 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 14921 12334 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 14921 12334 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 15002 12334 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 15002 12334 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 15083 12334 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 15083 12334 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 15164 12334 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 15164 12334 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 15245 12334 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 15245 12334 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 15326 12334 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 15326 12334 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 15407 12334 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 15407 12334 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 15488 12334 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 15488 12334 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 15569 12334 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 15569 12334 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 15650 12334 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 15650 12334 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 15731 12334 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 15731 12334 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 15812 12334 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 15812 12334 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 15893 12334 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 15893 12334 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 15974 12334 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 15974 12334 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 16055 12334 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 16055 12334 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 16136 12334 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 16136 12334 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 16217 12334 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 16217 12334 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 16298 12334 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 16298 12334 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 16379 12334 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 16379 12334 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12270 16460 12334 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12270 16460 12334 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 16559 12376 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 16559 12376 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 16641 12376 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 16641 12376 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 16723 12376 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 16723 12376 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 16805 12376 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 16805 12376 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 16887 12376 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 16887 12376 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 16969 12376 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 16969 12376 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17051 12376 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17051 12376 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17133 12376 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17133 12376 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17215 12376 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17215 12376 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17297 12376 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17297 12376 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17379 12376 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17379 12376 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17461 12376 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17461 12376 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17543 12376 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17543 12376 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17625 12376 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17625 12376 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17707 12376 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17707 12376 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17789 12376 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17789 12376 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17871 12376 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17871 12376 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17953 12376 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17953 12376 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 18035 12376 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 18035 12376 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 18117 12376 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 18117 12376 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 18199 12376 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 18199 12376 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 18281 12376 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 18281 12376 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 18363 12376 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 18363 12376 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 18445 12376 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 18445 12376 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 18527 12376 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 18527 12376 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12344 3560 12408 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12344 3560 12408 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12344 3646 12408 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12344 3646 12408 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12344 3732 12408 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12344 3732 12408 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12344 3818 12408 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12344 3818 12408 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12344 3904 12408 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12344 3904 12408 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12344 3990 12408 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12344 3990 12408 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12344 4076 12408 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12344 4076 12408 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12344 4162 12408 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12344 4162 12408 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12344 4248 12408 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12344 4248 12408 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12344 4334 12408 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12344 4334 12408 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12344 4420 12408 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12344 4420 12408 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 13613 12414 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 13613 12414 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 13695 12414 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 13695 12414 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 13777 12414 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 13777 12414 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 13859 12414 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 13859 12414 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 13941 12414 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 13941 12414 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 14023 12414 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 14023 12414 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 14105 12414 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 14105 12414 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 14187 12414 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 14187 12414 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 14269 12414 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 14269 12414 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 14351 12414 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 14351 12414 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 14433 12414 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 14433 12414 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 14515 12414 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 14515 12414 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 14597 12414 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 14597 12414 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 14678 12414 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 14678 12414 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 14759 12414 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 14759 12414 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 14840 12414 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 14840 12414 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 14921 12414 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 14921 12414 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 15002 12414 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 15002 12414 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 15083 12414 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 15083 12414 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 15164 12414 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 15164 12414 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 15245 12414 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 15245 12414 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 15326 12414 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 15326 12414 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 15407 12414 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 15407 12414 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 15488 12414 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 15488 12414 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 15569 12414 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 15569 12414 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 15650 12414 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 15650 12414 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 15731 12414 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 15731 12414 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 15812 12414 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 15812 12414 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 15893 12414 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 15893 12414 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 15974 12414 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 15974 12414 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 16055 12414 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 16055 12414 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 16136 12414 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 16136 12414 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 16217 12414 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 16217 12414 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 16298 12414 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 16298 12414 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 16379 12414 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 16379 12414 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12350 16460 12414 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12350 16460 12414 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 16559 12457 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 16559 12457 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 16641 12457 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 16641 12457 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 16723 12457 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 16723 12457 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 16805 12457 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 16805 12457 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 16887 12457 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 16887 12457 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 16969 12457 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 16969 12457 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17051 12457 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17051 12457 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17133 12457 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17133 12457 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17215 12457 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17215 12457 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17297 12457 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17297 12457 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17379 12457 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17379 12457 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17461 12457 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17461 12457 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17543 12457 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17543 12457 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17625 12457 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17625 12457 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17707 12457 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17707 12457 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17789 12457 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17789 12457 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17871 12457 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17871 12457 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17953 12457 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17953 12457 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 18035 12457 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 18035 12457 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 18117 12457 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 18117 12457 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 18199 12457 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 18199 12457 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 18281 12457 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 18281 12457 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 18363 12457 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 18363 12457 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 18445 12457 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 18445 12457 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 18527 12457 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 18527 12457 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12425 3560 12489 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12425 3560 12489 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12425 3646 12489 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12425 3646 12489 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12425 3732 12489 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12425 3732 12489 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12425 3818 12489 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12425 3818 12489 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12425 3904 12489 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12425 3904 12489 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12425 3990 12489 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12425 3990 12489 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12425 4076 12489 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12425 4076 12489 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12425 4162 12489 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12425 4162 12489 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12425 4248 12489 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12425 4248 12489 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12425 4334 12489 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12425 4334 12489 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12425 4420 12489 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12425 4420 12489 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 13613 12494 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 13613 12494 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 13695 12494 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 13695 12494 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 13777 12494 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 13777 12494 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 13859 12494 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 13859 12494 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 13941 12494 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 13941 12494 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 14023 12494 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 14023 12494 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 14105 12494 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 14105 12494 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 14187 12494 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 14187 12494 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 14269 12494 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 14269 12494 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 14351 12494 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 14351 12494 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 14433 12494 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 14433 12494 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 14515 12494 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 14515 12494 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 14597 12494 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 14597 12494 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 14678 12494 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 14678 12494 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 14759 12494 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 14759 12494 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 14840 12494 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 14840 12494 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 14921 12494 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 14921 12494 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 15002 12494 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 15002 12494 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 15083 12494 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 15083 12494 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 15164 12494 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 15164 12494 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 15245 12494 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 15245 12494 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 15326 12494 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 15326 12494 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 15407 12494 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 15407 12494 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 15488 12494 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 15488 12494 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 15569 12494 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 15569 12494 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 15650 12494 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 15650 12494 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 15731 12494 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 15731 12494 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 15812 12494 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 15812 12494 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 15893 12494 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 15893 12494 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 15974 12494 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 15974 12494 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 16055 12494 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 16055 12494 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 16136 12494 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 16136 12494 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 16217 12494 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 16217 12494 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 16298 12494 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 16298 12494 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 16379 12494 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 16379 12494 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12430 16460 12494 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12430 16460 12494 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 16559 12538 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 16559 12538 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 16641 12538 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 16641 12538 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 16723 12538 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 16723 12538 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 16805 12538 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 16805 12538 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 16887 12538 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 16887 12538 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 16969 12538 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 16969 12538 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17051 12538 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17051 12538 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17133 12538 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17133 12538 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17215 12538 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17215 12538 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17297 12538 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17297 12538 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17379 12538 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17379 12538 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17461 12538 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17461 12538 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17543 12538 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17543 12538 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17625 12538 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17625 12538 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17707 12538 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17707 12538 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17789 12538 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17789 12538 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17871 12538 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17871 12538 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17953 12538 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17953 12538 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 18035 12538 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 18035 12538 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 18117 12538 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 18117 12538 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 18199 12538 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 18199 12538 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 18281 12538 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 18281 12538 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 18363 12538 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 18363 12538 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 18445 12538 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 18445 12538 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 18527 12538 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 18527 12538 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12506 3560 12570 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12506 3560 12570 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12506 3646 12570 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12506 3646 12570 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12506 3732 12570 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12506 3732 12570 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12506 3818 12570 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12506 3818 12570 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12506 3904 12570 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12506 3904 12570 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12506 3990 12570 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12506 3990 12570 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12506 4076 12570 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12506 4076 12570 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12506 4162 12570 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12506 4162 12570 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12506 4248 12570 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12506 4248 12570 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12506 4334 12570 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12506 4334 12570 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12506 4420 12570 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12506 4420 12570 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 13613 12574 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 13613 12574 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 13695 12574 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 13695 12574 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 13777 12574 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 13777 12574 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 13859 12574 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 13859 12574 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 13941 12574 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 13941 12574 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 14023 12574 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 14023 12574 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 14105 12574 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 14105 12574 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 14187 12574 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 14187 12574 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 14269 12574 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 14269 12574 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 14351 12574 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 14351 12574 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 14433 12574 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 14433 12574 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 14515 12574 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 14515 12574 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 14597 12574 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 14597 12574 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 14678 12574 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 14678 12574 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 14759 12574 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 14759 12574 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 14840 12574 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 14840 12574 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 14921 12574 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 14921 12574 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 15002 12574 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 15002 12574 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 15083 12574 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 15083 12574 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 15164 12574 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 15164 12574 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 15245 12574 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 15245 12574 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 15326 12574 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 15326 12574 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 15407 12574 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 15407 12574 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 15488 12574 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 15488 12574 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 15569 12574 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 15569 12574 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 15650 12574 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 15650 12574 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 15731 12574 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 15731 12574 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 15812 12574 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 15812 12574 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 15893 12574 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 15893 12574 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 15974 12574 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 15974 12574 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 16055 12574 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 16055 12574 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 16136 12574 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 16136 12574 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 16217 12574 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 16217 12574 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 16298 12574 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 16298 12574 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 16379 12574 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 16379 12574 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12510 16460 12574 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12510 16460 12574 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 16559 12620 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 16559 12620 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 16641 12620 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 16641 12620 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 16723 12620 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 16723 12620 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 16805 12620 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 16805 12620 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 16887 12620 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 16887 12620 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 16969 12620 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 16969 12620 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17051 12620 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17051 12620 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17133 12620 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17133 12620 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17215 12620 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17215 12620 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17297 12620 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17297 12620 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17379 12620 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17379 12620 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17461 12620 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17461 12620 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17543 12620 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17543 12620 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17625 12620 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17625 12620 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17707 12620 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17707 12620 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17789 12620 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17789 12620 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17871 12620 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17871 12620 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17953 12620 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17953 12620 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 18035 12620 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 18035 12620 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 18117 12620 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 18117 12620 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 18199 12620 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 18199 12620 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 18281 12620 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 18281 12620 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 18363 12620 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 18363 12620 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 18445 12620 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 18445 12620 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 18527 12620 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 18527 12620 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12587 3560 12651 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12587 3560 12651 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12587 3646 12651 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12587 3646 12651 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12587 3732 12651 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12587 3732 12651 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12587 3818 12651 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12587 3818 12651 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12587 3904 12651 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12587 3904 12651 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12587 3990 12651 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12587 3990 12651 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12587 4076 12651 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12587 4076 12651 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12587 4162 12651 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12587 4162 12651 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12587 4248 12651 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12587 4248 12651 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12587 4334 12651 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12587 4334 12651 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12587 4420 12651 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12587 4420 12651 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 13613 12654 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 13613 12654 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 13695 12654 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 13695 12654 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 13777 12654 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 13777 12654 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 13859 12654 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 13859 12654 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 13941 12654 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 13941 12654 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 14023 12654 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 14023 12654 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 14105 12654 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 14105 12654 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 14187 12654 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 14187 12654 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 14269 12654 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 14269 12654 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 14351 12654 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 14351 12654 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 14433 12654 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 14433 12654 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 14515 12654 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 14515 12654 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 14597 12654 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 14597 12654 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 14678 12654 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 14678 12654 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 14759 12654 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 14759 12654 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 14840 12654 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 14840 12654 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 14921 12654 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 14921 12654 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 15002 12654 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 15002 12654 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 15083 12654 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 15083 12654 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 15164 12654 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 15164 12654 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 15245 12654 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 15245 12654 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 15326 12654 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 15326 12654 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 15407 12654 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 15407 12654 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 15488 12654 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 15488 12654 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 15569 12654 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 15569 12654 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 15650 12654 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 15650 12654 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 15731 12654 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 15731 12654 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 15812 12654 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 15812 12654 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 15893 12654 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 15893 12654 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 15974 12654 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 15974 12654 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 16055 12654 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 16055 12654 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 16136 12654 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 16136 12654 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 16217 12654 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 16217 12654 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 16298 12654 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 16298 12654 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 16379 12654 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 16379 12654 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12590 16460 12654 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12590 16460 12654 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 16559 12702 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 16559 12702 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 16641 12702 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 16641 12702 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 16723 12702 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 16723 12702 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 16805 12702 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 16805 12702 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 16887 12702 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 16887 12702 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 16969 12702 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 16969 12702 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17051 12702 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17051 12702 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17133 12702 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17133 12702 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17215 12702 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17215 12702 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17297 12702 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17297 12702 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17379 12702 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17379 12702 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17461 12702 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17461 12702 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17543 12702 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17543 12702 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17625 12702 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17625 12702 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17707 12702 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17707 12702 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17789 12702 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17789 12702 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17871 12702 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17871 12702 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17953 12702 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17953 12702 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 18035 12702 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 18035 12702 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 18117 12702 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 18117 12702 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 18199 12702 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 18199 12702 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 18281 12702 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 18281 12702 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 18363 12702 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 18363 12702 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 18445 12702 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 18445 12702 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 18527 12702 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 18527 12702 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12668 3560 12732 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12668 3560 12732 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12668 3646 12732 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12668 3646 12732 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12668 3732 12732 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12668 3732 12732 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12668 3818 12732 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12668 3818 12732 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12668 3904 12732 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12668 3904 12732 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12668 3990 12732 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12668 3990 12732 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12668 4076 12732 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12668 4076 12732 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12668 4162 12732 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12668 4162 12732 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12668 4248 12732 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12668 4248 12732 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12668 4334 12732 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12668 4334 12732 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12668 4420 12732 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12668 4420 12732 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 13613 12734 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 13613 12734 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 13695 12734 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 13695 12734 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 13777 12734 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 13777 12734 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 13859 12734 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 13859 12734 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 13941 12734 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 13941 12734 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 14023 12734 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 14023 12734 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 14105 12734 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 14105 12734 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 14187 12734 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 14187 12734 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 14269 12734 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 14269 12734 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 14351 12734 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 14351 12734 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 14433 12734 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 14433 12734 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 14515 12734 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 14515 12734 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 14597 12734 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 14597 12734 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 14678 12734 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 14678 12734 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 14759 12734 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 14759 12734 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 14840 12734 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 14840 12734 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 14921 12734 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 14921 12734 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 15002 12734 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 15002 12734 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 15083 12734 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 15083 12734 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 15164 12734 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 15164 12734 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 15245 12734 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 15245 12734 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 15326 12734 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 15326 12734 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 15407 12734 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 15407 12734 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 15488 12734 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 15488 12734 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 15569 12734 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 15569 12734 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 15650 12734 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 15650 12734 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 15731 12734 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 15731 12734 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 15812 12734 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 15812 12734 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 15893 12734 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 15893 12734 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 15974 12734 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 15974 12734 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 16055 12734 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 16055 12734 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 16136 12734 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 16136 12734 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 16217 12734 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 16217 12734 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 16298 12734 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 16298 12734 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 16379 12734 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 16379 12734 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12670 16460 12734 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12670 16460 12734 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 16559 12784 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 16559 12784 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 16641 12784 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 16641 12784 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 16723 12784 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 16723 12784 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 16805 12784 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 16805 12784 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 16887 12784 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 16887 12784 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 16969 12784 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 16969 12784 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17051 12784 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17051 12784 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17133 12784 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17133 12784 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17215 12784 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17215 12784 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17297 12784 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17297 12784 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17379 12784 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17379 12784 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17461 12784 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17461 12784 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17543 12784 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17543 12784 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17625 12784 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17625 12784 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17707 12784 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17707 12784 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17789 12784 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17789 12784 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17871 12784 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17871 12784 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17953 12784 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17953 12784 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 18035 12784 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 18035 12784 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 18117 12784 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 18117 12784 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 18199 12784 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 18199 12784 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 18281 12784 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 18281 12784 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 18363 12784 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 18363 12784 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 18445 12784 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 18445 12784 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 18527 12784 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 18527 12784 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12749 3560 12813 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12749 3560 12813 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12749 3646 12813 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12749 3646 12813 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12749 3732 12813 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12749 3732 12813 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12749 3818 12813 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12749 3818 12813 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12749 3904 12813 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12749 3904 12813 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12749 3990 12813 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12749 3990 12813 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12749 4076 12813 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12749 4076 12813 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12749 4162 12813 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12749 4162 12813 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12749 4248 12813 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12749 4248 12813 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12749 4334 12813 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12749 4334 12813 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12749 4420 12813 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12749 4420 12813 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 13613 12814 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 13613 12814 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 13695 12814 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 13695 12814 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 13777 12814 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 13777 12814 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 13859 12814 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 13859 12814 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 13941 12814 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 13941 12814 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 14023 12814 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 14023 12814 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 14105 12814 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 14105 12814 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 14187 12814 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 14187 12814 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 14269 12814 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 14269 12814 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 14351 12814 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 14351 12814 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 14433 12814 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 14433 12814 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 14515 12814 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 14515 12814 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 14597 12814 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 14597 12814 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 14678 12814 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 14678 12814 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 14759 12814 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 14759 12814 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 14840 12814 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 14840 12814 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 14921 12814 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 14921 12814 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 15002 12814 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 15002 12814 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 15083 12814 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 15083 12814 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 15164 12814 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 15164 12814 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 15245 12814 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 15245 12814 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 15326 12814 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 15326 12814 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 15407 12814 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 15407 12814 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 15488 12814 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 15488 12814 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 15569 12814 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 15569 12814 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 15650 12814 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 15650 12814 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 15731 12814 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 15731 12814 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 15812 12814 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 15812 12814 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 15893 12814 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 15893 12814 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 15974 12814 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 15974 12814 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 16055 12814 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 16055 12814 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 16136 12814 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 16136 12814 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 16217 12814 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 16217 12814 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 16298 12814 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 16298 12814 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 16379 12814 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 16379 12814 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12750 16460 12814 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12750 16460 12814 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 16559 12866 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 16559 12866 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 16641 12866 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 16641 12866 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 16723 12866 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 16723 12866 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 16805 12866 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 16805 12866 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 16887 12866 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 16887 12866 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 16969 12866 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 16969 12866 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17051 12866 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17051 12866 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17133 12866 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17133 12866 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17215 12866 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17215 12866 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17297 12866 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17297 12866 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17379 12866 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17379 12866 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17461 12866 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17461 12866 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17543 12866 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17543 12866 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17625 12866 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17625 12866 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17707 12866 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17707 12866 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17789 12866 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17789 12866 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17871 12866 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17871 12866 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17953 12866 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17953 12866 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 18035 12866 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 18035 12866 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 18117 12866 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 18117 12866 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 18199 12866 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 18199 12866 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 18281 12866 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 18281 12866 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 18363 12866 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 18363 12866 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 18445 12866 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 18445 12866 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 18527 12866 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 18527 12866 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 3560 12894 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 3560 12894 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 3646 12894 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 3646 12894 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 3732 12894 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 3732 12894 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 3818 12894 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 3818 12894 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 3904 12894 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 3904 12894 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 3990 12894 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 3990 12894 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 4076 12894 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 4076 12894 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 4162 12894 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 4162 12894 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 4248 12894 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 4248 12894 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 4334 12894 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 4334 12894 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 4420 12894 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 4420 12894 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 13613 12894 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 13613 12894 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 13695 12894 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 13695 12894 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 13777 12894 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 13777 12894 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 13859 12894 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 13859 12894 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 13941 12894 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 13941 12894 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 14023 12894 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 14023 12894 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 14105 12894 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 14105 12894 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 14187 12894 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 14187 12894 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 14269 12894 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 14269 12894 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 14351 12894 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 14351 12894 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 14433 12894 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 14433 12894 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 14515 12894 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 14515 12894 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 14597 12894 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 14597 12894 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 14678 12894 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 14678 12894 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 14759 12894 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 14759 12894 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 14840 12894 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 14840 12894 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 14921 12894 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 14921 12894 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 15002 12894 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 15002 12894 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 15083 12894 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 15083 12894 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 15164 12894 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 15164 12894 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 15245 12894 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 15245 12894 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 15326 12894 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 15326 12894 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 15407 12894 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 15407 12894 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 15488 12894 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 15488 12894 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 15569 12894 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 15569 12894 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 15650 12894 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 15650 12894 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 15731 12894 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 15731 12894 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 15812 12894 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 15812 12894 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 15893 12894 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 15893 12894 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 15974 12894 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 15974 12894 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 16055 12894 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 16055 12894 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 16136 12894 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 16136 12894 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 16217 12894 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 16217 12894 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 16298 12894 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 16298 12894 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 16379 12894 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 16379 12894 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12830 16460 12894 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12830 16460 12894 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 16559 12948 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 16559 12948 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 16641 12948 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 16641 12948 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 16723 12948 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 16723 12948 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 16805 12948 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 16805 12948 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 16887 12948 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 16887 12948 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 16969 12948 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 16969 12948 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17051 12948 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17051 12948 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17133 12948 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17133 12948 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17215 12948 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17215 12948 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17297 12948 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17297 12948 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17379 12948 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17379 12948 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17461 12948 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17461 12948 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17543 12948 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17543 12948 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17625 12948 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17625 12948 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17707 12948 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17707 12948 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17789 12948 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17789 12948 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17871 12948 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17871 12948 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17953 12948 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17953 12948 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 18035 12948 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 18035 12948 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 18117 12948 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 18117 12948 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 18199 12948 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 18199 12948 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 18281 12948 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 18281 12948 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 18363 12948 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 18363 12948 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 18445 12948 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 18445 12948 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 18527 12948 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 18527 12948 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 13613 12974 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 13613 12974 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 13695 12974 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 13695 12974 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 13777 12974 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 13777 12974 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 13859 12974 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 13859 12974 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 13941 12974 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 13941 12974 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 14023 12974 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 14023 12974 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 14105 12974 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 14105 12974 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 14187 12974 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 14187 12974 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 14269 12974 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 14269 12974 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 14351 12974 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 14351 12974 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 14433 12974 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 14433 12974 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 14515 12974 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 14515 12974 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 14597 12974 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 14597 12974 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 14678 12974 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 14678 12974 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 14759 12974 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 14759 12974 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 14840 12974 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 14840 12974 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 14921 12974 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 14921 12974 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 15002 12974 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 15002 12974 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 15083 12974 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 15083 12974 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 15164 12974 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 15164 12974 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 15245 12974 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 15245 12974 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 15326 12974 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 15326 12974 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 15407 12974 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 15407 12974 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 15488 12974 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 15488 12974 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 15569 12974 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 15569 12974 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 15650 12974 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 15650 12974 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 15731 12974 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 15731 12974 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 15812 12974 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 15812 12974 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 15893 12974 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 15893 12974 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 15974 12974 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 15974 12974 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 16055 12974 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 16055 12974 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 16136 12974 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 16136 12974 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 16217 12974 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 16217 12974 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 16298 12974 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 16298 12974 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 16379 12974 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 16379 12974 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12910 16460 12974 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12910 16460 12974 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12911 3560 12975 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12911 3560 12975 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12911 3646 12975 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12911 3646 12975 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12911 3732 12975 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12911 3732 12975 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12911 3818 12975 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12911 3818 12975 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12911 3904 12975 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12911 3904 12975 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12911 3990 12975 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12911 3990 12975 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12911 4076 12975 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12911 4076 12975 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12911 4162 12975 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12911 4162 12975 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12911 4248 12975 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12911 4248 12975 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12911 4334 12975 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12911 4334 12975 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12911 4420 12975 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12911 4420 12975 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 16559 13030 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 16559 13030 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 16641 13030 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 16641 13030 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 16723 13030 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 16723 13030 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 16805 13030 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 16805 13030 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 16887 13030 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 16887 13030 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 16969 13030 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 16969 13030 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17051 13030 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17051 13030 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17133 13030 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17133 13030 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17215 13030 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17215 13030 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17297 13030 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17297 13030 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17379 13030 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17379 13030 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17461 13030 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17461 13030 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17543 13030 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17543 13030 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17625 13030 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17625 13030 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17707 13030 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17707 13030 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17789 13030 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17789 13030 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17871 13030 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17871 13030 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17953 13030 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17953 13030 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 18035 13030 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 18035 13030 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 18117 13030 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 18117 13030 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 18199 13030 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 18199 13030 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 18281 13030 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 18281 13030 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 18363 13030 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 18363 13030 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 18445 13030 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 18445 13030 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 18527 13030 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 18527 13030 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 13613 13054 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 13613 13054 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 13695 13054 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 13695 13054 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 13777 13054 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 13777 13054 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 13859 13054 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 13859 13054 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 13941 13054 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 13941 13054 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 14023 13054 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 14023 13054 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 14105 13054 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 14105 13054 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 14187 13054 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 14187 13054 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 14269 13054 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 14269 13054 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 14351 13054 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 14351 13054 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 14433 13054 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 14433 13054 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 14515 13054 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 14515 13054 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 14597 13054 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 14597 13054 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 14678 13054 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 14678 13054 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 14759 13054 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 14759 13054 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 14840 13054 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 14840 13054 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 14921 13054 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 14921 13054 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 15002 13054 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 15002 13054 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 15083 13054 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 15083 13054 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 15164 13054 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 15164 13054 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 15245 13054 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 15245 13054 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 15326 13054 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 15326 13054 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 15407 13054 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 15407 13054 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 15488 13054 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 15488 13054 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 15569 13054 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 15569 13054 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 15650 13054 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 15650 13054 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 15731 13054 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 15731 13054 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 15812 13054 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 15812 13054 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 15893 13054 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 15893 13054 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 15974 13054 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 15974 13054 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 16055 13054 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 16055 13054 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 16136 13054 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 16136 13054 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 16217 13054 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 16217 13054 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 16298 13054 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 16298 13054 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 16379 13054 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 16379 13054 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12990 16460 13054 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12990 16460 13054 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12992 3560 13056 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12992 3560 13056 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12992 3646 13056 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12992 3646 13056 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12992 3732 13056 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12992 3732 13056 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12992 3818 13056 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12992 3818 13056 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12992 3904 13056 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12992 3904 13056 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12992 3990 13056 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12992 3990 13056 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12992 4076 13056 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12992 4076 13056 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12992 4162 13056 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12992 4162 13056 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12992 4248 13056 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12992 4248 13056 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12992 4334 13056 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12992 4334 13056 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12992 4420 13056 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12992 4420 13056 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 16559 13112 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 16559 13112 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 16641 13112 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 16641 13112 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 16723 13112 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 16723 13112 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 16805 13112 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 16805 13112 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 16887 13112 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 16887 13112 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 16969 13112 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 16969 13112 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17051 13112 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17051 13112 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17133 13112 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17133 13112 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17215 13112 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17215 13112 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17297 13112 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17297 13112 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17379 13112 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17379 13112 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17461 13112 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17461 13112 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17543 13112 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17543 13112 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17625 13112 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17625 13112 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17707 13112 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17707 13112 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17789 13112 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17789 13112 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17871 13112 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17871 13112 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17953 13112 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17953 13112 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 18035 13112 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 18035 13112 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 18117 13112 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 18117 13112 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 18199 13112 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 18199 13112 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 18281 13112 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 18281 13112 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 18363 13112 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 18363 13112 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 18445 13112 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 18445 13112 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 18527 13112 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 18527 13112 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 13613 13134 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 13613 13134 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 13695 13134 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 13695 13134 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 13777 13134 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 13777 13134 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 13859 13134 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 13859 13134 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 13941 13134 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 13941 13134 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 14023 13134 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 14023 13134 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 14105 13134 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 14105 13134 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 14187 13134 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 14187 13134 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 14269 13134 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 14269 13134 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 14351 13134 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 14351 13134 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 14433 13134 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 14433 13134 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 14515 13134 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 14515 13134 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 14597 13134 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 14597 13134 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 14678 13134 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 14678 13134 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 14759 13134 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 14759 13134 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 14840 13134 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 14840 13134 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 14921 13134 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 14921 13134 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 15002 13134 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 15002 13134 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 15083 13134 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 15083 13134 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 15164 13134 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 15164 13134 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 15245 13134 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 15245 13134 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 15326 13134 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 15326 13134 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 15407 13134 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 15407 13134 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 15488 13134 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 15488 13134 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 15569 13134 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 15569 13134 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 15650 13134 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 15650 13134 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 15731 13134 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 15731 13134 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 15812 13134 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 15812 13134 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 15893 13134 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 15893 13134 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 15974 13134 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 15974 13134 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 16055 13134 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 16055 13134 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 16136 13134 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 16136 13134 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 16217 13134 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 16217 13134 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 16298 13134 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 16298 13134 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 16379 13134 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 16379 13134 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13070 16460 13134 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13070 16460 13134 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13073 3560 13137 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13073 3560 13137 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13073 3646 13137 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13073 3646 13137 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13073 3732 13137 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13073 3732 13137 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13073 3818 13137 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13073 3818 13137 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13073 3904 13137 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13073 3904 13137 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13073 3990 13137 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13073 3990 13137 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13073 4076 13137 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13073 4076 13137 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13073 4162 13137 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13073 4162 13137 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13073 4248 13137 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13073 4248 13137 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13073 4334 13137 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13073 4334 13137 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13073 4420 13137 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13073 4420 13137 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 16559 13194 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 16559 13194 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 16641 13194 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 16641 13194 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 16723 13194 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 16723 13194 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 16805 13194 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 16805 13194 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 16887 13194 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 16887 13194 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 16969 13194 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 16969 13194 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17051 13194 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17051 13194 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17133 13194 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17133 13194 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17215 13194 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17215 13194 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17297 13194 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17297 13194 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17379 13194 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17379 13194 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17461 13194 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17461 13194 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17543 13194 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17543 13194 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17625 13194 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17625 13194 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17707 13194 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17707 13194 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17789 13194 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17789 13194 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17871 13194 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17871 13194 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17953 13194 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17953 13194 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 18035 13194 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 18035 13194 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 18117 13194 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 18117 13194 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 18199 13194 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 18199 13194 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 18281 13194 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 18281 13194 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 18363 13194 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 18363 13194 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 18445 13194 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 18445 13194 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 18527 13194 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 18527 13194 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 13613 13214 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 13613 13214 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 13695 13214 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 13695 13214 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 13777 13214 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 13777 13214 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 13859 13214 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 13859 13214 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 13941 13214 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 13941 13214 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 14023 13214 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 14023 13214 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 14105 13214 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 14105 13214 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 14187 13214 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 14187 13214 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 14269 13214 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 14269 13214 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 14351 13214 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 14351 13214 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 14433 13214 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 14433 13214 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 14515 13214 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 14515 13214 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 14597 13214 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 14597 13214 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 14678 13214 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 14678 13214 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 14759 13214 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 14759 13214 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 14840 13214 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 14840 13214 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 14921 13214 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 14921 13214 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 15002 13214 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 15002 13214 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 15083 13214 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 15083 13214 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 15164 13214 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 15164 13214 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 15245 13214 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 15245 13214 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 15326 13214 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 15326 13214 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 15407 13214 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 15407 13214 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 15488 13214 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 15488 13214 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 15569 13214 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 15569 13214 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 15650 13214 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 15650 13214 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 15731 13214 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 15731 13214 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 15812 13214 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 15812 13214 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 15893 13214 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 15893 13214 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 15974 13214 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 15974 13214 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 16055 13214 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 16055 13214 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 16136 13214 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 16136 13214 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 16217 13214 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 16217 13214 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 16298 13214 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 16298 13214 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 16379 13214 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 16379 13214 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13150 16460 13214 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13150 16460 13214 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13154 3560 13218 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13154 3560 13218 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13154 3646 13218 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13154 3646 13218 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13154 3732 13218 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13154 3732 13218 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13154 3818 13218 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13154 3818 13218 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13154 3904 13218 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13154 3904 13218 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13154 3990 13218 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13154 3990 13218 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13154 4076 13218 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13154 4076 13218 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13154 4162 13218 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13154 4162 13218 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13154 4248 13218 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13154 4248 13218 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13154 4334 13218 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13154 4334 13218 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13154 4420 13218 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13154 4420 13218 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 16559 13276 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 16559 13276 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 16641 13276 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 16641 13276 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 16723 13276 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 16723 13276 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 16805 13276 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 16805 13276 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 16887 13276 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 16887 13276 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 16969 13276 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 16969 13276 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17051 13276 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17051 13276 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17133 13276 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17133 13276 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17215 13276 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17215 13276 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17297 13276 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17297 13276 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17379 13276 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17379 13276 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17461 13276 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17461 13276 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17543 13276 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17543 13276 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17625 13276 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17625 13276 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17707 13276 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17707 13276 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17789 13276 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17789 13276 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17871 13276 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17871 13276 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17953 13276 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17953 13276 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 18035 13276 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 18035 13276 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 18117 13276 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 18117 13276 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 18199 13276 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 18199 13276 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 18281 13276 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 18281 13276 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 18363 13276 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 18363 13276 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 18445 13276 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 18445 13276 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 18527 13276 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 18527 13276 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 13613 13294 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 13613 13294 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 13695 13294 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 13695 13294 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 13777 13294 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 13777 13294 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 13859 13294 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 13859 13294 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 13941 13294 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 13941 13294 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 14023 13294 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 14023 13294 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 14105 13294 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 14105 13294 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 14187 13294 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 14187 13294 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 14269 13294 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 14269 13294 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 14351 13294 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 14351 13294 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 14433 13294 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 14433 13294 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 14515 13294 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 14515 13294 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 14597 13294 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 14597 13294 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 14678 13294 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 14678 13294 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 14759 13294 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 14759 13294 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 14840 13294 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 14840 13294 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 14921 13294 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 14921 13294 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 15002 13294 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 15002 13294 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 15083 13294 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 15083 13294 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 15164 13294 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 15164 13294 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 15245 13294 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 15245 13294 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 15326 13294 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 15326 13294 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 15407 13294 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 15407 13294 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 15488 13294 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 15488 13294 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 15569 13294 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 15569 13294 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 15650 13294 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 15650 13294 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 15731 13294 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 15731 13294 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 15812 13294 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 15812 13294 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 15893 13294 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 15893 13294 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 15974 13294 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 15974 13294 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 16055 13294 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 16055 13294 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 16136 13294 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 16136 13294 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 16217 13294 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 16217 13294 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 16298 13294 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 16298 13294 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 16379 13294 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 16379 13294 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13230 16460 13294 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13230 16460 13294 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13235 3560 13299 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13235 3560 13299 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13235 3646 13299 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13235 3646 13299 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13235 3732 13299 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13235 3732 13299 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13235 3818 13299 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13235 3818 13299 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13235 3904 13299 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13235 3904 13299 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13235 3990 13299 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13235 3990 13299 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13235 4076 13299 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13235 4076 13299 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13235 4162 13299 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13235 4162 13299 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13235 4248 13299 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13235 4248 13299 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13235 4334 13299 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13235 4334 13299 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13235 4420 13299 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13235 4420 13299 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 16559 13358 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 16559 13358 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 16641 13358 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 16641 13358 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 16723 13358 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 16723 13358 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 16805 13358 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 16805 13358 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 16887 13358 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 16887 13358 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 16969 13358 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 16969 13358 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17051 13358 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17051 13358 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17133 13358 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17133 13358 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17215 13358 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17215 13358 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17297 13358 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17297 13358 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17379 13358 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17379 13358 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17461 13358 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17461 13358 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17543 13358 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17543 13358 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17625 13358 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17625 13358 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17707 13358 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17707 13358 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17789 13358 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17789 13358 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17871 13358 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17871 13358 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17953 13358 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17953 13358 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 18035 13358 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 18035 13358 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 18117 13358 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 18117 13358 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 18199 13358 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 18199 13358 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 18281 13358 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 18281 13358 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 18363 13358 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 18363 13358 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 18445 13358 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 18445 13358 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 18527 13358 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 18527 13358 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 13613 13374 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 13613 13374 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 13695 13374 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 13695 13374 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 13777 13374 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 13777 13374 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 13859 13374 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 13859 13374 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 13941 13374 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 13941 13374 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 14023 13374 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 14023 13374 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 14105 13374 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 14105 13374 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 14187 13374 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 14187 13374 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 14269 13374 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 14269 13374 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 14351 13374 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 14351 13374 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 14433 13374 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 14433 13374 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 14515 13374 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 14515 13374 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 14597 13374 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 14597 13374 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 14678 13374 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 14678 13374 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 14759 13374 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 14759 13374 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 14840 13374 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 14840 13374 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 14921 13374 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 14921 13374 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 15002 13374 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 15002 13374 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 15083 13374 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 15083 13374 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 15164 13374 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 15164 13374 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 15245 13374 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 15245 13374 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 15326 13374 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 15326 13374 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 15407 13374 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 15407 13374 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 15488 13374 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 15488 13374 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 15569 13374 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 15569 13374 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 15650 13374 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 15650 13374 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 15731 13374 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 15731 13374 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 15812 13374 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 15812 13374 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 15893 13374 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 15893 13374 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 15974 13374 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 15974 13374 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 16055 13374 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 16055 13374 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 16136 13374 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 16136 13374 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 16217 13374 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 16217 13374 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 16298 13374 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 16298 13374 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 16379 13374 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 16379 13374 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13310 16460 13374 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13310 16460 13374 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13316 3560 13380 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13316 3560 13380 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13316 3646 13380 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13316 3646 13380 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13316 3732 13380 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13316 3732 13380 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13316 3818 13380 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13316 3818 13380 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13316 3904 13380 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13316 3904 13380 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13316 3990 13380 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13316 3990 13380 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13316 4076 13380 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13316 4076 13380 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13316 4162 13380 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13316 4162 13380 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13316 4248 13380 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13316 4248 13380 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13316 4334 13380 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13316 4334 13380 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13316 4420 13380 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13316 4420 13380 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 16559 13440 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 16559 13440 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 16641 13440 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 16641 13440 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 16723 13440 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 16723 13440 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 16805 13440 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 16805 13440 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 16887 13440 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 16887 13440 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 16969 13440 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 16969 13440 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17051 13440 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17051 13440 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17133 13440 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17133 13440 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17215 13440 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17215 13440 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17297 13440 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17297 13440 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17379 13440 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17379 13440 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17461 13440 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17461 13440 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17543 13440 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17543 13440 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17625 13440 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17625 13440 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17707 13440 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17707 13440 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17789 13440 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17789 13440 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17871 13440 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17871 13440 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17953 13440 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17953 13440 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 18035 13440 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 18035 13440 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 18117 13440 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 18117 13440 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 18199 13440 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 18199 13440 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 18281 13440 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 18281 13440 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 18363 13440 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 18363 13440 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 18445 13440 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 18445 13440 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 18527 13440 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 18527 13440 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 13613 13454 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 13613 13454 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 13695 13454 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 13695 13454 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 13777 13454 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 13777 13454 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 13859 13454 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 13859 13454 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 13941 13454 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 13941 13454 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 14023 13454 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 14023 13454 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 14105 13454 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 14105 13454 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 14187 13454 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 14187 13454 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 14269 13454 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 14269 13454 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 14351 13454 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 14351 13454 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 14433 13454 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 14433 13454 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 14515 13454 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 14515 13454 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 14597 13454 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 14597 13454 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 14678 13454 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 14678 13454 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 14759 13454 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 14759 13454 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 14840 13454 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 14840 13454 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 14921 13454 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 14921 13454 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 15002 13454 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 15002 13454 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 15083 13454 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 15083 13454 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 15164 13454 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 15164 13454 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 15245 13454 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 15245 13454 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 15326 13454 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 15326 13454 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 15407 13454 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 15407 13454 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 15488 13454 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 15488 13454 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 15569 13454 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 15569 13454 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 15650 13454 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 15650 13454 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 15731 13454 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 15731 13454 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 15812 13454 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 15812 13454 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 15893 13454 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 15893 13454 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 15974 13454 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 15974 13454 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 16055 13454 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 16055 13454 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 16136 13454 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 16136 13454 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 16217 13454 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 16217 13454 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 16298 13454 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 16298 13454 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 16379 13454 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 16379 13454 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13390 16460 13454 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13390 16460 13454 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13397 3560 13461 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13397 3560 13461 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13397 3646 13461 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13397 3646 13461 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13397 3732 13461 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13397 3732 13461 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13397 3818 13461 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13397 3818 13461 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13397 3904 13461 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13397 3904 13461 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13397 3990 13461 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13397 3990 13461 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13397 4076 13461 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13397 4076 13461 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13397 4162 13461 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13397 4162 13461 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13397 4248 13461 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13397 4248 13461 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13397 4334 13461 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13397 4334 13461 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13397 4420 13461 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13397 4420 13461 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 16559 13522 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 16559 13522 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 16641 13522 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 16641 13522 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 16723 13522 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 16723 13522 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 16805 13522 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 16805 13522 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 16887 13522 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 16887 13522 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 16969 13522 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 16969 13522 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17051 13522 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17051 13522 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17133 13522 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17133 13522 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17215 13522 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17215 13522 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17297 13522 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17297 13522 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17379 13522 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17379 13522 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17461 13522 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17461 13522 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17543 13522 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17543 13522 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17625 13522 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17625 13522 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17707 13522 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17707 13522 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17789 13522 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17789 13522 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17871 13522 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17871 13522 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17953 13522 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17953 13522 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 18035 13522 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 18035 13522 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 18117 13522 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 18117 13522 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 18199 13522 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 18199 13522 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 18281 13522 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 18281 13522 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 18363 13522 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 18363 13522 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 18445 13522 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 18445 13522 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 18527 13522 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 18527 13522 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 13613 13534 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 13613 13534 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 13695 13534 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 13695 13534 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 13777 13534 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 13777 13534 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 13859 13534 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 13859 13534 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 13941 13534 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 13941 13534 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 14023 13534 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 14023 13534 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 14105 13534 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 14105 13534 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 14187 13534 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 14187 13534 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 14269 13534 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 14269 13534 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 14351 13534 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 14351 13534 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 14433 13534 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 14433 13534 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 14515 13534 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 14515 13534 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 14597 13534 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 14597 13534 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 14678 13534 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 14678 13534 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 14759 13534 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 14759 13534 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 14840 13534 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 14840 13534 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 14921 13534 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 14921 13534 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 15002 13534 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 15002 13534 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 15083 13534 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 15083 13534 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 15164 13534 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 15164 13534 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 15245 13534 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 15245 13534 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 15326 13534 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 15326 13534 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 15407 13534 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 15407 13534 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 15488 13534 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 15488 13534 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 15569 13534 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 15569 13534 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 15650 13534 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 15650 13534 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 15731 13534 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 15731 13534 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 15812 13534 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 15812 13534 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 15893 13534 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 15893 13534 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 15974 13534 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 15974 13534 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 16055 13534 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16055 13534 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 16136 13534 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16136 13534 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 16217 13534 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16217 13534 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 16298 13534 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16298 13534 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 16379 13534 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16379 13534 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13470 16460 13534 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16460 13534 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13478 3560 13542 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13478 3560 13542 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13478 3646 13542 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13478 3646 13542 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13478 3732 13542 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13478 3732 13542 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13478 3818 13542 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13478 3818 13542 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13478 3904 13542 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13478 3904 13542 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13478 3990 13542 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13478 3990 13542 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13478 4076 13542 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13478 4076 13542 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13478 4162 13542 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13478 4162 13542 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13478 4248 13542 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13478 4248 13542 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13478 4334 13542 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13478 4334 13542 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13478 4420 13542 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13478 4420 13542 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 16559 13604 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 16559 13604 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 16641 13604 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 16641 13604 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 16723 13604 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 16723 13604 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 16805 13604 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 16805 13604 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 16887 13604 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 16887 13604 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 16969 13604 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 16969 13604 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17051 13604 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17051 13604 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17133 13604 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17133 13604 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17215 13604 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17215 13604 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17297 13604 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17297 13604 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17379 13604 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17379 13604 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17461 13604 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17461 13604 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17543 13604 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17543 13604 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17625 13604 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17625 13604 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17707 13604 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17707 13604 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17789 13604 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17789 13604 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17871 13604 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17871 13604 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17953 13604 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17953 13604 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 18035 13604 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 18035 13604 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 18117 13604 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 18117 13604 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 18199 13604 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 18199 13604 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 18281 13604 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 18281 13604 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 18363 13604 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 18363 13604 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 18445 13604 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 18445 13604 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 18527 13604 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 18527 13604 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 13613 13614 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 13613 13614 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 13695 13614 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 13695 13614 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 13777 13614 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 13777 13614 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 13859 13614 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 13859 13614 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 13941 13614 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 13941 13614 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 14023 13614 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 14023 13614 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 14105 13614 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 14105 13614 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 14187 13614 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 14187 13614 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 14269 13614 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 14269 13614 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 14351 13614 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 14351 13614 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 14433 13614 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 14433 13614 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 14515 13614 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 14515 13614 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 14597 13614 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 14597 13614 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 14678 13614 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 14678 13614 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 14759 13614 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 14759 13614 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 14840 13614 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 14840 13614 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 14921 13614 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 14921 13614 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 15002 13614 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 15002 13614 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 15083 13614 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 15083 13614 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 15164 13614 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 15164 13614 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 15245 13614 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 15245 13614 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 15326 13614 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 15326 13614 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 15407 13614 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 15407 13614 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 15488 13614 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 15488 13614 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 15569 13614 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 15569 13614 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 15650 13614 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 15650 13614 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 15731 13614 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 15731 13614 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 15812 13614 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 15812 13614 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 15893 13614 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 15893 13614 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 15974 13614 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 15974 13614 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 16055 13614 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 16055 13614 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 16136 13614 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 16136 13614 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 16217 13614 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 16217 13614 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 16298 13614 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 16298 13614 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 16379 13614 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 16379 13614 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13550 16460 13614 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13550 16460 13614 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13559 3560 13623 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13559 3560 13623 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13559 3646 13623 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13559 3646 13623 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13559 3732 13623 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13559 3732 13623 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13559 3818 13623 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13559 3818 13623 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13559 3904 13623 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13559 3904 13623 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13559 3990 13623 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13559 3990 13623 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13559 4076 13623 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13559 4076 13623 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13559 4162 13623 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13559 4162 13623 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13559 4248 13623 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13559 4248 13623 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13559 4334 13623 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13559 4334 13623 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13559 4420 13623 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13559 4420 13623 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 16559 13686 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 16559 13686 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 16641 13686 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 16641 13686 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 16723 13686 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 16723 13686 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 16805 13686 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 16805 13686 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 16887 13686 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 16887 13686 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 16969 13686 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 16969 13686 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17051 13686 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17051 13686 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17133 13686 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17133 13686 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17215 13686 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17215 13686 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17297 13686 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17297 13686 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17379 13686 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17379 13686 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17461 13686 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17461 13686 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17543 13686 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17543 13686 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17625 13686 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17625 13686 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17707 13686 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17707 13686 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17789 13686 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17789 13686 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17871 13686 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17871 13686 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17953 13686 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17953 13686 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 18035 13686 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 18035 13686 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 18117 13686 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 18117 13686 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 18199 13686 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 18199 13686 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 18281 13686 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 18281 13686 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 18363 13686 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 18363 13686 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 18445 13686 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 18445 13686 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 18527 13686 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 18527 13686 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 13613 13694 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 13613 13694 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 13695 13694 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 13695 13694 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 13777 13694 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 13777 13694 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 13859 13694 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 13859 13694 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 13941 13694 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 13941 13694 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 14023 13694 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 14023 13694 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 14105 13694 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 14105 13694 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 14187 13694 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 14187 13694 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 14269 13694 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 14269 13694 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 14351 13694 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 14351 13694 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 14433 13694 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 14433 13694 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 14515 13694 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 14515 13694 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 14597 13694 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 14597 13694 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 14678 13694 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 14678 13694 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 14759 13694 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 14759 13694 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 14840 13694 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 14840 13694 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 14921 13694 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 14921 13694 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 15002 13694 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 15002 13694 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 15083 13694 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 15083 13694 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 15164 13694 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 15164 13694 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 15245 13694 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 15245 13694 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 15326 13694 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 15326 13694 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 15407 13694 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 15407 13694 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 15488 13694 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 15488 13694 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 15569 13694 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 15569 13694 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 15650 13694 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 15650 13694 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 15731 13694 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 15731 13694 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 15812 13694 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 15812 13694 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 15893 13694 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 15893 13694 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 15974 13694 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 15974 13694 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 16055 13694 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 16055 13694 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 16136 13694 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 16136 13694 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 16217 13694 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 16217 13694 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 16298 13694 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 16298 13694 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 16379 13694 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 16379 13694 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13630 16460 13694 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13630 16460 13694 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13640 3560 13704 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13640 3560 13704 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13640 3646 13704 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13640 3646 13704 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13640 3732 13704 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13640 3732 13704 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13640 3818 13704 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13640 3818 13704 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13640 3904 13704 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13640 3904 13704 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13640 3990 13704 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13640 3990 13704 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13640 4076 13704 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13640 4076 13704 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13640 4162 13704 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13640 4162 13704 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13640 4248 13704 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13640 4248 13704 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13640 4334 13704 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13640 4334 13704 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13640 4420 13704 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13640 4420 13704 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 16559 13768 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 16559 13768 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 16641 13768 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 16641 13768 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 16723 13768 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 16723 13768 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 16805 13768 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 16805 13768 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 16887 13768 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 16887 13768 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 16969 13768 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 16969 13768 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17051 13768 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17051 13768 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17133 13768 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17133 13768 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17215 13768 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17215 13768 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17297 13768 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17297 13768 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17379 13768 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17379 13768 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17461 13768 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17461 13768 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17543 13768 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17543 13768 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17625 13768 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17625 13768 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17707 13768 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17707 13768 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17789 13768 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17789 13768 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17871 13768 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17871 13768 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17953 13768 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17953 13768 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 18035 13768 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 18035 13768 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 18117 13768 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 18117 13768 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 18199 13768 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 18199 13768 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 18281 13768 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 18281 13768 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 18363 13768 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 18363 13768 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 18445 13768 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 18445 13768 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 18527 13768 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 18527 13768 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 13613 13774 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 13613 13774 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 13695 13774 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 13695 13774 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 13777 13774 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 13777 13774 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 13859 13774 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 13859 13774 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 13941 13774 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 13941 13774 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 14023 13774 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 14023 13774 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 14105 13774 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 14105 13774 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 14187 13774 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 14187 13774 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 14269 13774 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 14269 13774 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 14351 13774 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 14351 13774 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 14433 13774 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 14433 13774 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 14515 13774 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 14515 13774 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 14597 13774 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 14597 13774 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 14678 13774 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 14678 13774 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 14759 13774 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 14759 13774 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 14840 13774 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 14840 13774 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 14921 13774 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 14921 13774 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 15002 13774 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 15002 13774 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 15083 13774 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 15083 13774 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 15164 13774 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 15164 13774 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 15245 13774 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 15245 13774 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 15326 13774 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 15326 13774 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 15407 13774 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 15407 13774 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 15488 13774 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 15488 13774 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 15569 13774 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 15569 13774 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 15650 13774 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 15650 13774 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 15731 13774 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 15731 13774 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 15812 13774 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 15812 13774 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 15893 13774 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 15893 13774 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 15974 13774 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 15974 13774 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 16055 13774 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 16055 13774 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 16136 13774 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 16136 13774 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 16217 13774 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 16217 13774 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 16298 13774 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 16298 13774 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 16379 13774 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 16379 13774 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13710 16460 13774 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13710 16460 13774 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13721 3560 13785 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13721 3560 13785 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13721 3646 13785 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13721 3646 13785 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13721 3732 13785 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13721 3732 13785 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13721 3818 13785 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13721 3818 13785 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13721 3904 13785 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13721 3904 13785 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13721 3990 13785 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13721 3990 13785 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13721 4076 13785 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13721 4076 13785 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13721 4162 13785 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13721 4162 13785 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13721 4248 13785 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13721 4248 13785 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13721 4334 13785 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13721 4334 13785 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13721 4420 13785 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13721 4420 13785 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 16559 13850 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 16559 13850 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 16641 13850 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 16641 13850 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 16723 13850 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 16723 13850 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 16805 13850 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 16805 13850 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 16887 13850 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 16887 13850 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 16969 13850 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 16969 13850 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17051 13850 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17051 13850 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17133 13850 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17133 13850 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17215 13850 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17215 13850 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17297 13850 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17297 13850 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17379 13850 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17379 13850 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17461 13850 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17461 13850 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17543 13850 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17543 13850 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17625 13850 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17625 13850 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17707 13850 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17707 13850 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17789 13850 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17789 13850 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17871 13850 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17871 13850 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17953 13850 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17953 13850 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 18035 13850 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 18035 13850 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 18117 13850 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 18117 13850 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 18199 13850 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 18199 13850 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 18281 13850 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 18281 13850 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 18363 13850 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 18363 13850 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 18445 13850 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 18445 13850 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 18527 13850 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 18527 13850 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 13613 13854 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 13613 13854 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 13695 13854 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 13695 13854 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 13777 13854 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 13777 13854 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 13859 13854 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 13859 13854 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 13941 13854 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 13941 13854 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 14023 13854 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 14023 13854 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 14105 13854 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 14105 13854 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 14187 13854 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 14187 13854 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 14269 13854 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 14269 13854 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 14351 13854 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 14351 13854 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 14433 13854 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 14433 13854 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 14515 13854 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 14515 13854 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 14597 13854 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 14597 13854 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 14678 13854 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 14678 13854 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 14759 13854 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 14759 13854 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 14840 13854 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 14840 13854 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 14921 13854 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 14921 13854 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 15002 13854 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 15002 13854 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 15083 13854 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 15083 13854 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 15164 13854 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 15164 13854 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 15245 13854 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 15245 13854 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 15326 13854 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 15326 13854 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 15407 13854 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 15407 13854 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 15488 13854 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 15488 13854 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 15569 13854 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 15569 13854 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 15650 13854 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 15650 13854 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 15731 13854 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 15731 13854 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 15812 13854 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 15812 13854 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 15893 13854 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 15893 13854 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 15974 13854 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 15974 13854 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 16055 13854 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 16055 13854 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 16136 13854 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 16136 13854 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 16217 13854 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 16217 13854 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 16298 13854 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 16298 13854 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 16379 13854 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 16379 13854 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13790 16460 13854 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13790 16460 13854 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13802 3560 13866 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 3560 13866 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13802 3646 13866 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 3646 13866 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13802 3732 13866 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 3732 13866 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13802 3818 13866 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 3818 13866 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13802 3904 13866 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 3904 13866 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13802 3990 13866 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 3990 13866 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13802 4076 13866 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 4076 13866 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13802 4162 13866 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 4162 13866 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13802 4248 13866 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 4248 13866 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13802 4334 13866 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 4334 13866 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13802 4420 13866 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 4420 13866 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 16559 13932 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 16559 13932 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 16641 13932 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 16641 13932 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 16723 13932 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 16723 13932 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 16805 13932 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 16805 13932 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 16887 13932 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 16887 13932 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 16969 13932 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 16969 13932 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17051 13932 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17051 13932 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17133 13932 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17133 13932 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17215 13932 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17215 13932 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17297 13932 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17297 13932 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17379 13932 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17379 13932 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17461 13932 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17461 13932 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17543 13932 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17543 13932 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17625 13932 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17625 13932 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17707 13932 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17707 13932 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17789 13932 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17789 13932 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17871 13932 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17871 13932 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17953 13932 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17953 13932 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 18035 13932 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 18035 13932 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 18117 13932 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 18117 13932 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 18199 13932 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 18199 13932 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 18281 13932 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 18281 13932 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 18363 13932 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 18363 13932 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 18445 13932 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 18445 13932 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 18527 13932 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 18527 13932 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 13613 13934 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 13613 13934 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 13695 13934 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 13695 13934 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 13777 13934 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 13777 13934 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 13859 13934 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 13859 13934 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 13941 13934 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 13941 13934 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 14023 13934 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 14023 13934 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 14105 13934 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 14105 13934 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 14187 13934 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 14187 13934 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 14269 13934 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 14269 13934 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 14351 13934 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 14351 13934 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 14433 13934 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 14433 13934 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 14515 13934 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 14515 13934 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 14597 13934 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 14597 13934 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 14678 13934 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 14678 13934 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 14759 13934 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 14759 13934 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 14840 13934 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 14840 13934 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 14921 13934 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 14921 13934 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 15002 13934 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 15002 13934 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 15083 13934 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 15083 13934 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 15164 13934 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 15164 13934 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 15245 13934 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 15245 13934 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 15326 13934 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 15326 13934 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 15407 13934 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 15407 13934 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 15488 13934 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 15488 13934 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 15569 13934 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 15569 13934 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 15650 13934 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 15650 13934 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 15731 13934 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 15731 13934 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 15812 13934 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 15812 13934 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 15893 13934 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 15893 13934 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 15974 13934 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 15974 13934 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 16055 13934 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 16055 13934 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 16136 13934 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 16136 13934 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 16217 13934 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 16217 13934 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 16298 13934 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 16298 13934 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 16379 13934 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 16379 13934 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13870 16460 13934 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13870 16460 13934 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13883 3560 13947 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13883 3560 13947 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13883 3646 13947 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13883 3646 13947 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13883 3732 13947 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13883 3732 13947 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13883 3818 13947 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13883 3818 13947 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13883 3904 13947 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13883 3904 13947 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13883 3990 13947 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13883 3990 13947 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13883 4076 13947 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13883 4076 13947 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13883 4162 13947 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13883 4162 13947 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13883 4248 13947 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13883 4248 13947 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13883 4334 13947 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13883 4334 13947 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13883 4420 13947 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13883 4420 13947 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 13613 14014 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 13613 14014 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 13695 14014 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 13695 14014 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 13777 14014 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 13777 14014 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 13859 14014 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 13859 14014 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 13941 14014 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 13941 14014 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 14023 14014 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 14023 14014 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 14105 14014 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 14105 14014 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 14187 14014 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 14187 14014 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 14269 14014 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 14269 14014 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 14351 14014 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 14351 14014 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 14433 14014 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 14433 14014 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 14515 14014 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 14515 14014 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 14597 14014 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 14597 14014 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 14678 14014 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 14678 14014 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 14759 14014 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 14759 14014 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 14840 14014 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 14840 14014 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 14921 14014 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 14921 14014 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 15002 14014 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 15002 14014 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 15083 14014 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 15083 14014 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 15164 14014 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 15164 14014 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 15245 14014 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 15245 14014 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 15326 14014 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 15326 14014 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 15407 14014 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 15407 14014 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 15488 14014 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 15488 14014 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 15569 14014 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 15569 14014 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 15650 14014 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 15650 14014 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 15731 14014 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 15731 14014 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 15812 14014 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 15812 14014 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 15893 14014 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 15893 14014 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 15974 14014 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 15974 14014 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16055 14014 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16055 14014 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16136 14014 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16136 14014 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16217 14014 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16217 14014 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16298 14014 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16298 14014 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16379 14014 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16379 14014 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16460 14014 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16460 14014 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16559 14014 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16559 14014 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16641 14014 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16641 14014 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16723 14014 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16723 14014 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16805 14014 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16805 14014 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16887 14014 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16887 14014 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16969 14014 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16969 14014 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17051 14014 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17051 14014 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17133 14014 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17133 14014 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17215 14014 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17215 14014 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17297 14014 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17297 14014 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17379 14014 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17379 14014 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17461 14014 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17461 14014 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17543 14014 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17543 14014 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17625 14014 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17625 14014 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17707 14014 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17707 14014 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17789 14014 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17789 14014 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17871 14014 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17871 14014 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17953 14014 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17953 14014 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 18035 14014 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 18035 14014 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 18117 14014 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 18117 14014 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 18199 14014 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 18199 14014 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 18281 14014 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 18281 14014 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 18363 14014 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 18363 14014 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 18445 14014 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 18445 14014 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 18527 14014 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 18527 14014 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13964 3560 14028 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13964 3560 14028 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13964 3646 14028 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13964 3646 14028 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13964 3732 14028 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13964 3732 14028 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13964 3818 14028 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13964 3818 14028 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13964 3904 14028 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13964 3904 14028 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13964 3990 14028 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13964 3990 14028 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13964 4076 14028 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13964 4076 14028 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13964 4162 14028 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13964 4162 14028 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13964 4248 14028 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13964 4248 14028 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13964 4334 14028 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13964 4334 14028 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13964 4420 14028 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13964 4420 14028 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1422 3560 1486 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1422 3560 1486 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1422 3646 1486 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1422 3646 1486 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1422 3732 1486 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1422 3732 1486 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1422 3818 1486 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1422 3818 1486 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1422 3904 1486 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1422 3904 1486 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1422 3990 1486 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1422 3990 1486 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1422 4076 1486 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1422 4076 1486 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1422 4162 1486 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1422 4162 1486 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1422 4248 1486 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1422 4248 1486 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1422 4334 1486 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1422 4334 1486 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1422 4420 1486 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1422 4420 1486 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 13613 1501 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 13613 1501 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 13695 1501 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 13695 1501 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 13777 1501 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 13777 1501 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 13859 1501 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 13859 1501 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 13941 1501 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 13941 1501 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14023 1501 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14023 1501 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14105 1501 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14105 1501 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14187 1501 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14187 1501 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14269 1501 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14269 1501 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14351 1501 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14351 1501 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14433 1501 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14433 1501 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14515 1501 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14515 1501 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14597 1501 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14597 1501 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14678 1501 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14678 1501 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14759 1501 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14759 1501 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14840 1501 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14840 1501 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14921 1501 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14921 1501 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15002 1501 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15002 1501 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15083 1501 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15083 1501 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15164 1501 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15164 1501 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15245 1501 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15245 1501 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15326 1501 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15326 1501 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15407 1501 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15407 1501 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15488 1501 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15488 1501 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15569 1501 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15569 1501 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15650 1501 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15650 1501 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15731 1501 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15731 1501 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15812 1501 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15812 1501 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15893 1501 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15893 1501 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15974 1501 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15974 1501 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 16055 1501 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16055 1501 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 16136 1501 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16136 1501 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 16217 1501 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16217 1501 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 16298 1501 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16298 1501 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 16379 1501 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16379 1501 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 16460 1501 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16460 1501 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 16559 1511 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16559 1511 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 16641 1511 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16641 1511 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 16723 1511 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16723 1511 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 16805 1511 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16805 1511 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 16887 1511 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16887 1511 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 16969 1511 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16969 1511 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17051 1511 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17051 1511 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17133 1511 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17133 1511 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17215 1511 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17215 1511 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17297 1511 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17297 1511 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17379 1511 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17379 1511 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17461 1511 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17461 1511 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17543 1511 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17543 1511 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17625 1511 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17625 1511 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17707 1511 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17707 1511 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17789 1511 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17789 1511 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17871 1511 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17871 1511 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17953 1511 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17953 1511 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 18035 1511 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18035 1511 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 18117 1511 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18117 1511 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 18199 1511 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18199 1511 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 18281 1511 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18281 1511 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 18363 1511 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18363 1511 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 18445 1511 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18445 1511 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 18527 1511 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18527 1511 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1503 3560 1567 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1503 3560 1567 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1503 3646 1567 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1503 3646 1567 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1503 3732 1567 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1503 3732 1567 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1503 3818 1567 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1503 3818 1567 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1503 3904 1567 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1503 3904 1567 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1503 3990 1567 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1503 3990 1567 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1503 4076 1567 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1503 4076 1567 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1503 4162 1567 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1503 4162 1567 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1503 4248 1567 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1503 4248 1567 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1503 4334 1567 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1503 4334 1567 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1503 4420 1567 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1503 4420 1567 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 13613 1581 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 13613 1581 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 13695 1581 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 13695 1581 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 13777 1581 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 13777 1581 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 13859 1581 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 13859 1581 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 13941 1581 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 13941 1581 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14023 1581 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14023 1581 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14105 1581 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14105 1581 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14187 1581 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14187 1581 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14269 1581 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14269 1581 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14351 1581 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14351 1581 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14433 1581 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14433 1581 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14515 1581 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14515 1581 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14597 1581 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14597 1581 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14678 1581 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14678 1581 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14759 1581 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14759 1581 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14840 1581 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14840 1581 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14921 1581 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14921 1581 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15002 1581 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15002 1581 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15083 1581 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15083 1581 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15164 1581 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15164 1581 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15245 1581 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15245 1581 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15326 1581 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15326 1581 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15407 1581 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15407 1581 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15488 1581 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15488 1581 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15569 1581 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15569 1581 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15650 1581 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15650 1581 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15731 1581 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15731 1581 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15812 1581 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15812 1581 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15893 1581 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15893 1581 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15974 1581 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15974 1581 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 16055 1581 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16055 1581 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 16136 1581 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16136 1581 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 16217 1581 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16217 1581 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 16298 1581 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16298 1581 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 16379 1581 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16379 1581 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 16460 1581 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16460 1581 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 16559 1593 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16559 1593 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 16641 1593 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16641 1593 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 16723 1593 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16723 1593 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 16805 1593 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16805 1593 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 16887 1593 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16887 1593 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 16969 1593 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16969 1593 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17051 1593 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17051 1593 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17133 1593 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17133 1593 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17215 1593 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17215 1593 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17297 1593 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17297 1593 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17379 1593 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17379 1593 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17461 1593 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17461 1593 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17543 1593 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17543 1593 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17625 1593 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17625 1593 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17707 1593 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17707 1593 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17789 1593 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17789 1593 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17871 1593 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17871 1593 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17953 1593 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17953 1593 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 18035 1593 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18035 1593 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 18117 1593 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18117 1593 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 18199 1593 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18199 1593 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 18281 1593 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18281 1593 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 18363 1593 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18363 1593 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 18445 1593 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18445 1593 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 18527 1593 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18527 1593 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1584 3560 1648 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1584 3560 1648 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1584 3646 1648 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1584 3646 1648 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1584 3732 1648 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1584 3732 1648 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1584 3818 1648 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1584 3818 1648 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1584 3904 1648 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1584 3904 1648 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1584 3990 1648 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1584 3990 1648 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1584 4076 1648 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1584 4076 1648 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1584 4162 1648 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1584 4162 1648 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1584 4248 1648 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1584 4248 1648 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1584 4334 1648 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1584 4334 1648 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1584 4420 1648 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1584 4420 1648 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 13613 1661 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 13613 1661 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 13695 1661 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 13695 1661 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 13777 1661 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 13777 1661 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 13859 1661 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 13859 1661 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 13941 1661 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 13941 1661 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14023 1661 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14023 1661 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14105 1661 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14105 1661 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14187 1661 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14187 1661 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14269 1661 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14269 1661 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14351 1661 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14351 1661 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14433 1661 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14433 1661 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14515 1661 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14515 1661 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14597 1661 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14597 1661 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14678 1661 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14678 1661 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14759 1661 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14759 1661 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14840 1661 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14840 1661 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14921 1661 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14921 1661 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15002 1661 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15002 1661 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15083 1661 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15083 1661 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15164 1661 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15164 1661 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15245 1661 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15245 1661 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15326 1661 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15326 1661 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15407 1661 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15407 1661 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15488 1661 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15488 1661 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15569 1661 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15569 1661 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15650 1661 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15650 1661 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15731 1661 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15731 1661 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15812 1661 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15812 1661 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15893 1661 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15893 1661 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15974 1661 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15974 1661 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 16055 1661 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16055 1661 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 16136 1661 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16136 1661 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 16217 1661 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16217 1661 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 16298 1661 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16298 1661 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 16379 1661 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16379 1661 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 16460 1661 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16460 1661 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 13613 14094 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 13613 14094 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 13695 14094 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 13695 14094 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 13777 14094 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 13777 14094 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 13859 14094 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 13859 14094 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 13941 14094 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 13941 14094 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 14023 14094 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 14023 14094 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 14105 14094 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 14105 14094 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 14187 14094 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 14187 14094 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 14269 14094 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 14269 14094 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 14351 14094 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 14351 14094 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 14433 14094 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 14433 14094 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 14515 14094 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 14515 14094 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 14597 14094 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 14597 14094 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 14678 14094 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 14678 14094 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 14759 14094 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 14759 14094 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 14840 14094 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 14840 14094 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 14921 14094 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 14921 14094 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 15002 14094 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 15002 14094 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 15083 14094 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 15083 14094 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 15164 14094 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 15164 14094 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 15245 14094 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 15245 14094 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 15326 14094 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 15326 14094 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 15407 14094 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 15407 14094 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 15488 14094 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 15488 14094 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 15569 14094 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 15569 14094 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 15650 14094 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 15650 14094 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 15731 14094 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 15731 14094 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 15812 14094 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 15812 14094 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 15893 14094 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 15893 14094 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 15974 14094 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 15974 14094 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 16055 14094 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 16055 14094 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 16136 14094 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 16136 14094 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 16217 14094 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 16217 14094 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 16298 14094 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 16298 14094 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 16379 14094 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 16379 14094 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14030 16460 14094 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14030 16460 14094 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 16559 14096 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 16559 14096 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 16641 14096 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 16641 14096 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 16723 14096 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 16723 14096 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 16805 14096 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 16805 14096 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 16887 14096 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 16887 14096 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 16969 14096 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 16969 14096 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17051 14096 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17051 14096 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17133 14096 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17133 14096 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17215 14096 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17215 14096 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17297 14096 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17297 14096 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17379 14096 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17379 14096 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17461 14096 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17461 14096 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17543 14096 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17543 14096 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17625 14096 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17625 14096 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17707 14096 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17707 14096 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17789 14096 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17789 14096 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17871 14096 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17871 14096 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17953 14096 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17953 14096 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 18035 14096 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 18035 14096 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 18117 14096 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 18117 14096 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 18199 14096 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 18199 14096 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 18281 14096 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 18281 14096 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 18363 14096 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 18363 14096 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 18445 14096 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 18445 14096 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 18527 14096 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 18527 14096 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14045 3560 14109 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14045 3560 14109 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14045 3646 14109 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14045 3646 14109 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14045 3732 14109 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14045 3732 14109 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14045 3818 14109 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14045 3818 14109 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14045 3904 14109 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14045 3904 14109 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14045 3990 14109 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14045 3990 14109 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14045 4076 14109 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14045 4076 14109 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14045 4162 14109 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14045 4162 14109 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14045 4248 14109 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14045 4248 14109 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14045 4334 14109 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14045 4334 14109 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14045 4420 14109 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14045 4420 14109 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 13613 14174 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 13613 14174 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 13695 14174 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 13695 14174 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 13777 14174 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 13777 14174 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 13859 14174 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 13859 14174 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 13941 14174 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 13941 14174 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 14023 14174 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 14023 14174 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 14105 14174 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 14105 14174 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 14187 14174 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 14187 14174 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 14269 14174 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 14269 14174 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 14351 14174 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 14351 14174 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 14433 14174 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 14433 14174 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 14515 14174 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 14515 14174 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 14597 14174 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 14597 14174 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 14678 14174 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 14678 14174 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 14759 14174 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 14759 14174 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 14840 14174 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 14840 14174 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 14921 14174 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 14921 14174 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 15002 14174 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 15002 14174 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 15083 14174 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 15083 14174 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 15164 14174 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 15164 14174 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 15245 14174 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 15245 14174 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 15326 14174 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 15326 14174 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 15407 14174 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 15407 14174 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 15488 14174 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 15488 14174 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 15569 14174 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 15569 14174 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 15650 14174 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 15650 14174 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 15731 14174 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 15731 14174 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 15812 14174 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 15812 14174 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 15893 14174 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 15893 14174 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 15974 14174 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 15974 14174 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 16055 14174 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 16055 14174 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 16136 14174 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 16136 14174 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 16217 14174 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 16217 14174 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 16298 14174 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 16298 14174 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 16379 14174 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 16379 14174 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14110 16460 14174 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14110 16460 14174 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 16559 14178 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 16559 14178 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 16641 14178 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 16641 14178 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 16723 14178 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 16723 14178 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 16805 14178 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 16805 14178 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 16887 14178 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 16887 14178 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 16969 14178 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 16969 14178 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17051 14178 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17051 14178 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17133 14178 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17133 14178 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17215 14178 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17215 14178 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17297 14178 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17297 14178 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17379 14178 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17379 14178 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17461 14178 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17461 14178 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17543 14178 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17543 14178 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17625 14178 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17625 14178 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17707 14178 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17707 14178 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17789 14178 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17789 14178 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17871 14178 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17871 14178 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17953 14178 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17953 14178 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 18035 14178 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 18035 14178 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 18117 14178 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 18117 14178 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 18199 14178 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 18199 14178 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 18281 14178 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 18281 14178 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 18363 14178 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 18363 14178 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 18445 14178 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 18445 14178 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 18527 14178 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 18527 14178 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14126 3560 14190 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 3560 14190 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14126 3646 14190 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 3646 14190 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14126 3732 14190 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 3732 14190 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14126 3818 14190 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 3818 14190 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14126 3904 14190 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 3904 14190 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14126 3990 14190 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 3990 14190 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14126 4076 14190 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 4076 14190 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14126 4162 14190 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 4162 14190 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14126 4248 14190 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 4248 14190 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14126 4334 14190 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 4334 14190 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14126 4420 14190 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 4420 14190 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 13613 14254 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 13613 14254 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 13695 14254 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 13695 14254 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 13777 14254 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 13777 14254 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 13859 14254 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 13859 14254 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 13941 14254 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 13941 14254 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 14023 14254 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 14023 14254 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 14105 14254 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 14105 14254 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 14187 14254 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 14187 14254 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 14269 14254 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 14269 14254 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 14351 14254 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 14351 14254 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 14433 14254 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 14433 14254 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 14515 14254 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 14515 14254 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 14597 14254 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 14597 14254 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 14678 14254 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 14678 14254 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 14759 14254 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 14759 14254 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 14840 14254 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 14840 14254 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 14921 14254 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 14921 14254 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 15002 14254 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 15002 14254 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 15083 14254 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 15083 14254 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 15164 14254 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 15164 14254 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 15245 14254 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 15245 14254 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 15326 14254 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 15326 14254 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 15407 14254 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 15407 14254 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 15488 14254 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 15488 14254 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 15569 14254 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 15569 14254 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 15650 14254 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 15650 14254 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 15731 14254 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 15731 14254 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 15812 14254 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 15812 14254 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 15893 14254 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 15893 14254 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 15974 14254 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 15974 14254 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 16055 14254 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 16055 14254 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 16136 14254 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 16136 14254 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 16217 14254 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 16217 14254 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 16298 14254 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 16298 14254 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 16379 14254 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 16379 14254 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14190 16460 14254 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14190 16460 14254 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 16559 14260 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 16559 14260 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 16641 14260 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 16641 14260 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 16723 14260 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 16723 14260 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 16805 14260 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 16805 14260 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 16887 14260 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 16887 14260 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 16969 14260 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 16969 14260 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17051 14260 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17051 14260 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17133 14260 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17133 14260 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17215 14260 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17215 14260 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17297 14260 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17297 14260 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17379 14260 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17379 14260 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17461 14260 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17461 14260 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17543 14260 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17543 14260 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17625 14260 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17625 14260 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17707 14260 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17707 14260 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17789 14260 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17789 14260 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17871 14260 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17871 14260 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17953 14260 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17953 14260 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 18035 14260 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 18035 14260 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 18117 14260 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 18117 14260 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 18199 14260 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 18199 14260 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 18281 14260 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 18281 14260 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 18363 14260 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 18363 14260 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 18445 14260 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 18445 14260 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 18527 14260 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 18527 14260 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14207 3560 14271 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14207 3560 14271 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14207 3646 14271 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14207 3646 14271 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14207 3732 14271 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14207 3732 14271 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14207 3818 14271 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14207 3818 14271 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14207 3904 14271 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14207 3904 14271 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14207 3990 14271 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14207 3990 14271 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14207 4076 14271 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14207 4076 14271 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14207 4162 14271 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14207 4162 14271 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14207 4248 14271 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14207 4248 14271 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14207 4334 14271 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14207 4334 14271 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14207 4420 14271 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14207 4420 14271 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 13613 14334 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 13613 14334 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 13695 14334 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 13695 14334 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 13777 14334 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 13777 14334 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 13859 14334 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 13859 14334 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 13941 14334 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 13941 14334 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 14023 14334 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 14023 14334 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 14105 14334 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 14105 14334 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 14187 14334 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 14187 14334 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 14269 14334 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 14269 14334 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 14351 14334 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 14351 14334 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 14433 14334 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 14433 14334 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 14515 14334 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 14515 14334 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 14597 14334 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 14597 14334 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 14678 14334 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 14678 14334 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 14759 14334 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 14759 14334 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 14840 14334 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 14840 14334 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 14921 14334 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 14921 14334 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 15002 14334 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 15002 14334 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 15083 14334 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 15083 14334 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 15164 14334 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 15164 14334 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 15245 14334 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 15245 14334 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 15326 14334 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 15326 14334 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 15407 14334 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 15407 14334 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 15488 14334 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 15488 14334 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 15569 14334 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 15569 14334 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 15650 14334 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 15650 14334 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 15731 14334 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 15731 14334 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 15812 14334 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 15812 14334 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 15893 14334 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 15893 14334 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 15974 14334 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 15974 14334 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 16055 14334 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 16055 14334 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 16136 14334 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 16136 14334 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 16217 14334 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 16217 14334 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 16298 14334 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 16298 14334 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 16379 14334 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 16379 14334 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14270 16460 14334 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14270 16460 14334 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 16559 14342 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 16559 14342 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 16641 14342 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 16641 14342 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 16723 14342 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 16723 14342 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 16805 14342 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 16805 14342 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 16887 14342 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 16887 14342 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 16969 14342 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 16969 14342 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17051 14342 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17051 14342 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17133 14342 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17133 14342 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17215 14342 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17215 14342 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17297 14342 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17297 14342 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17379 14342 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17379 14342 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17461 14342 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17461 14342 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17543 14342 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17543 14342 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17625 14342 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17625 14342 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17707 14342 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17707 14342 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17789 14342 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17789 14342 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17871 14342 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17871 14342 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17953 14342 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17953 14342 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 18035 14342 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 18035 14342 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 18117 14342 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 18117 14342 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 18199 14342 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 18199 14342 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 18281 14342 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 18281 14342 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 18363 14342 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 18363 14342 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 18445 14342 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 18445 14342 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 18527 14342 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 18527 14342 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14288 3560 14352 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14288 3560 14352 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14288 3646 14352 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14288 3646 14352 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14288 3732 14352 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14288 3732 14352 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14288 3818 14352 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14288 3818 14352 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14288 3904 14352 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14288 3904 14352 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14288 3990 14352 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14288 3990 14352 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14288 4076 14352 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14288 4076 14352 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14288 4162 14352 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14288 4162 14352 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14288 4248 14352 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14288 4248 14352 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14288 4334 14352 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14288 4334 14352 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14288 4420 14352 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14288 4420 14352 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 13613 14414 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 13613 14414 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 13695 14414 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 13695 14414 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 13777 14414 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 13777 14414 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 13859 14414 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 13859 14414 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 13941 14414 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 13941 14414 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 14023 14414 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 14023 14414 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 14105 14414 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 14105 14414 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 14187 14414 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 14187 14414 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 14269 14414 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 14269 14414 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 14351 14414 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 14351 14414 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 14433 14414 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 14433 14414 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 14515 14414 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 14515 14414 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 14597 14414 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 14597 14414 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 14678 14414 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 14678 14414 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 14759 14414 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 14759 14414 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 14840 14414 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 14840 14414 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 14921 14414 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 14921 14414 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 15002 14414 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 15002 14414 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 15083 14414 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 15083 14414 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 15164 14414 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 15164 14414 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 15245 14414 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 15245 14414 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 15326 14414 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 15326 14414 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 15407 14414 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 15407 14414 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 15488 14414 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 15488 14414 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 15569 14414 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 15569 14414 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 15650 14414 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 15650 14414 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 15731 14414 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 15731 14414 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 15812 14414 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 15812 14414 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 15893 14414 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 15893 14414 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 15974 14414 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 15974 14414 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 16055 14414 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 16055 14414 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 16136 14414 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 16136 14414 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 16217 14414 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 16217 14414 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 16298 14414 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 16298 14414 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 16379 14414 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 16379 14414 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14350 16460 14414 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14350 16460 14414 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 16559 14424 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 16559 14424 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 16641 14424 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 16641 14424 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 16723 14424 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 16723 14424 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 16805 14424 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 16805 14424 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 16887 14424 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 16887 14424 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 16969 14424 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 16969 14424 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17051 14424 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17051 14424 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17133 14424 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17133 14424 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17215 14424 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17215 14424 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17297 14424 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17297 14424 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17379 14424 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17379 14424 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17461 14424 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17461 14424 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17543 14424 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17543 14424 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17625 14424 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17625 14424 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17707 14424 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17707 14424 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17789 14424 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17789 14424 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17871 14424 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17871 14424 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17953 14424 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17953 14424 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 18035 14424 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 18035 14424 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 18117 14424 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 18117 14424 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 18199 14424 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 18199 14424 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 18281 14424 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 18281 14424 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 18363 14424 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 18363 14424 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 18445 14424 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 18445 14424 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 18527 14424 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 18527 14424 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14369 3560 14433 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14369 3560 14433 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14369 3646 14433 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14369 3646 14433 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14369 3732 14433 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14369 3732 14433 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14369 3818 14433 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14369 3818 14433 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14369 3904 14433 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14369 3904 14433 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14369 3990 14433 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14369 3990 14433 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14369 4076 14433 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14369 4076 14433 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14369 4162 14433 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14369 4162 14433 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14369 4248 14433 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14369 4248 14433 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14369 4334 14433 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14369 4334 14433 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14369 4420 14433 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14369 4420 14433 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 13613 14494 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 13613 14494 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 13695 14494 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 13695 14494 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 13777 14494 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 13777 14494 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 13859 14494 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 13859 14494 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 13941 14494 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 13941 14494 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 14023 14494 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 14023 14494 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 14105 14494 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 14105 14494 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 14187 14494 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 14187 14494 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 14269 14494 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 14269 14494 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 14351 14494 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 14351 14494 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 14433 14494 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 14433 14494 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 14515 14494 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 14515 14494 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 14597 14494 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 14597 14494 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 14678 14494 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 14678 14494 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 14759 14494 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 14759 14494 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 14840 14494 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 14840 14494 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 14921 14494 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 14921 14494 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 15002 14494 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 15002 14494 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 15083 14494 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 15083 14494 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 15164 14494 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 15164 14494 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 15245 14494 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 15245 14494 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 15326 14494 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 15326 14494 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 15407 14494 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 15407 14494 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 15488 14494 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 15488 14494 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 15569 14494 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 15569 14494 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 15650 14494 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 15650 14494 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 15731 14494 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 15731 14494 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 15812 14494 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 15812 14494 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 15893 14494 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 15893 14494 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 15974 14494 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 15974 14494 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 16055 14494 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 16055 14494 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 16136 14494 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 16136 14494 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 16217 14494 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 16217 14494 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 16298 14494 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 16298 14494 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 16379 14494 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 16379 14494 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14430 16460 14494 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14430 16460 14494 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 16559 14506 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16559 14506 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 16641 14506 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16641 14506 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 16723 14506 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16723 14506 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 16805 14506 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16805 14506 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 16887 14506 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16887 14506 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 16969 14506 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16969 14506 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17051 14506 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17051 14506 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17133 14506 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17133 14506 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17215 14506 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17215 14506 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17297 14506 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17297 14506 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17379 14506 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17379 14506 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17461 14506 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17461 14506 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17543 14506 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17543 14506 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17625 14506 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17625 14506 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17707 14506 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17707 14506 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17789 14506 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17789 14506 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17871 14506 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17871 14506 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17953 14506 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17953 14506 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 18035 14506 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 18035 14506 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 18117 14506 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 18117 14506 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 18199 14506 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 18199 14506 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 18281 14506 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 18281 14506 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 18363 14506 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 18363 14506 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 18445 14506 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 18445 14506 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 18527 14506 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 18527 14506 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14451 3560 14515 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14451 3560 14515 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14451 3646 14515 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14451 3646 14515 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14451 3732 14515 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14451 3732 14515 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14451 3818 14515 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14451 3818 14515 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14451 3904 14515 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14451 3904 14515 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14451 3990 14515 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14451 3990 14515 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14451 4076 14515 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14451 4076 14515 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14451 4162 14515 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14451 4162 14515 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14451 4248 14515 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14451 4248 14515 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14451 4334 14515 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14451 4334 14515 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14451 4420 14515 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14451 4420 14515 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 13613 14574 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 13613 14574 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 13695 14574 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 13695 14574 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 13777 14574 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 13777 14574 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 13859 14574 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 13859 14574 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 13941 14574 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 13941 14574 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 14023 14574 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 14023 14574 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 14105 14574 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 14105 14574 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 14187 14574 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 14187 14574 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 14269 14574 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 14269 14574 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 14351 14574 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 14351 14574 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 14433 14574 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 14433 14574 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 14515 14574 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 14515 14574 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 14597 14574 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 14597 14574 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 14678 14574 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 14678 14574 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 14759 14574 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 14759 14574 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 14840 14574 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 14840 14574 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 14921 14574 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 14921 14574 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 15002 14574 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 15002 14574 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 15083 14574 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 15083 14574 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 15164 14574 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 15164 14574 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 15245 14574 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 15245 14574 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 15326 14574 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 15326 14574 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 15407 14574 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 15407 14574 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 15488 14574 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 15488 14574 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 15569 14574 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 15569 14574 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 15650 14574 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 15650 14574 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 15731 14574 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 15731 14574 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 15812 14574 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 15812 14574 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 15893 14574 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 15893 14574 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 15974 14574 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 15974 14574 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 16055 14574 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 16055 14574 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 16136 14574 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 16136 14574 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 16217 14574 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 16217 14574 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 16298 14574 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 16298 14574 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 16379 14574 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 16379 14574 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14510 16460 14574 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14510 16460 14574 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 16559 14588 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 16559 14588 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 16641 14588 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 16641 14588 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 16723 14588 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 16723 14588 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 16805 14588 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 16805 14588 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 16887 14588 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 16887 14588 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 16969 14588 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 16969 14588 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17051 14588 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17051 14588 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17133 14588 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17133 14588 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17215 14588 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17215 14588 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17297 14588 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17297 14588 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17379 14588 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17379 14588 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17461 14588 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17461 14588 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17543 14588 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17543 14588 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17625 14588 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17625 14588 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17707 14588 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17707 14588 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17789 14588 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17789 14588 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17871 14588 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17871 14588 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17953 14588 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17953 14588 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 18035 14588 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 18035 14588 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 18117 14588 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 18117 14588 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 18199 14588 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 18199 14588 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 18281 14588 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 18281 14588 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 18363 14588 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 18363 14588 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 18445 14588 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 18445 14588 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 18527 14588 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 18527 14588 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14533 3560 14597 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14533 3560 14597 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14533 3646 14597 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14533 3646 14597 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14533 3732 14597 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14533 3732 14597 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14533 3818 14597 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14533 3818 14597 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14533 3904 14597 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14533 3904 14597 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14533 3990 14597 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14533 3990 14597 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14533 4076 14597 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14533 4076 14597 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14533 4162 14597 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14533 4162 14597 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14533 4248 14597 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14533 4248 14597 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14533 4334 14597 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14533 4334 14597 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14533 4420 14597 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14533 4420 14597 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 13613 14654 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 13613 14654 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 13695 14654 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 13695 14654 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 13777 14654 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 13777 14654 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 13859 14654 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 13859 14654 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 13941 14654 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 13941 14654 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 14023 14654 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 14023 14654 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 14105 14654 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 14105 14654 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 14187 14654 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 14187 14654 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 14269 14654 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 14269 14654 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 14351 14654 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 14351 14654 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 14433 14654 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 14433 14654 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 14515 14654 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 14515 14654 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 14597 14654 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 14597 14654 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 14678 14654 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 14678 14654 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 14759 14654 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 14759 14654 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 14840 14654 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 14840 14654 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 14921 14654 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 14921 14654 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 15002 14654 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 15002 14654 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 15083 14654 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 15083 14654 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 15164 14654 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 15164 14654 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 15245 14654 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 15245 14654 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 15326 14654 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 15326 14654 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 15407 14654 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 15407 14654 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 15488 14654 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 15488 14654 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 15569 14654 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 15569 14654 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 15650 14654 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 15650 14654 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 15731 14654 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 15731 14654 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 15812 14654 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 15812 14654 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 15893 14654 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 15893 14654 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 15974 14654 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 15974 14654 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 16055 14654 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 16055 14654 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 16136 14654 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 16136 14654 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 16217 14654 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 16217 14654 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 16298 14654 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 16298 14654 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 16379 14654 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 16379 14654 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14590 16460 14654 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14590 16460 14654 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 16559 14670 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 16559 14670 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 16641 14670 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 16641 14670 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 16723 14670 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 16723 14670 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 16805 14670 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 16805 14670 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 16887 14670 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 16887 14670 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 16969 14670 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 16969 14670 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17051 14670 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17051 14670 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17133 14670 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17133 14670 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17215 14670 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17215 14670 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17297 14670 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17297 14670 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17379 14670 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17379 14670 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17461 14670 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17461 14670 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17543 14670 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17543 14670 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17625 14670 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17625 14670 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17707 14670 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17707 14670 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17789 14670 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17789 14670 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17871 14670 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17871 14670 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17953 14670 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17953 14670 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 18035 14670 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 18035 14670 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 18117 14670 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 18117 14670 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 18199 14670 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 18199 14670 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 18281 14670 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 18281 14670 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 18363 14670 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 18363 14670 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 18445 14670 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 18445 14670 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 18527 14670 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 18527 14670 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14615 3560 14679 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14615 3560 14679 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14615 3646 14679 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14615 3646 14679 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14615 3732 14679 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14615 3732 14679 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14615 3818 14679 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14615 3818 14679 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14615 3904 14679 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14615 3904 14679 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14615 3990 14679 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14615 3990 14679 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14615 4076 14679 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14615 4076 14679 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14615 4162 14679 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14615 4162 14679 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14615 4248 14679 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14615 4248 14679 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14615 4334 14679 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14615 4334 14679 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14615 4420 14679 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14615 4420 14679 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 13613 14734 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 13613 14734 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 13695 14734 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 13695 14734 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 13777 14734 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 13777 14734 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 13859 14734 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 13859 14734 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 13941 14734 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 13941 14734 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 14023 14734 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 14023 14734 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 14105 14734 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 14105 14734 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 14187 14734 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 14187 14734 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 14269 14734 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 14269 14734 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 14351 14734 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 14351 14734 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 14433 14734 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 14433 14734 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 14515 14734 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 14515 14734 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 14597 14734 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 14597 14734 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 14678 14734 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 14678 14734 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 14759 14734 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 14759 14734 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 14840 14734 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 14840 14734 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 14921 14734 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 14921 14734 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 15002 14734 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 15002 14734 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 15083 14734 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 15083 14734 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 15164 14734 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 15164 14734 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 15245 14734 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 15245 14734 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 15326 14734 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 15326 14734 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 15407 14734 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 15407 14734 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 15488 14734 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 15488 14734 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 15569 14734 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 15569 14734 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 15650 14734 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 15650 14734 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 15731 14734 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 15731 14734 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 15812 14734 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 15812 14734 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 15893 14734 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 15893 14734 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 15974 14734 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 15974 14734 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 16055 14734 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 16055 14734 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 16136 14734 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 16136 14734 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 16217 14734 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 16217 14734 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 16298 14734 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 16298 14734 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 16379 14734 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 16379 14734 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14670 16460 14734 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14670 16460 14734 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 16559 14752 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 16559 14752 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 16641 14752 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 16641 14752 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 16723 14752 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 16723 14752 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 16805 14752 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 16805 14752 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 16887 14752 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 16887 14752 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 16969 14752 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 16969 14752 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17051 14752 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17051 14752 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17133 14752 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17133 14752 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17215 14752 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17215 14752 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17297 14752 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17297 14752 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17379 14752 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17379 14752 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17461 14752 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17461 14752 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17543 14752 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17543 14752 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17625 14752 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17625 14752 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17707 14752 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17707 14752 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17789 14752 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17789 14752 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17871 14752 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17871 14752 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17953 14752 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17953 14752 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 18035 14752 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 18035 14752 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 18117 14752 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 18117 14752 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 18199 14752 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 18199 14752 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 18281 14752 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 18281 14752 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 18363 14752 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 18363 14752 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 18445 14752 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 18445 14752 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 18527 14752 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 18527 14752 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14697 3560 14761 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14697 3560 14761 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14697 3646 14761 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14697 3646 14761 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14697 3732 14761 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14697 3732 14761 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14697 3818 14761 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14697 3818 14761 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14697 3904 14761 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14697 3904 14761 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14697 3990 14761 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14697 3990 14761 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14697 4076 14761 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14697 4076 14761 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14697 4162 14761 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14697 4162 14761 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14697 4248 14761 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14697 4248 14761 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14697 4334 14761 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14697 4334 14761 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14697 4420 14761 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14697 4420 14761 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 13613 14814 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 13613 14814 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 13695 14814 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 13695 14814 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 13777 14814 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 13777 14814 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 13859 14814 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 13859 14814 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 13941 14814 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 13941 14814 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 14023 14814 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 14023 14814 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 14105 14814 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 14105 14814 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 14187 14814 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 14187 14814 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 14269 14814 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 14269 14814 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 14351 14814 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 14351 14814 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 14433 14814 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 14433 14814 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 14515 14814 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 14515 14814 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 14597 14814 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 14597 14814 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 14678 14814 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 14678 14814 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 14759 14814 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 14759 14814 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 14840 14814 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 14840 14814 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 14921 14814 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 14921 14814 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 15002 14814 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 15002 14814 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 15083 14814 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 15083 14814 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 15164 14814 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 15164 14814 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 15245 14814 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 15245 14814 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 15326 14814 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 15326 14814 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 15407 14814 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 15407 14814 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 15488 14814 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 15488 14814 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 15569 14814 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 15569 14814 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 15650 14814 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 15650 14814 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 15731 14814 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 15731 14814 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 15812 14814 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 15812 14814 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 15893 14814 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 15893 14814 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 15974 14814 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 15974 14814 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 16055 14814 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 16055 14814 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 16136 14814 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 16136 14814 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 16217 14814 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 16217 14814 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 16298 14814 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 16298 14814 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 16379 14814 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 16379 14814 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14750 16460 14814 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14750 16460 14814 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 16559 14834 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 16559 14834 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 16641 14834 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 16641 14834 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 16723 14834 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 16723 14834 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 16805 14834 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 16805 14834 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 16887 14834 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 16887 14834 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 16969 14834 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 16969 14834 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 17051 14834 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17051 14834 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 17133 14834 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17133 14834 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 17215 14834 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17215 14834 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 17297 14834 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17297 14834 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 17379 14834 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17379 14834 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 17461 14834 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17461 14834 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 17543 14834 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17543 14834 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 17625 14834 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17625 14834 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 17707 14834 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17707 14834 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 17789 14834 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17789 14834 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 17871 14834 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17871 14834 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 17953 14834 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17953 14834 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 18035 14834 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 18035 14834 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 18117 14834 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 18117 14834 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 18199 14834 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 18199 14834 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 18281 14834 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 18281 14834 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 18363 14834 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 18363 14834 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 18445 14834 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 18445 14834 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14770 18527 14834 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 18527 14834 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14779 3560 14843 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14779 3560 14843 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14779 3646 14843 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14779 3646 14843 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14779 3732 14843 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14779 3732 14843 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14779 3818 14843 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14779 3818 14843 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14779 3904 14843 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14779 3904 14843 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14779 3990 14843 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14779 3990 14843 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14779 4076 14843 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14779 4076 14843 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14779 4162 14843 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14779 4162 14843 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14779 4248 14843 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14779 4248 14843 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14779 4334 14843 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14779 4334 14843 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14779 4420 14843 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14779 4420 14843 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 13613 14894 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 13613 14894 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 13695 14894 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 13695 14894 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 13777 14894 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 13777 14894 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 13859 14894 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 13859 14894 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 13941 14894 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 13941 14894 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 14023 14894 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 14023 14894 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 14105 14894 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 14105 14894 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 14187 14894 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 14187 14894 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 14269 14894 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 14269 14894 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 14351 14894 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 14351 14894 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 14433 14894 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 14433 14894 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 14515 14894 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 14515 14894 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 14597 14894 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 14597 14894 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 14678 14894 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 14678 14894 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 14759 14894 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 14759 14894 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 14840 14894 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 14840 14894 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 14921 14894 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 14921 14894 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 15002 14894 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 15002 14894 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 15083 14894 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 15083 14894 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 15164 14894 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 15164 14894 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 15245 14894 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 15245 14894 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 15326 14894 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 15326 14894 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 15407 14894 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 15407 14894 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 15488 14894 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 15488 14894 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 15569 14894 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 15569 14894 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 15650 14894 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 15650 14894 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 15731 14894 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 15731 14894 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 15812 14894 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 15812 14894 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 15893 14894 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 15893 14894 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 15974 14894 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 15974 14894 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 16055 14894 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 16055 14894 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 16136 14894 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 16136 14894 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 16217 14894 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 16217 14894 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 16298 14894 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 16298 14894 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 16379 14894 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 16379 14894 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14830 16460 14894 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14830 16460 14894 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 16559 14916 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 16559 14916 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 16641 14916 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 16641 14916 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 16723 14916 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 16723 14916 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 16805 14916 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 16805 14916 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 16887 14916 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 16887 14916 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 16969 14916 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 16969 14916 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 17051 14916 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17051 14916 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 17133 14916 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17133 14916 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 17215 14916 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17215 14916 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 17297 14916 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17297 14916 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 17379 14916 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17379 14916 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 17461 14916 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17461 14916 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 17543 14916 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17543 14916 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 17625 14916 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17625 14916 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 17707 14916 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17707 14916 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 17789 14916 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17789 14916 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 17871 14916 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17871 14916 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 17953 14916 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17953 14916 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 18035 14916 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 18035 14916 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 18117 14916 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 18117 14916 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 18199 14916 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 18199 14916 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 18281 14916 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 18281 14916 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 18363 14916 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 18363 14916 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 18445 14916 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 18445 14916 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14852 18527 14916 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 18527 14916 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14861 3560 14925 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14861 3560 14925 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14861 3646 14925 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14861 3646 14925 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14861 3732 14925 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14861 3732 14925 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14861 3818 14925 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14861 3818 14925 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14861 3904 14925 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14861 3904 14925 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14861 3990 14925 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14861 3990 14925 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14861 4076 14925 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14861 4076 14925 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14861 4162 14925 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14861 4162 14925 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14861 4248 14925 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14861 4248 14925 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14861 4334 14925 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14861 4334 14925 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14861 4420 14925 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14861 4420 14925 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 16559 1675 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16559 1675 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 16641 1675 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16641 1675 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 16723 1675 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16723 1675 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 16805 1675 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16805 1675 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 16887 1675 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16887 1675 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 16969 1675 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16969 1675 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17051 1675 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17051 1675 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17133 1675 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17133 1675 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17215 1675 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17215 1675 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17297 1675 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17297 1675 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17379 1675 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17379 1675 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17461 1675 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17461 1675 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17543 1675 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17543 1675 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17625 1675 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17625 1675 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17707 1675 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17707 1675 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17789 1675 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17789 1675 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17871 1675 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17871 1675 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17953 1675 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17953 1675 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 18035 1675 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18035 1675 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 18117 1675 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18117 1675 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 18199 1675 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18199 1675 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 18281 1675 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18281 1675 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 18363 1675 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18363 1675 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 18445 1675 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18445 1675 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 18527 1675 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18527 1675 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1665 3560 1729 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1665 3560 1729 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1665 3646 1729 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1665 3646 1729 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1665 3732 1729 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1665 3732 1729 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1665 3818 1729 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1665 3818 1729 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1665 3904 1729 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1665 3904 1729 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1665 3990 1729 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1665 3990 1729 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1665 4076 1729 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1665 4076 1729 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1665 4162 1729 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1665 4162 1729 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1665 4248 1729 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1665 4248 1729 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1665 4334 1729 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1665 4334 1729 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1665 4420 1729 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1665 4420 1729 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 13613 1741 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 13613 1741 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 13695 1741 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 13695 1741 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 13777 1741 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 13777 1741 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 13859 1741 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 13859 1741 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 13941 1741 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 13941 1741 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14023 1741 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14023 1741 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14105 1741 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14105 1741 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14187 1741 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14187 1741 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14269 1741 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14269 1741 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14351 1741 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14351 1741 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14433 1741 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14433 1741 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14515 1741 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14515 1741 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14597 1741 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14597 1741 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14678 1741 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14678 1741 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14759 1741 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14759 1741 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14840 1741 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14840 1741 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14921 1741 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14921 1741 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15002 1741 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15002 1741 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15083 1741 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15083 1741 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15164 1741 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15164 1741 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15245 1741 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15245 1741 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15326 1741 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15326 1741 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15407 1741 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15407 1741 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15488 1741 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15488 1741 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15569 1741 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15569 1741 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15650 1741 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15650 1741 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15731 1741 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15731 1741 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15812 1741 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15812 1741 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15893 1741 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15893 1741 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15974 1741 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15974 1741 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 16055 1741 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16055 1741 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 16136 1741 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16136 1741 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 16217 1741 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16217 1741 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 16298 1741 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16298 1741 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 16379 1741 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16379 1741 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 16460 1741 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16460 1741 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 16559 1757 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16559 1757 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 16641 1757 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16641 1757 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 16723 1757 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16723 1757 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 16805 1757 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16805 1757 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 16887 1757 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16887 1757 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 16969 1757 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16969 1757 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17051 1757 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17051 1757 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17133 1757 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17133 1757 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17215 1757 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17215 1757 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17297 1757 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17297 1757 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17379 1757 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17379 1757 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17461 1757 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17461 1757 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17543 1757 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17543 1757 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17625 1757 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17625 1757 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17707 1757 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17707 1757 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17789 1757 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17789 1757 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17871 1757 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17871 1757 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17953 1757 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17953 1757 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 18035 1757 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18035 1757 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 18117 1757 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18117 1757 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 18199 1757 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18199 1757 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 18281 1757 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18281 1757 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 18363 1757 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18363 1757 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 18445 1757 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18445 1757 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 18527 1757 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18527 1757 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1746 3560 1810 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1746 3560 1810 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1746 3646 1810 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1746 3646 1810 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1746 3732 1810 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1746 3732 1810 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1746 3818 1810 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1746 3818 1810 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1746 3904 1810 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1746 3904 1810 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1746 3990 1810 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1746 3990 1810 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1746 4076 1810 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1746 4076 1810 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1746 4162 1810 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1746 4162 1810 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1746 4248 1810 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1746 4248 1810 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1746 4334 1810 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1746 4334 1810 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1746 4420 1810 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1746 4420 1810 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 13613 1821 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 13613 1821 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 13695 1821 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 13695 1821 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 13777 1821 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 13777 1821 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 13859 1821 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 13859 1821 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 13941 1821 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 13941 1821 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14023 1821 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14023 1821 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14105 1821 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14105 1821 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14187 1821 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14187 1821 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14269 1821 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14269 1821 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14351 1821 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14351 1821 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14433 1821 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14433 1821 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14515 1821 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14515 1821 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14597 1821 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14597 1821 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14678 1821 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14678 1821 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14759 1821 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14759 1821 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14840 1821 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14840 1821 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14921 1821 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14921 1821 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15002 1821 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15002 1821 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15083 1821 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15083 1821 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15164 1821 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15164 1821 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15245 1821 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15245 1821 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15326 1821 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15326 1821 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15407 1821 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15407 1821 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15488 1821 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15488 1821 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15569 1821 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15569 1821 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15650 1821 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15650 1821 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15731 1821 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15731 1821 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15812 1821 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15812 1821 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15893 1821 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15893 1821 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15974 1821 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15974 1821 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 16055 1821 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16055 1821 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 16136 1821 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16136 1821 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 16217 1821 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16217 1821 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 16298 1821 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16298 1821 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 16379 1821 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16379 1821 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 16460 1821 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16460 1821 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 16559 1839 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16559 1839 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 16641 1839 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16641 1839 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 16723 1839 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16723 1839 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 16805 1839 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16805 1839 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 16887 1839 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16887 1839 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 16969 1839 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16969 1839 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17051 1839 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17051 1839 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17133 1839 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17133 1839 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17215 1839 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17215 1839 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17297 1839 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17297 1839 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17379 1839 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17379 1839 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17461 1839 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17461 1839 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17543 1839 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17543 1839 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17625 1839 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17625 1839 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17707 1839 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17707 1839 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17789 1839 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17789 1839 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17871 1839 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17871 1839 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17953 1839 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17953 1839 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 18035 1839 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18035 1839 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 18117 1839 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18117 1839 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 18199 1839 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18199 1839 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 18281 1839 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18281 1839 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 18363 1839 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18363 1839 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 18445 1839 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18445 1839 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 18527 1839 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18527 1839 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1827 3560 1891 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1827 3560 1891 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1827 3646 1891 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1827 3646 1891 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1827 3732 1891 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1827 3732 1891 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1827 3818 1891 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1827 3818 1891 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1827 3904 1891 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1827 3904 1891 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1827 3990 1891 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1827 3990 1891 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1827 4076 1891 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1827 4076 1891 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1827 4162 1891 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1827 4162 1891 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1827 4248 1891 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1827 4248 1891 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1827 4334 1891 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1827 4334 1891 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1827 4420 1891 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1827 4420 1891 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 13613 1901 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 13613 1901 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 13695 1901 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 13695 1901 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 13777 1901 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 13777 1901 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 13859 1901 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 13859 1901 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 13941 1901 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 13941 1901 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14023 1901 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14023 1901 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14105 1901 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14105 1901 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14187 1901 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14187 1901 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14269 1901 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14269 1901 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14351 1901 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14351 1901 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14433 1901 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14433 1901 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14515 1901 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14515 1901 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14597 1901 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14597 1901 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14678 1901 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14678 1901 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14759 1901 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14759 1901 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14840 1901 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14840 1901 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14921 1901 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14921 1901 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15002 1901 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15002 1901 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15083 1901 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15083 1901 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15164 1901 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15164 1901 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15245 1901 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15245 1901 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15326 1901 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15326 1901 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15407 1901 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15407 1901 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15488 1901 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15488 1901 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15569 1901 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15569 1901 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15650 1901 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15650 1901 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15731 1901 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15731 1901 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15812 1901 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15812 1901 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15893 1901 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15893 1901 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15974 1901 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15974 1901 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 16055 1901 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16055 1901 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 16136 1901 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16136 1901 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 16217 1901 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16217 1901 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 16298 1901 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16298 1901 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 16379 1901 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16379 1901 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 16460 1901 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16460 1901 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 16559 1921 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16559 1921 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 16641 1921 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16641 1921 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 16723 1921 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16723 1921 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 16805 1921 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16805 1921 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 16887 1921 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16887 1921 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 16969 1921 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16969 1921 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17051 1921 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17051 1921 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17133 1921 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17133 1921 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17215 1921 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17215 1921 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17297 1921 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17297 1921 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17379 1921 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17379 1921 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17461 1921 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17461 1921 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17543 1921 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17543 1921 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17625 1921 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17625 1921 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17707 1921 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17707 1921 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17789 1921 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17789 1921 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17871 1921 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17871 1921 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17953 1921 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17953 1921 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 18035 1921 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18035 1921 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 18117 1921 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18117 1921 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 18199 1921 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18199 1921 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 18281 1921 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18281 1921 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 18363 1921 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18363 1921 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 18445 1921 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18445 1921 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 18527 1921 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18527 1921 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1908 3560 1972 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1908 3560 1972 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1908 3646 1972 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1908 3646 1972 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1908 3732 1972 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1908 3732 1972 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1908 3818 1972 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1908 3818 1972 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1908 3904 1972 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1908 3904 1972 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1908 3990 1972 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1908 3990 1972 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1908 4076 1972 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1908 4076 1972 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1908 4162 1972 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1908 4162 1972 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1908 4248 1972 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1908 4248 1972 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1908 4334 1972 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1908 4334 1972 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1908 4420 1972 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1908 4420 1972 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 13613 1981 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 13613 1981 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 13695 1981 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 13695 1981 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 13777 1981 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 13777 1981 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 13859 1981 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 13859 1981 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 13941 1981 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 13941 1981 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14023 1981 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14023 1981 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14105 1981 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14105 1981 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14187 1981 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14187 1981 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14269 1981 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14269 1981 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14351 1981 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14351 1981 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14433 1981 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14433 1981 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14515 1981 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14515 1981 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14597 1981 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14597 1981 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14678 1981 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14678 1981 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14759 1981 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14759 1981 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14840 1981 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14840 1981 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14921 1981 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14921 1981 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15002 1981 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15002 1981 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15083 1981 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15083 1981 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15164 1981 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15164 1981 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15245 1981 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15245 1981 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15326 1981 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15326 1981 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15407 1981 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15407 1981 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15488 1981 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15488 1981 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15569 1981 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15569 1981 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15650 1981 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15650 1981 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15731 1981 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15731 1981 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15812 1981 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15812 1981 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15893 1981 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15893 1981 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15974 1981 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15974 1981 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 16055 1981 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16055 1981 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 16136 1981 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16136 1981 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 16217 1981 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16217 1981 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 16298 1981 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16298 1981 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 16379 1981 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16379 1981 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 16460 1981 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16460 1981 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 16559 2003 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16559 2003 16623 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 16641 2003 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16641 2003 16705 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 16723 2003 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16723 2003 16787 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 16805 2003 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16805 2003 16869 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 16887 2003 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16887 2003 16951 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 16969 2003 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16969 2003 17033 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17051 2003 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17051 2003 17115 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17133 2003 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17133 2003 17197 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17215 2003 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17215 2003 17279 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17297 2003 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17297 2003 17361 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17379 2003 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17379 2003 17443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17461 2003 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17461 2003 17525 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17543 2003 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17543 2003 17607 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17625 2003 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17625 2003 17689 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17707 2003 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17707 2003 17771 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17789 2003 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17789 2003 17853 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17871 2003 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17871 2003 17935 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17953 2003 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17953 2003 18017 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 18035 2003 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18035 2003 18099 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 18117 2003 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18117 2003 18181 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 18199 2003 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18199 2003 18263 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 18281 2003 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18281 2003 18345 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 18363 2003 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18363 2003 18427 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 18445 2003 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18445 2003 18509 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 18527 2003 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18527 2003 18591 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1989 3560 2053 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1989 3560 2053 3624 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1989 3646 2053 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1989 3646 2053 3710 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1989 3732 2053 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1989 3732 2053 3796 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1989 3818 2053 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1989 3818 2053 3882 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1989 3904 2053 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1989 3904 2053 3968 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1989 3990 2053 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1989 3990 2053 4054 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1989 4076 2053 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1989 4076 2053 4140 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1989 4162 2053 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1989 4162 2053 4226 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1989 4248 2053 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1989 4248 2053 4312 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1989 4334 2053 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1989 4334 2053 4398 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1989 4420 2053 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1989 4420 2053 4484 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 13613 2061 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 13613 2061 13677 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 13695 2061 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 13695 2061 13759 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 13777 2061 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 13777 2061 13841 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 13859 2061 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 13859 2061 13923 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 13941 2061 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 13941 2061 14005 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14023 2061 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14023 2061 14087 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14105 2061 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14105 2061 14169 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14187 2061 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14187 2061 14251 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14269 2061 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14269 2061 14333 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14351 2061 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14351 2061 14415 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14433 2061 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14433 2061 14497 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14515 2061 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14515 2061 14579 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14597 2061 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14597 2061 14661 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14678 2061 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14678 2061 14742 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14759 2061 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14759 2061 14823 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14840 2061 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14840 2061 14904 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14921 2061 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14921 2061 14985 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15002 2061 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15002 2061 15066 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15083 2061 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15083 2061 15147 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15164 2061 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15164 2061 15228 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15245 2061 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15245 2061 15309 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15326 2061 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15326 2061 15390 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15407 2061 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15407 2061 15471 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15488 2061 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15488 2061 15552 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15569 2061 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15569 2061 15633 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15650 2061 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15650 2061 15714 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15731 2061 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15731 2061 15795 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15812 2061 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15812 2061 15876 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15893 2061 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15893 2061 15957 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15974 2061 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15974 2061 16038 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 16055 2061 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16055 2061 16119 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 16136 2061 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16136 2061 16200 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 16217 2061 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16217 2061 16281 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 16298 2061 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16298 2061 16362 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 16379 2061 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16379 2061 16443 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 16460 2061 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16460 2061 16524 1 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 126 12502 190 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12502 190 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 126 12584 190 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12584 190 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 126 12666 190 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12666 190 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 126 12748 190 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12748 190 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 126 12830 190 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12830 190 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 126 12912 190 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12912 190 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 126 12994 190 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12994 190 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 126 13076 190 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 13076 190 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 126 13158 190 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 13158 190 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 126 13240 190 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 13240 190 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 207 12420 271 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12420 271 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 207 12502 271 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12502 271 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 207 12584 271 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12584 271 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 207 12666 271 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12666 271 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 207 12748 271 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12748 271 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 207 12830 271 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12830 271 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 207 12912 271 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12912 271 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 207 12994 271 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12994 271 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 207 13076 271 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 13076 271 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 207 13158 271 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 13158 271 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 207 13240 271 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 13240 271 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 12420 352 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12420 352 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 12502 352 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12502 352 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 12584 352 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12584 352 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 12666 352 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12666 352 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 12748 352 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12748 352 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 12830 352 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12830 352 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 12912 352 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12912 352 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 12994 352 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12994 352 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 13076 352 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 13076 352 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 13158 352 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 13158 352 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 13240 352 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 13240 352 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 12420 433 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12420 433 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 12502 433 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12502 433 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 12584 433 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12584 433 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 12666 433 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12666 433 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 12748 433 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12748 433 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 12830 433 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12830 433 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 12912 433 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12912 433 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 12994 433 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12994 433 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 13076 433 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 13076 433 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 13158 433 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 13158 433 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 13240 433 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 13240 433 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 12420 2134 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12420 2134 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 12502 2134 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12502 2134 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 12584 2134 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12584 2134 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 12666 2134 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12666 2134 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 12748 2134 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12748 2134 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 12830 2134 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12830 2134 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 12912 2134 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12912 2134 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 12994 2134 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12994 2134 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 13076 2134 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 13076 2134 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 13158 2134 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 13158 2134 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 13240 2134 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 13240 2134 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 12420 2215 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12420 2215 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 12502 2215 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12502 2215 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 12584 2215 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12584 2215 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 12666 2215 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12666 2215 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 12748 2215 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12748 2215 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 12830 2215 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12830 2215 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 12912 2215 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12912 2215 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 12994 2215 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12994 2215 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 13076 2215 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 13076 2215 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 13158 2215 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 13158 2215 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 13240 2215 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 13240 2215 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 12420 2296 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12420 2296 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 12502 2296 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12502 2296 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 12584 2296 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12584 2296 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 12666 2296 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12666 2296 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 12748 2296 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12748 2296 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 12830 2296 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12830 2296 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 12912 2296 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12912 2296 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 12994 2296 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12994 2296 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 13076 2296 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 13076 2296 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 13158 2296 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 13158 2296 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 13240 2296 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 13240 2296 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 12420 2377 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12420 2377 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 12502 2377 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12502 2377 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 12584 2377 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12584 2377 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 12666 2377 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12666 2377 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 12748 2377 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12748 2377 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 12830 2377 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12830 2377 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 12912 2377 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12912 2377 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 12994 2377 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12994 2377 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 13076 2377 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 13076 2377 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 13158 2377 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 13158 2377 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 13240 2377 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 13240 2377 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 12420 2458 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12420 2458 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 12502 2458 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12502 2458 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 12584 2458 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12584 2458 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 12666 2458 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12666 2458 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 12748 2458 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12748 2458 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 12830 2458 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12830 2458 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 12912 2458 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12912 2458 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 12994 2458 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12994 2458 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 13076 2458 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 13076 2458 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 13158 2458 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 13158 2458 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 13240 2458 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 13240 2458 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 12420 2539 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12420 2539 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 12502 2539 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12502 2539 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 12584 2539 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12584 2539 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 12666 2539 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12666 2539 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 12748 2539 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12748 2539 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 12830 2539 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12830 2539 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 12912 2539 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12912 2539 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 12994 2539 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12994 2539 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 13076 2539 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 13076 2539 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 13158 2539 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 13158 2539 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 13240 2539 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 13240 2539 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 12420 2620 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12420 2620 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 12502 2620 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12502 2620 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 12584 2620 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12584 2620 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 12666 2620 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12666 2620 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 12748 2620 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12748 2620 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 12830 2620 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12830 2620 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 12912 2620 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12912 2620 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 12994 2620 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12994 2620 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 13076 2620 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 13076 2620 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 13158 2620 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 13158 2620 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 13240 2620 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 13240 2620 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 12420 2701 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12420 2701 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 12502 2701 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12502 2701 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 12584 2701 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12584 2701 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 12666 2701 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12666 2701 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 12748 2701 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12748 2701 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 12830 2701 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12830 2701 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 12912 2701 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12912 2701 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 12994 2701 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12994 2701 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 13076 2701 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 13076 2701 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 13158 2701 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 13158 2701 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 13240 2701 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 13240 2701 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 12420 2782 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12420 2782 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 12502 2782 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12502 2782 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 12584 2782 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12584 2782 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 12666 2782 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12666 2782 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 12748 2782 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12748 2782 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 12830 2782 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12830 2782 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 12912 2782 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12912 2782 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 12994 2782 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12994 2782 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 13076 2782 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 13076 2782 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 13158 2782 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 13158 2782 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 13240 2782 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 13240 2782 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 12420 2863 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12420 2863 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 12502 2863 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12502 2863 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 12584 2863 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12584 2863 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 12666 2863 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12666 2863 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 12748 2863 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12748 2863 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 12830 2863 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12830 2863 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 12912 2863 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12912 2863 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 12994 2863 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12994 2863 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 13076 2863 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 13076 2863 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 13158 2863 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 13158 2863 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 13240 2863 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 13240 2863 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 12420 2944 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12420 2944 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 12502 2944 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12502 2944 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 12584 2944 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12584 2944 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 12666 2944 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12666 2944 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 12748 2944 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12748 2944 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 12830 2944 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12830 2944 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 12912 2944 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12912 2944 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 12994 2944 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12994 2944 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 13076 2944 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 13076 2944 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 13158 2944 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 13158 2944 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 13240 2944 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 13240 2944 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 12420 3025 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12420 3025 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 12502 3025 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12502 3025 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 12584 3025 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12584 3025 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 12666 3025 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12666 3025 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 12748 3025 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12748 3025 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 12830 3025 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12830 3025 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 12912 3025 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12912 3025 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 12994 3025 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12994 3025 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 13076 3025 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 13076 3025 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 13158 3025 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 13158 3025 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 13240 3025 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 13240 3025 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 12420 3106 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12420 3106 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 12502 3106 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12502 3106 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 12584 3106 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12584 3106 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 12666 3106 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12666 3106 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 12748 3106 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12748 3106 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 12830 3106 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12830 3106 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 12912 3106 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12912 3106 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 12994 3106 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12994 3106 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 13076 3106 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 13076 3106 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 13158 3106 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 13158 3106 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 13240 3106 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 13240 3106 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 12420 3187 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12420 3187 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 12502 3187 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12502 3187 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 12584 3187 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12584 3187 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 12666 3187 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12666 3187 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 12748 3187 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12748 3187 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 12830 3187 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12830 3187 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 12912 3187 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12912 3187 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 12994 3187 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12994 3187 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 13076 3187 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 13076 3187 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 13158 3187 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 13158 3187 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 13240 3187 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 13240 3187 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 12420 3268 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12420 3268 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 12502 3268 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12502 3268 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 12584 3268 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12584 3268 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 12666 3268 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12666 3268 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 12748 3268 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12748 3268 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 12830 3268 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12830 3268 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 12912 3268 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12912 3268 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 12994 3268 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12994 3268 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 13076 3268 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 13076 3268 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 13158 3268 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 13158 3268 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 13240 3268 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 13240 3268 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 12420 3349 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12420 3349 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 12502 3349 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12502 3349 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 12584 3349 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12584 3349 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 12666 3349 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12666 3349 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 12748 3349 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12748 3349 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 12830 3349 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12830 3349 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 12912 3349 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12912 3349 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 12994 3349 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12994 3349 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 13076 3349 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 13076 3349 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 13158 3349 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 13158 3349 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 13240 3349 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 13240 3349 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 12420 3430 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12420 3430 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 12502 3430 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12502 3430 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 12584 3430 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12584 3430 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 12666 3430 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12666 3430 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 12748 3430 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12748 3430 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 12830 3430 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12830 3430 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 12912 3430 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12912 3430 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 12994 3430 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12994 3430 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 13076 3430 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 13076 3430 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 13158 3430 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 13158 3430 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 13240 3430 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 13240 3430 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 12420 3511 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12420 3511 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 12502 3511 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12502 3511 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 12584 3511 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12584 3511 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 12666 3511 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12666 3511 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 12748 3511 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12748 3511 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 12830 3511 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12830 3511 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 12912 3511 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12912 3511 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 12994 3511 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12994 3511 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 13076 3511 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 13076 3511 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 13158 3511 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 13158 3511 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 13240 3511 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 13240 3511 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 12420 3592 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12420 3592 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 12502 3592 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12502 3592 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 12584 3592 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12584 3592 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 12666 3592 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12666 3592 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 12748 3592 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12748 3592 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 12830 3592 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12830 3592 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 12912 3592 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12912 3592 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 12994 3592 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12994 3592 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 13076 3592 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 13076 3592 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 13158 3592 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 13158 3592 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 13240 3592 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 13240 3592 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 12420 3673 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12420 3673 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 12502 3673 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12502 3673 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 12584 3673 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12584 3673 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 12666 3673 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12666 3673 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 12748 3673 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12748 3673 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 12830 3673 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12830 3673 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 12912 3673 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12912 3673 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 12994 3673 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12994 3673 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 13076 3673 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 13076 3673 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 13158 3673 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 13158 3673 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 13240 3673 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 13240 3673 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 12420 3754 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12420 3754 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 12502 3754 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12502 3754 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 12584 3754 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12584 3754 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 12666 3754 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12666 3754 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 12748 3754 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12748 3754 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 12830 3754 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12830 3754 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 12912 3754 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12912 3754 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 12994 3754 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12994 3754 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 13076 3754 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 13076 3754 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 13158 3754 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 13158 3754 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 13240 3754 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 13240 3754 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 12420 3835 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12420 3835 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 12502 3835 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12502 3835 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 12584 3835 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12584 3835 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 12666 3835 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12666 3835 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 12748 3835 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12748 3835 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 12830 3835 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12830 3835 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 12912 3835 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12912 3835 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 12994 3835 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12994 3835 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 13076 3835 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 13076 3835 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 13158 3835 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 13158 3835 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 13240 3835 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 13240 3835 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 12420 3916 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12420 3916 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 12502 3916 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12502 3916 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 12584 3916 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12584 3916 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 12666 3916 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12666 3916 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 12748 3916 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12748 3916 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 12830 3916 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12830 3916 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 12912 3916 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12912 3916 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 12994 3916 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12994 3916 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 13076 3916 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 13076 3916 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 13158 3916 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 13158 3916 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 13240 3916 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 13240 3916 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 12420 3997 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12420 3997 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 12502 3997 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12502 3997 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 12584 3997 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12584 3997 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 12666 3997 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12666 3997 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 12748 3997 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12748 3997 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 12830 3997 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12830 3997 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 12912 3997 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12912 3997 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 12994 3997 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12994 3997 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 13076 3997 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 13076 3997 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 13158 3997 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 13158 3997 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 13240 3997 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 13240 3997 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 12420 514 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12420 514 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 12502 514 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12502 514 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 12584 514 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12584 514 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 12666 514 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12666 514 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 12748 514 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12748 514 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 12830 514 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12830 514 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 12912 514 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12912 514 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 12994 514 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12994 514 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 13076 514 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 13076 514 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 13158 514 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 13158 514 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 13240 514 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 13240 514 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 12420 595 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12420 595 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 12502 595 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12502 595 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 12584 595 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12584 595 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 12666 595 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12666 595 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 12748 595 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12748 595 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 12830 595 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12830 595 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 12912 595 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12912 595 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 12994 595 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12994 595 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 13076 595 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 13076 595 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 13158 595 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 13158 595 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 13240 595 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 13240 595 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 12420 4078 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12420 4078 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 12502 4078 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12502 4078 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 12584 4078 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12584 4078 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 12666 4078 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12666 4078 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 12748 4078 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12748 4078 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 12830 4078 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12830 4078 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 12912 4078 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12912 4078 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 12994 4078 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12994 4078 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 13076 4078 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 13076 4078 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 13158 4078 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 13158 4078 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 13240 4078 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 13240 4078 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 12420 4159 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12420 4159 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 12502 4159 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12502 4159 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 12584 4159 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12584 4159 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 12666 4159 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12666 4159 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 12748 4159 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12748 4159 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 12830 4159 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12830 4159 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 12912 4159 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12912 4159 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 12994 4159 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12994 4159 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 13076 4159 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 13076 4159 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 13158 4159 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 13158 4159 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 13240 4159 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 13240 4159 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 12420 4240 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12420 4240 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 12502 4240 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12502 4240 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 12584 4240 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12584 4240 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 12666 4240 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12666 4240 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 12748 4240 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12748 4240 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 12830 4240 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12830 4240 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 12912 4240 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12912 4240 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 12994 4240 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12994 4240 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 13076 4240 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 13076 4240 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 13158 4240 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 13158 4240 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 13240 4240 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 13240 4240 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 12420 4321 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12420 4321 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 12502 4321 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12502 4321 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 12584 4321 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12584 4321 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 12666 4321 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12666 4321 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 12748 4321 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12748 4321 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 12830 4321 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12830 4321 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 12912 4321 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12912 4321 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 12994 4321 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12994 4321 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 13076 4321 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 13076 4321 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 13158 4321 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 13158 4321 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 13240 4321 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 13240 4321 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 12420 4402 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12420 4402 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 12502 4402 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12502 4402 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 12584 4402 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12584 4402 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 12666 4402 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12666 4402 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 12748 4402 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12748 4402 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 12830 4402 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12830 4402 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 12912 4402 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12912 4402 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 12994 4402 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12994 4402 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 13076 4402 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 13076 4402 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 13158 4402 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 13158 4402 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 13240 4402 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 13240 4402 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 12420 4484 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12420 4484 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 12502 4484 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12502 4484 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 12584 4484 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12584 4484 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 12666 4484 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12666 4484 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 12748 4484 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12748 4484 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 12830 4484 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12830 4484 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 12912 4484 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12912 4484 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 12994 4484 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12994 4484 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 13076 4484 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 13076 4484 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 13158 4484 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 13158 4484 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 13240 4484 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 13240 4484 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 12420 4566 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12420 4566 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 12502 4566 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12502 4566 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 12584 4566 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12584 4566 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 12666 4566 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12666 4566 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 12748 4566 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12748 4566 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 12830 4566 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12830 4566 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 12912 4566 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12912 4566 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 12994 4566 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12994 4566 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 13076 4566 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 13076 4566 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 13158 4566 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 13158 4566 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 13240 4566 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 13240 4566 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 12420 4648 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12420 4648 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 12502 4648 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12502 4648 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 12584 4648 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12584 4648 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 12666 4648 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12666 4648 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 12748 4648 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12748 4648 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 12830 4648 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12830 4648 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 12912 4648 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12912 4648 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 12994 4648 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12994 4648 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 13076 4648 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 13076 4648 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 13158 4648 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 13158 4648 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 13240 4648 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 13240 4648 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 12420 4730 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12420 4730 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 12502 4730 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12502 4730 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 12584 4730 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12584 4730 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 12666 4730 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12666 4730 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 12748 4730 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12748 4730 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 12830 4730 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12830 4730 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 12912 4730 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12912 4730 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 12994 4730 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12994 4730 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 13076 4730 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 13076 4730 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 13158 4730 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 13158 4730 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 13240 4730 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 13240 4730 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 12420 4812 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12420 4812 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 12502 4812 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12502 4812 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 12584 4812 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12584 4812 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 12666 4812 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12666 4812 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 12748 4812 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12748 4812 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 12830 4812 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12830 4812 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 12912 4812 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12912 4812 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 12994 4812 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12994 4812 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 13076 4812 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 13076 4812 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 13158 4812 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 13158 4812 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 13240 4812 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 13240 4812 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 12420 4894 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12420 4894 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 12502 4894 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12502 4894 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 12584 4894 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12584 4894 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 12666 4894 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12666 4894 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 12748 4894 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12748 4894 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 12830 4894 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12830 4894 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 12912 4894 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12912 4894 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 12994 4894 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12994 4894 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 13076 4894 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 13076 4894 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 13158 4894 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 13158 4894 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 13240 4894 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 13240 4894 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 12420 676 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12420 676 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 12502 676 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12502 676 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 12584 676 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12584 676 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 12666 676 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12666 676 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 12748 676 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12748 676 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 12830 676 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12830 676 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 12912 676 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12912 676 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 12994 676 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12994 676 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 13076 676 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 13076 676 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 13158 676 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 13158 676 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 13240 676 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 13240 676 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 12420 757 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12420 757 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 12502 757 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12502 757 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 12584 757 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12584 757 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 12666 757 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12666 757 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 12748 757 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12748 757 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 12830 757 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12830 757 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 12912 757 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12912 757 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 12994 757 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12994 757 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 13076 757 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 13076 757 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 13158 757 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 13158 757 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 13240 757 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 13240 757 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 12420 838 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12420 838 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 12502 838 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12502 838 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 12584 838 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12584 838 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 12666 838 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12666 838 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 12748 838 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12748 838 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 12830 838 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12830 838 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 12912 838 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12912 838 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 12994 838 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12994 838 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 13076 838 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 13076 838 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 13158 838 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 13158 838 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 13240 838 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 13240 838 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 12420 919 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12420 919 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 12502 919 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12502 919 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 12584 919 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12584 919 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 12666 919 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12666 919 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 12748 919 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12748 919 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 12830 919 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12830 919 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 12912 919 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12912 919 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 12994 919 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12994 919 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 13076 919 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 13076 919 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 13158 919 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 13158 919 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 13240 919 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 13240 919 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 12420 1000 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12420 1000 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 12502 1000 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12502 1000 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 12584 1000 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12584 1000 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 12666 1000 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12666 1000 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 12748 1000 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12748 1000 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 12830 1000 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12830 1000 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 12912 1000 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12912 1000 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 12994 1000 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12994 1000 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 13076 1000 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 13076 1000 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 13158 1000 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 13158 1000 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 13240 1000 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 13240 1000 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 12420 1081 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12420 1081 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 12502 1081 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12502 1081 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 12584 1081 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12584 1081 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 12666 1081 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12666 1081 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 12748 1081 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12748 1081 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 12830 1081 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12830 1081 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 12912 1081 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12912 1081 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 12994 1081 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12994 1081 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 13076 1081 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 13076 1081 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 13158 1081 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 13158 1081 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 13240 1081 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 13240 1081 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 12420 1162 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12420 1162 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 12502 1162 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12502 1162 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 12584 1162 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12584 1162 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 12666 1162 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12666 1162 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 12748 1162 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12748 1162 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 12830 1162 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12830 1162 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 12912 1162 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12912 1162 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 12994 1162 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12994 1162 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 13076 1162 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 13076 1162 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 13158 1162 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 13158 1162 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 13240 1162 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 13240 1162 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 12420 1243 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12420 1243 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 12502 1243 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12502 1243 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 12584 1243 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12584 1243 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 12666 1243 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12666 1243 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 12748 1243 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12748 1243 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 12830 1243 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12830 1243 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 12912 1243 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12912 1243 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 12994 1243 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12994 1243 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 13076 1243 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 13076 1243 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 13158 1243 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 13158 1243 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 13240 1243 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 13240 1243 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10157 12420 10221 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10157 12420 10221 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10157 12502 10221 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10157 12502 10221 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10157 12584 10221 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10157 12584 10221 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10157 12666 10221 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10157 12666 10221 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10157 12748 10221 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10157 12748 10221 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10157 12830 10221 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10157 12830 10221 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10157 12912 10221 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10157 12912 10221 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10157 12994 10221 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10157 12994 10221 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10157 13076 10221 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10157 13076 10221 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10157 13158 10221 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10157 13158 10221 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10157 13240 10221 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10157 13240 10221 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10238 12420 10302 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10238 12420 10302 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10238 12502 10302 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10238 12502 10302 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10238 12584 10302 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10238 12584 10302 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10238 12666 10302 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10238 12666 10302 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10238 12748 10302 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10238 12748 10302 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10238 12830 10302 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10238 12830 10302 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10238 12912 10302 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10238 12912 10302 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10238 12994 10302 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10238 12994 10302 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10238 13076 10302 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10238 13076 10302 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10238 13158 10302 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10238 13158 10302 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10238 13240 10302 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10238 13240 10302 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10319 12420 10383 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10319 12420 10383 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10319 12502 10383 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10319 12502 10383 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10319 12584 10383 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10319 12584 10383 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10319 12666 10383 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10319 12666 10383 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10319 12748 10383 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10319 12748 10383 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10319 12830 10383 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10319 12830 10383 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10319 12912 10383 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10319 12912 10383 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10319 12994 10383 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10319 12994 10383 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10319 13076 10383 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10319 13076 10383 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10319 13158 10383 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10319 13158 10383 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10319 13240 10383 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10319 13240 10383 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10400 12420 10464 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10400 12420 10464 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10400 12502 10464 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10400 12502 10464 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10400 12584 10464 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10400 12584 10464 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10400 12666 10464 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10400 12666 10464 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10400 12748 10464 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10400 12748 10464 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10400 12830 10464 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10400 12830 10464 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10400 12912 10464 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10400 12912 10464 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10400 12994 10464 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10400 12994 10464 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10400 13076 10464 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10400 13076 10464 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10400 13158 10464 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10400 13158 10464 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10400 13240 10464 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10400 13240 10464 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10481 12420 10545 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10481 12420 10545 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10481 12502 10545 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10481 12502 10545 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10481 12584 10545 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10481 12584 10545 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10481 12666 10545 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10481 12666 10545 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10481 12748 10545 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10481 12748 10545 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10481 12830 10545 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10481 12830 10545 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10481 12912 10545 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10481 12912 10545 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10481 12994 10545 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10481 12994 10545 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10481 13076 10545 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10481 13076 10545 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10481 13158 10545 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10481 13158 10545 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10481 13240 10545 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10481 13240 10545 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10562 12420 10626 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10562 12420 10626 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10562 12502 10626 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10562 12502 10626 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10562 12584 10626 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10562 12584 10626 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10562 12666 10626 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10562 12666 10626 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10562 12748 10626 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10562 12748 10626 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10562 12830 10626 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10562 12830 10626 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10562 12912 10626 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10562 12912 10626 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10562 12994 10626 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10562 12994 10626 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10562 13076 10626 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10562 13076 10626 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10562 13158 10626 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10562 13158 10626 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10562 13240 10626 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10562 13240 10626 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10643 12420 10707 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10643 12420 10707 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10643 12502 10707 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10643 12502 10707 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10643 12584 10707 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10643 12584 10707 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10643 12666 10707 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10643 12666 10707 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10643 12748 10707 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10643 12748 10707 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10643 12830 10707 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10643 12830 10707 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10643 12912 10707 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10643 12912 10707 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10643 12994 10707 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10643 12994 10707 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10643 13076 10707 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10643 13076 10707 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10643 13158 10707 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10643 13158 10707 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10643 13240 10707 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10643 13240 10707 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10724 12420 10788 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10724 12420 10788 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10724 12502 10788 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10724 12502 10788 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10724 12584 10788 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10724 12584 10788 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10724 12666 10788 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10724 12666 10788 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10724 12748 10788 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10724 12748 10788 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10724 12830 10788 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10724 12830 10788 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10724 12912 10788 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10724 12912 10788 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10724 12994 10788 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10724 12994 10788 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10724 13076 10788 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10724 13076 10788 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10724 13158 10788 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10724 13158 10788 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10724 13240 10788 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10724 13240 10788 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10805 12420 10869 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10805 12420 10869 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10805 12502 10869 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10805 12502 10869 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10805 12584 10869 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10805 12584 10869 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10805 12666 10869 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10805 12666 10869 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10805 12748 10869 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10805 12748 10869 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10805 12830 10869 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10805 12830 10869 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10805 12912 10869 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10805 12912 10869 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10805 12994 10869 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10805 12994 10869 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10805 13076 10869 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10805 13076 10869 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10805 13158 10869 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10805 13158 10869 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10805 13240 10869 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10805 13240 10869 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10886 12420 10950 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10886 12420 10950 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10886 12502 10950 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10886 12502 10950 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10886 12584 10950 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10886 12584 10950 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10886 12666 10950 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10886 12666 10950 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10886 12748 10950 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10886 12748 10950 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10886 12830 10950 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10886 12830 10950 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10886 12912 10950 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10886 12912 10950 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10886 12994 10950 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10886 12994 10950 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10886 13076 10950 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10886 13076 10950 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10886 13158 10950 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10886 13158 10950 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10886 13240 10950 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10886 13240 10950 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10967 12420 11031 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10967 12420 11031 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10967 12502 11031 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10967 12502 11031 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10967 12584 11031 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10967 12584 11031 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10967 12666 11031 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10967 12666 11031 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10967 12748 11031 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10967 12748 11031 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10967 12830 11031 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10967 12830 11031 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10967 12912 11031 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10967 12912 11031 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10967 12994 11031 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10967 12994 11031 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10967 13076 11031 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10967 13076 11031 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10967 13158 11031 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10967 13158 11031 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10967 13240 11031 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10967 13240 11031 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11048 12420 11112 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11048 12420 11112 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11048 12502 11112 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11048 12502 11112 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11048 12584 11112 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11048 12584 11112 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11048 12666 11112 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11048 12666 11112 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11048 12748 11112 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11048 12748 11112 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11048 12830 11112 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11048 12830 11112 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11048 12912 11112 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11048 12912 11112 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11048 12994 11112 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11048 12994 11112 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11048 13076 11112 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11048 13076 11112 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11048 13158 11112 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11048 13158 11112 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11048 13240 11112 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11048 13240 11112 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11129 12420 11193 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11129 12420 11193 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11129 12502 11193 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11129 12502 11193 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11129 12584 11193 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11129 12584 11193 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11129 12666 11193 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11129 12666 11193 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11129 12748 11193 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11129 12748 11193 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11129 12830 11193 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11129 12830 11193 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11129 12912 11193 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11129 12912 11193 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11129 12994 11193 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11129 12994 11193 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11129 13076 11193 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11129 13076 11193 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11129 13158 11193 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11129 13158 11193 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11129 13240 11193 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11129 13240 11193 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11210 12420 11274 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11210 12420 11274 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11210 12502 11274 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11210 12502 11274 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11210 12584 11274 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11210 12584 11274 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11210 12666 11274 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11210 12666 11274 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11210 12748 11274 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11210 12748 11274 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11210 12830 11274 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11210 12830 11274 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11210 12912 11274 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11210 12912 11274 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11210 12994 11274 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11210 12994 11274 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11210 13076 11274 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11210 13076 11274 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11210 13158 11274 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11210 13158 11274 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11210 13240 11274 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11210 13240 11274 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11291 12420 11355 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11291 12420 11355 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11291 12502 11355 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11291 12502 11355 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11291 12584 11355 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11291 12584 11355 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11291 12666 11355 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11291 12666 11355 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11291 12748 11355 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11291 12748 11355 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11291 12830 11355 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11291 12830 11355 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11291 12912 11355 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11291 12912 11355 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11291 12994 11355 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11291 12994 11355 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11291 13076 11355 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11291 13076 11355 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11291 13158 11355 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11291 13158 11355 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11291 13240 11355 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11291 13240 11355 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11372 12420 11436 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11372 12420 11436 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11372 12502 11436 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11372 12502 11436 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11372 12584 11436 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11372 12584 11436 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11372 12666 11436 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11372 12666 11436 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11372 12748 11436 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11372 12748 11436 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11372 12830 11436 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11372 12830 11436 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11372 12912 11436 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11372 12912 11436 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11372 12994 11436 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11372 12994 11436 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11372 13076 11436 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11372 13076 11436 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11372 13158 11436 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11372 13158 11436 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11372 13240 11436 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11372 13240 11436 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11453 12420 11517 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11453 12420 11517 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11453 12502 11517 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11453 12502 11517 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11453 12584 11517 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11453 12584 11517 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11453 12666 11517 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11453 12666 11517 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11453 12748 11517 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11453 12748 11517 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11453 12830 11517 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11453 12830 11517 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11453 12912 11517 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11453 12912 11517 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11453 12994 11517 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11453 12994 11517 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11453 13076 11517 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11453 13076 11517 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11453 13158 11517 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11453 13158 11517 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11453 13240 11517 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11453 13240 11517 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11534 12420 11598 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11534 12420 11598 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11534 12502 11598 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11534 12502 11598 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11534 12584 11598 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11534 12584 11598 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11534 12666 11598 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11534 12666 11598 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11534 12748 11598 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11534 12748 11598 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11534 12830 11598 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11534 12830 11598 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11534 12912 11598 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11534 12912 11598 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11534 12994 11598 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11534 12994 11598 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11534 13076 11598 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11534 13076 11598 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11534 13158 11598 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11534 13158 11598 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11534 13240 11598 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11534 13240 11598 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11615 12420 11679 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11615 12420 11679 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11615 12502 11679 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11615 12502 11679 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11615 12584 11679 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11615 12584 11679 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11615 12666 11679 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11615 12666 11679 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11615 12748 11679 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11615 12748 11679 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11615 12830 11679 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11615 12830 11679 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11615 12912 11679 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11615 12912 11679 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11615 12994 11679 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11615 12994 11679 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11615 13076 11679 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11615 13076 11679 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11615 13158 11679 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11615 13158 11679 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11615 13240 11679 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11615 13240 11679 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11696 12420 11760 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11696 12420 11760 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11696 12502 11760 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11696 12502 11760 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11696 12584 11760 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11696 12584 11760 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11696 12666 11760 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11696 12666 11760 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11696 12748 11760 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11696 12748 11760 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11696 12830 11760 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11696 12830 11760 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11696 12912 11760 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11696 12912 11760 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11696 12994 11760 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11696 12994 11760 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11696 13076 11760 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11696 13076 11760 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11696 13158 11760 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11696 13158 11760 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11696 13240 11760 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11696 13240 11760 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11777 12420 11841 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11777 12420 11841 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11777 12502 11841 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11777 12502 11841 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11777 12584 11841 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11777 12584 11841 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11777 12666 11841 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11777 12666 11841 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11777 12748 11841 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11777 12748 11841 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11777 12830 11841 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11777 12830 11841 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11777 12912 11841 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11777 12912 11841 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11777 12994 11841 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11777 12994 11841 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11777 13076 11841 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11777 13076 11841 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11777 13158 11841 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11777 13158 11841 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11777 13240 11841 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11777 13240 11841 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11858 12420 11922 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11858 12420 11922 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11858 12502 11922 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11858 12502 11922 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11858 12584 11922 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11858 12584 11922 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11858 12666 11922 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11858 12666 11922 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11858 12748 11922 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11858 12748 11922 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11858 12830 11922 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11858 12830 11922 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11858 12912 11922 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11858 12912 11922 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11858 12994 11922 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11858 12994 11922 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11858 13076 11922 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11858 13076 11922 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11858 13158 11922 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11858 13158 11922 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11858 13240 11922 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11858 13240 11922 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11939 12420 12003 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11939 12420 12003 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11939 12502 12003 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11939 12502 12003 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11939 12584 12003 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11939 12584 12003 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11939 12666 12003 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11939 12666 12003 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11939 12748 12003 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11939 12748 12003 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11939 12830 12003 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11939 12830 12003 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11939 12912 12003 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11939 12912 12003 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11939 12994 12003 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11939 12994 12003 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11939 13076 12003 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11939 13076 12003 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11939 13158 12003 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11939 13158 12003 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 11939 13240 12003 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11939 13240 12003 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 12420 1324 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12420 1324 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 12502 1324 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12502 1324 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 12584 1324 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12584 1324 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 12666 1324 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12666 1324 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 12748 1324 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12748 1324 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 12830 1324 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12830 1324 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 12912 1324 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12912 1324 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 12994 1324 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12994 1324 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 13076 1324 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 13076 1324 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 13158 1324 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 13158 1324 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 13240 1324 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 13240 1324 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 12420 1405 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12420 1405 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 12502 1405 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12502 1405 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 12584 1405 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12584 1405 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 12666 1405 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12666 1405 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 12748 1405 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12748 1405 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 12830 1405 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12830 1405 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 12912 1405 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12912 1405 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 12994 1405 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12994 1405 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 13076 1405 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 13076 1405 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 13158 1405 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 13158 1405 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 13240 1405 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 13240 1405 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12020 12420 12084 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12020 12420 12084 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12020 12502 12084 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12020 12502 12084 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12020 12584 12084 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12020 12584 12084 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12020 12666 12084 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12020 12666 12084 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12020 12748 12084 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12020 12748 12084 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12020 12830 12084 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12020 12830 12084 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12020 12912 12084 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12020 12912 12084 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12020 12994 12084 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12020 12994 12084 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12020 13076 12084 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12020 13076 12084 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12020 13158 12084 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12020 13158 12084 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12020 13240 12084 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12020 13240 12084 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12101 12420 12165 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12101 12420 12165 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12101 12502 12165 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12101 12502 12165 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12101 12584 12165 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12101 12584 12165 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12101 12666 12165 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12101 12666 12165 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12101 12748 12165 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12101 12748 12165 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12101 12830 12165 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12101 12830 12165 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12101 12912 12165 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12101 12912 12165 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12101 12994 12165 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12101 12994 12165 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12101 13076 12165 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12101 13076 12165 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12101 13158 12165 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12101 13158 12165 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12101 13240 12165 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12101 13240 12165 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12182 12420 12246 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12182 12420 12246 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12182 12502 12246 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12182 12502 12246 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12182 12584 12246 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12182 12584 12246 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12182 12666 12246 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12182 12666 12246 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12182 12748 12246 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12182 12748 12246 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12182 12830 12246 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12182 12830 12246 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12182 12912 12246 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12182 12912 12246 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12182 12994 12246 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12182 12994 12246 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12182 13076 12246 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12182 13076 12246 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12182 13158 12246 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12182 13158 12246 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12182 13240 12246 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12182 13240 12246 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12263 12420 12327 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12263 12420 12327 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12263 12502 12327 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12263 12502 12327 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12263 12584 12327 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12263 12584 12327 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12263 12666 12327 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12263 12666 12327 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12263 12748 12327 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12263 12748 12327 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12263 12830 12327 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12263 12830 12327 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12263 12912 12327 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12263 12912 12327 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12263 12994 12327 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12263 12994 12327 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12263 13076 12327 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12263 13076 12327 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12263 13158 12327 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12263 13158 12327 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12263 13240 12327 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12263 13240 12327 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12344 12420 12408 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12344 12420 12408 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12344 12502 12408 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12344 12502 12408 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12344 12584 12408 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12344 12584 12408 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12344 12666 12408 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12344 12666 12408 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12344 12748 12408 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12344 12748 12408 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12344 12830 12408 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12344 12830 12408 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12344 12912 12408 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12344 12912 12408 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12344 12994 12408 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12344 12994 12408 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12344 13076 12408 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12344 13076 12408 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12344 13158 12408 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12344 13158 12408 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12344 13240 12408 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12344 13240 12408 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12425 12420 12489 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12425 12420 12489 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12425 12502 12489 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12425 12502 12489 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12425 12584 12489 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12425 12584 12489 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12425 12666 12489 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12425 12666 12489 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12425 12748 12489 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12425 12748 12489 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12425 12830 12489 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12425 12830 12489 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12425 12912 12489 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12425 12912 12489 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12425 12994 12489 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12425 12994 12489 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12425 13076 12489 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12425 13076 12489 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12425 13158 12489 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12425 13158 12489 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12425 13240 12489 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12425 13240 12489 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12506 12420 12570 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12506 12420 12570 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12506 12502 12570 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12506 12502 12570 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12506 12584 12570 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12506 12584 12570 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12506 12666 12570 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12506 12666 12570 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12506 12748 12570 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12506 12748 12570 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12506 12830 12570 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12506 12830 12570 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12506 12912 12570 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12506 12912 12570 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12506 12994 12570 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12506 12994 12570 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12506 13076 12570 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12506 13076 12570 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12506 13158 12570 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12506 13158 12570 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12506 13240 12570 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12506 13240 12570 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12587 12420 12651 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12587 12420 12651 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12587 12502 12651 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12587 12502 12651 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12587 12584 12651 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12587 12584 12651 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12587 12666 12651 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12587 12666 12651 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12587 12748 12651 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12587 12748 12651 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12587 12830 12651 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12587 12830 12651 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12587 12912 12651 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12587 12912 12651 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12587 12994 12651 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12587 12994 12651 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12587 13076 12651 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12587 13076 12651 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12587 13158 12651 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12587 13158 12651 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12587 13240 12651 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12587 13240 12651 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12668 12420 12732 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12668 12420 12732 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12668 12502 12732 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12668 12502 12732 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12668 12584 12732 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12668 12584 12732 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12668 12666 12732 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12668 12666 12732 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12668 12748 12732 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12668 12748 12732 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12668 12830 12732 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12668 12830 12732 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12668 12912 12732 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12668 12912 12732 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12668 12994 12732 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12668 12994 12732 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12668 13076 12732 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12668 13076 12732 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12668 13158 12732 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12668 13158 12732 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12668 13240 12732 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12668 13240 12732 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12749 12420 12813 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12749 12420 12813 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12749 12502 12813 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12749 12502 12813 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12749 12584 12813 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12749 12584 12813 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12749 12666 12813 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12749 12666 12813 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12749 12748 12813 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12749 12748 12813 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12749 12830 12813 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12749 12830 12813 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12749 12912 12813 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12749 12912 12813 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12749 12994 12813 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12749 12994 12813 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12749 13076 12813 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12749 13076 12813 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12749 13158 12813 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12749 13158 12813 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12749 13240 12813 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12749 13240 12813 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12830 12420 12894 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12830 12420 12894 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12830 12502 12894 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12830 12502 12894 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12830 12584 12894 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12830 12584 12894 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12830 12666 12894 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12830 12666 12894 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12830 12748 12894 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12830 12748 12894 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12830 12830 12894 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12830 12830 12894 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12830 12912 12894 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12830 12912 12894 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12830 12994 12894 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12830 12994 12894 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12830 13076 12894 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12830 13076 12894 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12830 13158 12894 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12830 13158 12894 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12830 13240 12894 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12830 13240 12894 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12911 12420 12975 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12911 12420 12975 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12911 12502 12975 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12911 12502 12975 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12911 12584 12975 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12911 12584 12975 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12911 12666 12975 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12911 12666 12975 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12911 12748 12975 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12911 12748 12975 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12911 12830 12975 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12911 12830 12975 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12911 12912 12975 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12911 12912 12975 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12911 12994 12975 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12911 12994 12975 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12911 13076 12975 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12911 13076 12975 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12911 13158 12975 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12911 13158 12975 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12911 13240 12975 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12911 13240 12975 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12992 12420 13056 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12992 12420 13056 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12992 12502 13056 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12992 12502 13056 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12992 12584 13056 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12992 12584 13056 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12992 12666 13056 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12992 12666 13056 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12992 12748 13056 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12992 12748 13056 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12992 12830 13056 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12992 12830 13056 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12992 12912 13056 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12992 12912 13056 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12992 12994 13056 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12992 12994 13056 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12992 13076 13056 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12992 13076 13056 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12992 13158 13056 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12992 13158 13056 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 12992 13240 13056 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12992 13240 13056 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13073 12420 13137 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13073 12420 13137 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13073 12502 13137 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13073 12502 13137 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13073 12584 13137 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13073 12584 13137 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13073 12666 13137 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13073 12666 13137 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13073 12748 13137 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13073 12748 13137 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13073 12830 13137 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13073 12830 13137 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13073 12912 13137 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13073 12912 13137 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13073 12994 13137 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13073 12994 13137 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13073 13076 13137 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13073 13076 13137 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13073 13158 13137 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13073 13158 13137 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13073 13240 13137 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13073 13240 13137 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13154 12420 13218 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13154 12420 13218 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13154 12502 13218 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13154 12502 13218 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13154 12584 13218 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13154 12584 13218 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13154 12666 13218 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13154 12666 13218 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13154 12748 13218 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13154 12748 13218 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13154 12830 13218 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13154 12830 13218 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13154 12912 13218 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13154 12912 13218 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13154 12994 13218 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13154 12994 13218 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13154 13076 13218 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13154 13076 13218 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13154 13158 13218 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13154 13158 13218 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13154 13240 13218 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13154 13240 13218 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13235 12420 13299 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13235 12420 13299 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13235 12502 13299 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13235 12502 13299 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13235 12584 13299 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13235 12584 13299 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13235 12666 13299 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13235 12666 13299 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13235 12748 13299 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13235 12748 13299 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13235 12830 13299 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13235 12830 13299 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13235 12912 13299 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13235 12912 13299 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13235 12994 13299 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13235 12994 13299 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13235 13076 13299 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13235 13076 13299 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13235 13158 13299 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13235 13158 13299 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13235 13240 13299 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13235 13240 13299 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13316 12420 13380 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13316 12420 13380 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13316 12502 13380 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13316 12502 13380 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13316 12584 13380 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13316 12584 13380 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13316 12666 13380 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13316 12666 13380 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13316 12748 13380 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13316 12748 13380 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13316 12830 13380 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13316 12830 13380 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13316 12912 13380 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13316 12912 13380 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13316 12994 13380 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13316 12994 13380 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13316 13076 13380 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13316 13076 13380 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13316 13158 13380 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13316 13158 13380 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13316 13240 13380 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13316 13240 13380 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13397 12420 13461 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13397 12420 13461 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13397 12502 13461 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13397 12502 13461 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13397 12584 13461 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13397 12584 13461 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13397 12666 13461 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13397 12666 13461 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13397 12748 13461 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13397 12748 13461 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13397 12830 13461 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13397 12830 13461 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13397 12912 13461 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13397 12912 13461 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13397 12994 13461 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13397 12994 13461 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13397 13076 13461 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13397 13076 13461 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13397 13158 13461 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13397 13158 13461 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13397 13240 13461 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13397 13240 13461 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13478 12420 13542 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13478 12420 13542 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13478 12502 13542 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13478 12502 13542 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13478 12584 13542 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13478 12584 13542 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13478 12666 13542 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13478 12666 13542 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13478 12748 13542 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13478 12748 13542 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13478 12830 13542 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13478 12830 13542 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13478 12912 13542 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13478 12912 13542 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13478 12994 13542 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13478 12994 13542 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13478 13076 13542 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13478 13076 13542 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13478 13158 13542 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13478 13158 13542 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13478 13240 13542 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13478 13240 13542 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13559 12420 13623 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13559 12420 13623 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13559 12502 13623 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13559 12502 13623 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13559 12584 13623 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13559 12584 13623 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13559 12666 13623 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13559 12666 13623 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13559 12748 13623 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13559 12748 13623 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13559 12830 13623 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13559 12830 13623 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13559 12912 13623 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13559 12912 13623 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13559 12994 13623 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13559 12994 13623 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13559 13076 13623 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13559 13076 13623 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13559 13158 13623 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13559 13158 13623 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13559 13240 13623 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13559 13240 13623 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13640 12420 13704 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13640 12420 13704 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13640 12502 13704 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13640 12502 13704 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13640 12584 13704 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13640 12584 13704 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13640 12666 13704 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13640 12666 13704 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13640 12748 13704 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13640 12748 13704 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13640 12830 13704 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13640 12830 13704 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13640 12912 13704 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13640 12912 13704 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13640 12994 13704 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13640 12994 13704 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13640 13076 13704 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13640 13076 13704 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13640 13158 13704 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13640 13158 13704 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13640 13240 13704 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13640 13240 13704 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13721 12420 13785 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13721 12420 13785 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13721 12502 13785 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13721 12502 13785 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13721 12584 13785 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13721 12584 13785 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13721 12666 13785 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13721 12666 13785 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13721 12748 13785 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13721 12748 13785 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13721 12830 13785 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13721 12830 13785 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13721 12912 13785 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13721 12912 13785 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13721 12994 13785 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13721 12994 13785 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13721 13076 13785 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13721 13076 13785 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13721 13158 13785 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13721 13158 13785 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13721 13240 13785 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13721 13240 13785 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13802 12420 13866 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13802 12420 13866 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13802 12502 13866 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13802 12502 13866 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13802 12584 13866 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13802 12584 13866 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13802 12666 13866 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13802 12666 13866 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13802 12748 13866 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13802 12748 13866 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13802 12830 13866 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13802 12830 13866 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13802 12912 13866 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13802 12912 13866 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13802 12994 13866 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13802 12994 13866 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13802 13076 13866 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13802 13076 13866 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13802 13158 13866 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13802 13158 13866 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13802 13240 13866 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13802 13240 13866 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13883 12420 13947 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13883 12420 13947 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13883 12502 13947 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13883 12502 13947 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13883 12584 13947 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13883 12584 13947 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13883 12666 13947 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13883 12666 13947 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13883 12748 13947 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13883 12748 13947 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13883 12830 13947 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13883 12830 13947 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13883 12912 13947 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13883 12912 13947 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13883 12994 13947 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13883 12994 13947 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13883 13076 13947 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13883 13076 13947 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13883 13158 13947 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13883 13158 13947 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13883 13240 13947 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13883 13240 13947 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13964 12420 14028 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13964 12420 14028 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13964 12502 14028 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13964 12502 14028 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13964 12584 14028 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13964 12584 14028 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13964 12666 14028 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13964 12666 14028 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13964 12748 14028 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13964 12748 14028 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13964 12830 14028 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13964 12830 14028 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13964 12912 14028 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13964 12912 14028 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13964 12994 14028 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13964 12994 14028 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13964 13076 14028 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13964 13076 14028 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13964 13158 14028 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13964 13158 14028 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 13964 13240 14028 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13964 13240 14028 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 12420 1486 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12420 1486 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 12502 1486 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12502 1486 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 12584 1486 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12584 1486 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 12666 1486 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12666 1486 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 12748 1486 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12748 1486 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 12830 1486 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12830 1486 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 12912 1486 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12912 1486 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 12994 1486 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12994 1486 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 13076 1486 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 13076 1486 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 13158 1486 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 13158 1486 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 13240 1486 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 13240 1486 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 12420 1567 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12420 1567 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 12502 1567 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12502 1567 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 12584 1567 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12584 1567 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 12666 1567 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12666 1567 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 12748 1567 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12748 1567 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 12830 1567 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12830 1567 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 12912 1567 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12912 1567 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 12994 1567 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12994 1567 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 13076 1567 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 13076 1567 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 13158 1567 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 13158 1567 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 13240 1567 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 13240 1567 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 12420 1648 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12420 1648 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 12502 1648 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12502 1648 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 12584 1648 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12584 1648 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 12666 1648 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12666 1648 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 12748 1648 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12748 1648 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 12830 1648 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12830 1648 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 12912 1648 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12912 1648 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 12994 1648 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12994 1648 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 13076 1648 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 13076 1648 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 13158 1648 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 13158 1648 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 13240 1648 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 13240 1648 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14045 12420 14109 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14045 12420 14109 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14045 12502 14109 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14045 12502 14109 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14045 12584 14109 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14045 12584 14109 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14045 12666 14109 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14045 12666 14109 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14045 12748 14109 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14045 12748 14109 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14045 12830 14109 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14045 12830 14109 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14045 12912 14109 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14045 12912 14109 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14045 12994 14109 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14045 12994 14109 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14045 13076 14109 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14045 13076 14109 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14045 13158 14109 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14045 13158 14109 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14045 13240 14109 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14045 13240 14109 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14126 12420 14190 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14126 12420 14190 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14126 12502 14190 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14126 12502 14190 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14126 12584 14190 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14126 12584 14190 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14126 12666 14190 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14126 12666 14190 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14126 12748 14190 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14126 12748 14190 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14126 12830 14190 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14126 12830 14190 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14126 12912 14190 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14126 12912 14190 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14126 12994 14190 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14126 12994 14190 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14126 13076 14190 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14126 13076 14190 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14126 13158 14190 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14126 13158 14190 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14126 13240 14190 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14126 13240 14190 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14207 12420 14271 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14207 12420 14271 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14207 12502 14271 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14207 12502 14271 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14207 12584 14271 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14207 12584 14271 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14207 12666 14271 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14207 12666 14271 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14207 12748 14271 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14207 12748 14271 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14207 12830 14271 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14207 12830 14271 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14207 12912 14271 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14207 12912 14271 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14207 12994 14271 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14207 12994 14271 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14207 13076 14271 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14207 13076 14271 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14207 13158 14271 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14207 13158 14271 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14207 13240 14271 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14207 13240 14271 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14288 12420 14352 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14288 12420 14352 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14288 12502 14352 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14288 12502 14352 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14288 12584 14352 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14288 12584 14352 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14288 12666 14352 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14288 12666 14352 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14288 12748 14352 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14288 12748 14352 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14288 12830 14352 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14288 12830 14352 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14288 12912 14352 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14288 12912 14352 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14288 12994 14352 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14288 12994 14352 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14288 13076 14352 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14288 13076 14352 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14288 13158 14352 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14288 13158 14352 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14288 13240 14352 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14288 13240 14352 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14369 12420 14433 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14369 12420 14433 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14369 12502 14433 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14369 12502 14433 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14369 12584 14433 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14369 12584 14433 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14369 12666 14433 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14369 12666 14433 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14369 12748 14433 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14369 12748 14433 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14369 12830 14433 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14369 12830 14433 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14369 12912 14433 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14369 12912 14433 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14369 12994 14433 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14369 12994 14433 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14369 13076 14433 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14369 13076 14433 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14369 13158 14433 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14369 13158 14433 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14369 13240 14433 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14369 13240 14433 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14451 12420 14515 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14451 12420 14515 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14451 12502 14515 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14451 12502 14515 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14451 12584 14515 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14451 12584 14515 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14451 12666 14515 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14451 12666 14515 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14451 12748 14515 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14451 12748 14515 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14451 12830 14515 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14451 12830 14515 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14451 12912 14515 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14451 12912 14515 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14451 12994 14515 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14451 12994 14515 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14451 13076 14515 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14451 13076 14515 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14451 13158 14515 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14451 13158 14515 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14451 13240 14515 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14451 13240 14515 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14533 12420 14597 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14533 12420 14597 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14533 12502 14597 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14533 12502 14597 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14533 12584 14597 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14533 12584 14597 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14533 12666 14597 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14533 12666 14597 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14533 12748 14597 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14533 12748 14597 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14533 12830 14597 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14533 12830 14597 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14533 12912 14597 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14533 12912 14597 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14533 12994 14597 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14533 12994 14597 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14533 13076 14597 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14533 13076 14597 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14533 13158 14597 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14533 13158 14597 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14533 13240 14597 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14533 13240 14597 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14615 12420 14679 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14615 12420 14679 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14615 12502 14679 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14615 12502 14679 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14615 12584 14679 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14615 12584 14679 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14615 12666 14679 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14615 12666 14679 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14615 12748 14679 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14615 12748 14679 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14615 12830 14679 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14615 12830 14679 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14615 12912 14679 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14615 12912 14679 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14615 12994 14679 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14615 12994 14679 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14615 13076 14679 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14615 13076 14679 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14615 13158 14679 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14615 13158 14679 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14615 13240 14679 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14615 13240 14679 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14697 12420 14761 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14697 12420 14761 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14697 12502 14761 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14697 12502 14761 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14697 12584 14761 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14697 12584 14761 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14697 12666 14761 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14697 12666 14761 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14697 12748 14761 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14697 12748 14761 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14697 12830 14761 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14697 12830 14761 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14697 12912 14761 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14697 12912 14761 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14697 12994 14761 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14697 12994 14761 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14697 13076 14761 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14697 13076 14761 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14697 13158 14761 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14697 13158 14761 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14697 13240 14761 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14697 13240 14761 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14779 12420 14843 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14779 12420 14843 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14779 12502 14843 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14779 12502 14843 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14779 12584 14843 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14779 12584 14843 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14779 12666 14843 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14779 12666 14843 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14779 12748 14843 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14779 12748 14843 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14779 12830 14843 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14779 12830 14843 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14779 12912 14843 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14779 12912 14843 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14779 12994 14843 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14779 12994 14843 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14779 13076 14843 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14779 13076 14843 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14779 13158 14843 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14779 13158 14843 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14779 13240 14843 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14779 13240 14843 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14861 12420 14925 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14861 12420 14925 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14861 12502 14925 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14861 12502 14925 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14861 12584 14925 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14861 12584 14925 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14861 12666 14925 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14861 12666 14925 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14861 12748 14925 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14861 12748 14925 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14861 12830 14925 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14861 12830 14925 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14861 12912 14925 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14861 12912 14925 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14861 12994 14925 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14861 12994 14925 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14861 13076 14925 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14861 13076 14925 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14861 13158 14925 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14861 13158 14925 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14861 13240 14925 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14861 13240 14925 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 12420 1729 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12420 1729 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 12502 1729 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12502 1729 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 12584 1729 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12584 1729 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 12666 1729 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12666 1729 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 12748 1729 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12748 1729 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 12830 1729 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12830 1729 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 12912 1729 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12912 1729 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 12994 1729 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12994 1729 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 13076 1729 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 13076 1729 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 13158 1729 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 13158 1729 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 13240 1729 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 13240 1729 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 12420 1810 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12420 1810 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 12502 1810 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12502 1810 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 12584 1810 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12584 1810 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 12666 1810 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12666 1810 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 12748 1810 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12748 1810 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 12830 1810 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12830 1810 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 12912 1810 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12912 1810 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 12994 1810 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12994 1810 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 13076 1810 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 13076 1810 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 13158 1810 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 13158 1810 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 13240 1810 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 13240 1810 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 12420 1891 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12420 1891 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 12502 1891 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12502 1891 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 12584 1891 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12584 1891 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 12666 1891 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12666 1891 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 12748 1891 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12748 1891 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 12830 1891 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12830 1891 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 12912 1891 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12912 1891 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 12994 1891 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12994 1891 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 13076 1891 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 13076 1891 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 13158 1891 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 13158 1891 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 13240 1891 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 13240 1891 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 12420 1972 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12420 1972 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 12502 1972 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12502 1972 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 12584 1972 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12584 1972 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 12666 1972 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12666 1972 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 12748 1972 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12748 1972 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 12830 1972 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12830 1972 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 12912 1972 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12912 1972 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 12994 1972 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12994 1972 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 13076 1972 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 13076 1972 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 13158 1972 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 13158 1972 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 13240 1972 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 13240 1972 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 12420 2053 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12420 2053 12484 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 12502 2053 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12502 2053 12566 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 12584 2053 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12584 2053 12648 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 12666 2053 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12666 2053 12730 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 12748 2053 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12748 2053 12812 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 12830 2053 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12830 2053 12894 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 12912 2053 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12912 2053 12976 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 12994 2053 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12994 2053 13058 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 13076 2053 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 13076 2053 13140 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 13158 2053 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 13158 2053 13222 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 13240 2053 13304 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 13240 2053 13304 1 VDDIO_Q
port 1 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 15000 39600
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string LEFsymmetry X Y R90
string GDS_END 5947526
string GDS_START 5363942
<< end >>
