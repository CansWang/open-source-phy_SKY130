magic
tech sky130A
magscale 1 2
timestamp 1619862920
<< checkpaint >>
rect -3546 -2154 18508 4578
<< dnwell >>
rect 11876 1604 17168 3110
<< nwell >>
rect 366 1613 4775 3116
rect 5290 1613 6758 3116
rect 7158 1613 8896 3116
rect 11796 3116 17248 3190
rect 9436 2904 17248 3116
rect 9436 1810 12082 2904
rect 14468 1810 14636 2904
rect 16962 1810 17248 2904
rect 9436 1613 17248 1810
rect 11796 1524 17248 1613
rect 1457 965 2403 1133
rect 2887 965 3498 1133
rect 3898 4 5716 1184
<< pwell >>
rect 184 3212 9078 3298
rect 184 2864 270 3212
rect -135 2212 270 2864
rect 184 1517 270 2212
rect 4870 1517 5159 3212
rect 6851 1517 7059 3212
rect 8992 1517 9078 3212
rect 12182 2718 14253 2804
rect 12192 1884 14244 2718
rect 14827 2718 16898 2804
rect 14836 1884 16888 2718
rect 184 1431 9078 1517
rect 1473 22 2343 108
rect 2953 22 3432 108
rect 5866 522 16038 1174
rect 5866 220 6616 522
rect 5890 100 6616 220
rect 7202 100 15130 522
rect 15504 122 16038 522
rect 15504 100 16024 122
rect 5890 14 16024 100
<< pmos >>
rect 3987 148 4037 1148
rect 4093 148 4143 1148
rect 4199 148 4249 1148
rect 4305 148 4355 1148
rect 4411 148 4461 1148
rect 4517 148 4567 1148
rect 4623 148 4673 1148
rect 4729 148 4779 1148
rect 4835 148 4885 1148
rect 4941 148 4991 1148
rect 5047 148 5097 1148
rect 5153 148 5203 1148
rect 5259 148 5309 1148
rect 5365 148 5415 1148
rect 5471 148 5521 1148
rect 5577 148 5627 1148
<< mvnmos >>
rect -56 2238 44 2838
rect 5945 948 6105 1148
rect 6161 948 6321 1148
rect 6377 948 6537 1148
rect 5945 618 6105 818
rect 6161 618 6321 818
rect 6377 618 6537 818
rect 6703 548 6803 1148
rect 6859 548 6959 1148
rect 7015 548 7115 1148
rect 5945 246 6105 446
rect 6161 246 6321 446
rect 6377 246 6537 446
rect 7281 148 7381 1148
rect 7547 148 7707 1148
rect 7763 148 7923 1148
rect 7979 148 8139 1148
rect 8195 148 8355 1148
rect 8411 148 8571 1148
rect 8627 148 8787 1148
rect 8843 148 9003 1148
rect 9059 148 9219 1148
rect 9275 148 9435 1148
rect 9491 148 9651 1148
rect 9707 148 9867 1148
rect 9923 148 10083 1148
rect 10139 148 10299 1148
rect 10355 148 10515 1148
rect 10571 148 10731 1148
rect 10787 148 10947 1148
rect 11003 148 11163 1148
rect 11219 148 11379 1148
rect 11435 148 11595 1148
rect 11651 148 11811 1148
rect 11867 148 12027 1148
rect 12083 148 12243 1148
rect 12299 148 12459 1148
rect 12515 148 12675 1148
rect 12731 148 12891 1148
rect 12947 148 13107 1148
rect 13163 148 13323 1148
rect 13379 148 13539 1148
rect 13595 148 13755 1148
rect 13811 148 13971 1148
rect 14027 148 14187 1148
rect 14243 148 14403 1148
rect 14459 148 14619 1148
rect 14675 148 14835 1148
rect 14891 148 15051 1148
rect 15217 548 15417 1148
rect 15583 148 15743 1148
rect 15799 148 15959 1148
<< mvpmos >>
rect 765 1921 865 2921
rect 921 1921 1021 2921
rect 1187 1921 1287 2921
rect 1343 1921 1443 2921
rect 1499 1921 1599 2921
rect 1655 1921 1755 2921
rect 1811 1921 1911 2921
rect 1967 1921 2067 2921
rect 2123 1921 2223 2921
rect 2279 1921 2379 2921
rect 2435 1921 2535 2921
rect 2591 1921 2691 2921
rect 2747 1921 2847 2921
rect 2903 1921 3003 2921
rect 3059 1921 3159 2921
rect 3215 1921 3315 2921
rect 3371 1921 3471 2921
rect 3527 1921 3627 2921
rect 3683 1921 3783 2921
rect 3839 1921 3939 2921
rect 3995 1921 4095 2921
rect 4261 1921 4361 2521
rect 4417 1921 4517 2521
rect 5547 1921 5647 2921
rect 5703 1921 5803 2921
rect 5859 1921 6019 2921
rect 6075 1921 6235 2921
rect 6401 2321 6501 2521
rect 7415 1921 7575 2921
rect 7631 1921 7791 2921
rect 7847 1921 8007 2921
rect 8063 1921 8163 2921
rect 8219 1921 8319 2921
rect 8375 1921 8475 2921
rect 8531 1921 8631 2921
rect 9693 1921 9793 2921
rect 9849 1921 9949 2921
rect 10005 1921 10105 2921
rect 10161 1921 10261 2921
rect 10317 1921 10417 2921
rect 10473 1921 10573 2921
rect 10629 1921 10729 2921
rect 10785 1921 10885 2921
rect 10941 1921 11041 2921
rect 11097 1921 11197 2921
rect 11253 1921 11353 2921
rect 11409 1921 11509 2921
<< mvnnmos >>
rect 12218 2435 14218 2615
rect 12218 2199 14218 2379
rect 12218 1963 14218 2143
rect 14862 2435 16862 2615
rect 14862 2199 16862 2379
rect 14862 1963 16862 2143
<< pdiff >>
rect 3934 1078 3987 1148
rect 3934 1044 3942 1078
rect 3976 1044 3987 1078
rect 3934 1010 3987 1044
rect 3934 976 3942 1010
rect 3976 976 3987 1010
rect 3934 942 3987 976
rect 3934 908 3942 942
rect 3976 908 3987 942
rect 3934 874 3987 908
rect 3934 840 3942 874
rect 3976 840 3987 874
rect 3934 806 3987 840
rect 3934 772 3942 806
rect 3976 772 3987 806
rect 3934 738 3987 772
rect 3934 704 3942 738
rect 3976 704 3987 738
rect 3934 670 3987 704
rect 3934 636 3942 670
rect 3976 636 3987 670
rect 3934 602 3987 636
rect 3934 568 3942 602
rect 3976 568 3987 602
rect 3934 534 3987 568
rect 3934 500 3942 534
rect 3976 500 3987 534
rect 3934 466 3987 500
rect 3934 432 3942 466
rect 3976 432 3987 466
rect 3934 398 3987 432
rect 3934 364 3942 398
rect 3976 364 3987 398
rect 3934 330 3987 364
rect 3934 296 3942 330
rect 3976 296 3987 330
rect 3934 262 3987 296
rect 3934 228 3942 262
rect 3976 228 3987 262
rect 3934 194 3987 228
rect 3934 160 3942 194
rect 3976 160 3987 194
rect 3934 148 3987 160
rect 4037 1078 4093 1148
rect 4037 1044 4048 1078
rect 4082 1044 4093 1078
rect 4037 1010 4093 1044
rect 4037 976 4048 1010
rect 4082 976 4093 1010
rect 4037 942 4093 976
rect 4037 908 4048 942
rect 4082 908 4093 942
rect 4037 874 4093 908
rect 4037 840 4048 874
rect 4082 840 4093 874
rect 4037 806 4093 840
rect 4037 772 4048 806
rect 4082 772 4093 806
rect 4037 738 4093 772
rect 4037 704 4048 738
rect 4082 704 4093 738
rect 4037 670 4093 704
rect 4037 636 4048 670
rect 4082 636 4093 670
rect 4037 602 4093 636
rect 4037 568 4048 602
rect 4082 568 4093 602
rect 4037 534 4093 568
rect 4037 500 4048 534
rect 4082 500 4093 534
rect 4037 466 4093 500
rect 4037 432 4048 466
rect 4082 432 4093 466
rect 4037 398 4093 432
rect 4037 364 4048 398
rect 4082 364 4093 398
rect 4037 330 4093 364
rect 4037 296 4048 330
rect 4082 296 4093 330
rect 4037 262 4093 296
rect 4037 228 4048 262
rect 4082 228 4093 262
rect 4037 194 4093 228
rect 4037 160 4048 194
rect 4082 160 4093 194
rect 4037 148 4093 160
rect 4143 1078 4199 1148
rect 4143 1044 4154 1078
rect 4188 1044 4199 1078
rect 4143 1010 4199 1044
rect 4143 976 4154 1010
rect 4188 976 4199 1010
rect 4143 942 4199 976
rect 4143 908 4154 942
rect 4188 908 4199 942
rect 4143 874 4199 908
rect 4143 840 4154 874
rect 4188 840 4199 874
rect 4143 806 4199 840
rect 4143 772 4154 806
rect 4188 772 4199 806
rect 4143 738 4199 772
rect 4143 704 4154 738
rect 4188 704 4199 738
rect 4143 670 4199 704
rect 4143 636 4154 670
rect 4188 636 4199 670
rect 4143 602 4199 636
rect 4143 568 4154 602
rect 4188 568 4199 602
rect 4143 534 4199 568
rect 4143 500 4154 534
rect 4188 500 4199 534
rect 4143 466 4199 500
rect 4143 432 4154 466
rect 4188 432 4199 466
rect 4143 398 4199 432
rect 4143 364 4154 398
rect 4188 364 4199 398
rect 4143 330 4199 364
rect 4143 296 4154 330
rect 4188 296 4199 330
rect 4143 262 4199 296
rect 4143 228 4154 262
rect 4188 228 4199 262
rect 4143 194 4199 228
rect 4143 160 4154 194
rect 4188 160 4199 194
rect 4143 148 4199 160
rect 4249 1078 4305 1148
rect 4249 1044 4260 1078
rect 4294 1044 4305 1078
rect 4249 1010 4305 1044
rect 4249 976 4260 1010
rect 4294 976 4305 1010
rect 4249 942 4305 976
rect 4249 908 4260 942
rect 4294 908 4305 942
rect 4249 874 4305 908
rect 4249 840 4260 874
rect 4294 840 4305 874
rect 4249 806 4305 840
rect 4249 772 4260 806
rect 4294 772 4305 806
rect 4249 738 4305 772
rect 4249 704 4260 738
rect 4294 704 4305 738
rect 4249 670 4305 704
rect 4249 636 4260 670
rect 4294 636 4305 670
rect 4249 602 4305 636
rect 4249 568 4260 602
rect 4294 568 4305 602
rect 4249 534 4305 568
rect 4249 500 4260 534
rect 4294 500 4305 534
rect 4249 466 4305 500
rect 4249 432 4260 466
rect 4294 432 4305 466
rect 4249 398 4305 432
rect 4249 364 4260 398
rect 4294 364 4305 398
rect 4249 330 4305 364
rect 4249 296 4260 330
rect 4294 296 4305 330
rect 4249 262 4305 296
rect 4249 228 4260 262
rect 4294 228 4305 262
rect 4249 194 4305 228
rect 4249 160 4260 194
rect 4294 160 4305 194
rect 4249 148 4305 160
rect 4355 1078 4411 1148
rect 4355 1044 4366 1078
rect 4400 1044 4411 1078
rect 4355 1010 4411 1044
rect 4355 976 4366 1010
rect 4400 976 4411 1010
rect 4355 942 4411 976
rect 4355 908 4366 942
rect 4400 908 4411 942
rect 4355 874 4411 908
rect 4355 840 4366 874
rect 4400 840 4411 874
rect 4355 806 4411 840
rect 4355 772 4366 806
rect 4400 772 4411 806
rect 4355 738 4411 772
rect 4355 704 4366 738
rect 4400 704 4411 738
rect 4355 670 4411 704
rect 4355 636 4366 670
rect 4400 636 4411 670
rect 4355 602 4411 636
rect 4355 568 4366 602
rect 4400 568 4411 602
rect 4355 534 4411 568
rect 4355 500 4366 534
rect 4400 500 4411 534
rect 4355 466 4411 500
rect 4355 432 4366 466
rect 4400 432 4411 466
rect 4355 398 4411 432
rect 4355 364 4366 398
rect 4400 364 4411 398
rect 4355 330 4411 364
rect 4355 296 4366 330
rect 4400 296 4411 330
rect 4355 262 4411 296
rect 4355 228 4366 262
rect 4400 228 4411 262
rect 4355 194 4411 228
rect 4355 160 4366 194
rect 4400 160 4411 194
rect 4355 148 4411 160
rect 4461 1078 4517 1148
rect 4461 1044 4472 1078
rect 4506 1044 4517 1078
rect 4461 1010 4517 1044
rect 4461 976 4472 1010
rect 4506 976 4517 1010
rect 4461 942 4517 976
rect 4461 908 4472 942
rect 4506 908 4517 942
rect 4461 874 4517 908
rect 4461 840 4472 874
rect 4506 840 4517 874
rect 4461 806 4517 840
rect 4461 772 4472 806
rect 4506 772 4517 806
rect 4461 738 4517 772
rect 4461 704 4472 738
rect 4506 704 4517 738
rect 4461 670 4517 704
rect 4461 636 4472 670
rect 4506 636 4517 670
rect 4461 602 4517 636
rect 4461 568 4472 602
rect 4506 568 4517 602
rect 4461 534 4517 568
rect 4461 500 4472 534
rect 4506 500 4517 534
rect 4461 466 4517 500
rect 4461 432 4472 466
rect 4506 432 4517 466
rect 4461 398 4517 432
rect 4461 364 4472 398
rect 4506 364 4517 398
rect 4461 330 4517 364
rect 4461 296 4472 330
rect 4506 296 4517 330
rect 4461 262 4517 296
rect 4461 228 4472 262
rect 4506 228 4517 262
rect 4461 194 4517 228
rect 4461 160 4472 194
rect 4506 160 4517 194
rect 4461 148 4517 160
rect 4567 1078 4623 1148
rect 4567 1044 4578 1078
rect 4612 1044 4623 1078
rect 4567 1010 4623 1044
rect 4567 976 4578 1010
rect 4612 976 4623 1010
rect 4567 942 4623 976
rect 4567 908 4578 942
rect 4612 908 4623 942
rect 4567 874 4623 908
rect 4567 840 4578 874
rect 4612 840 4623 874
rect 4567 806 4623 840
rect 4567 772 4578 806
rect 4612 772 4623 806
rect 4567 738 4623 772
rect 4567 704 4578 738
rect 4612 704 4623 738
rect 4567 670 4623 704
rect 4567 636 4578 670
rect 4612 636 4623 670
rect 4567 602 4623 636
rect 4567 568 4578 602
rect 4612 568 4623 602
rect 4567 534 4623 568
rect 4567 500 4578 534
rect 4612 500 4623 534
rect 4567 466 4623 500
rect 4567 432 4578 466
rect 4612 432 4623 466
rect 4567 398 4623 432
rect 4567 364 4578 398
rect 4612 364 4623 398
rect 4567 330 4623 364
rect 4567 296 4578 330
rect 4612 296 4623 330
rect 4567 262 4623 296
rect 4567 228 4578 262
rect 4612 228 4623 262
rect 4567 194 4623 228
rect 4567 160 4578 194
rect 4612 160 4623 194
rect 4567 148 4623 160
rect 4673 1078 4729 1148
rect 4673 1044 4684 1078
rect 4718 1044 4729 1078
rect 4673 1010 4729 1044
rect 4673 976 4684 1010
rect 4718 976 4729 1010
rect 4673 942 4729 976
rect 4673 908 4684 942
rect 4718 908 4729 942
rect 4673 874 4729 908
rect 4673 840 4684 874
rect 4718 840 4729 874
rect 4673 806 4729 840
rect 4673 772 4684 806
rect 4718 772 4729 806
rect 4673 738 4729 772
rect 4673 704 4684 738
rect 4718 704 4729 738
rect 4673 670 4729 704
rect 4673 636 4684 670
rect 4718 636 4729 670
rect 4673 602 4729 636
rect 4673 568 4684 602
rect 4718 568 4729 602
rect 4673 534 4729 568
rect 4673 500 4684 534
rect 4718 500 4729 534
rect 4673 466 4729 500
rect 4673 432 4684 466
rect 4718 432 4729 466
rect 4673 398 4729 432
rect 4673 364 4684 398
rect 4718 364 4729 398
rect 4673 330 4729 364
rect 4673 296 4684 330
rect 4718 296 4729 330
rect 4673 262 4729 296
rect 4673 228 4684 262
rect 4718 228 4729 262
rect 4673 194 4729 228
rect 4673 160 4684 194
rect 4718 160 4729 194
rect 4673 148 4729 160
rect 4779 1078 4835 1148
rect 4779 1044 4790 1078
rect 4824 1044 4835 1078
rect 4779 1010 4835 1044
rect 4779 976 4790 1010
rect 4824 976 4835 1010
rect 4779 942 4835 976
rect 4779 908 4790 942
rect 4824 908 4835 942
rect 4779 874 4835 908
rect 4779 840 4790 874
rect 4824 840 4835 874
rect 4779 806 4835 840
rect 4779 772 4790 806
rect 4824 772 4835 806
rect 4779 738 4835 772
rect 4779 704 4790 738
rect 4824 704 4835 738
rect 4779 670 4835 704
rect 4779 636 4790 670
rect 4824 636 4835 670
rect 4779 602 4835 636
rect 4779 568 4790 602
rect 4824 568 4835 602
rect 4779 534 4835 568
rect 4779 500 4790 534
rect 4824 500 4835 534
rect 4779 466 4835 500
rect 4779 432 4790 466
rect 4824 432 4835 466
rect 4779 398 4835 432
rect 4779 364 4790 398
rect 4824 364 4835 398
rect 4779 330 4835 364
rect 4779 296 4790 330
rect 4824 296 4835 330
rect 4779 262 4835 296
rect 4779 228 4790 262
rect 4824 228 4835 262
rect 4779 194 4835 228
rect 4779 160 4790 194
rect 4824 160 4835 194
rect 4779 148 4835 160
rect 4885 1078 4941 1148
rect 4885 1044 4896 1078
rect 4930 1044 4941 1078
rect 4885 1010 4941 1044
rect 4885 976 4896 1010
rect 4930 976 4941 1010
rect 4885 942 4941 976
rect 4885 908 4896 942
rect 4930 908 4941 942
rect 4885 874 4941 908
rect 4885 840 4896 874
rect 4930 840 4941 874
rect 4885 806 4941 840
rect 4885 772 4896 806
rect 4930 772 4941 806
rect 4885 738 4941 772
rect 4885 704 4896 738
rect 4930 704 4941 738
rect 4885 670 4941 704
rect 4885 636 4896 670
rect 4930 636 4941 670
rect 4885 602 4941 636
rect 4885 568 4896 602
rect 4930 568 4941 602
rect 4885 534 4941 568
rect 4885 500 4896 534
rect 4930 500 4941 534
rect 4885 466 4941 500
rect 4885 432 4896 466
rect 4930 432 4941 466
rect 4885 398 4941 432
rect 4885 364 4896 398
rect 4930 364 4941 398
rect 4885 330 4941 364
rect 4885 296 4896 330
rect 4930 296 4941 330
rect 4885 262 4941 296
rect 4885 228 4896 262
rect 4930 228 4941 262
rect 4885 194 4941 228
rect 4885 160 4896 194
rect 4930 160 4941 194
rect 4885 148 4941 160
rect 4991 1078 5047 1148
rect 4991 1044 5002 1078
rect 5036 1044 5047 1078
rect 4991 1010 5047 1044
rect 4991 976 5002 1010
rect 5036 976 5047 1010
rect 4991 942 5047 976
rect 4991 908 5002 942
rect 5036 908 5047 942
rect 4991 874 5047 908
rect 4991 840 5002 874
rect 5036 840 5047 874
rect 4991 806 5047 840
rect 4991 772 5002 806
rect 5036 772 5047 806
rect 4991 738 5047 772
rect 4991 704 5002 738
rect 5036 704 5047 738
rect 4991 670 5047 704
rect 4991 636 5002 670
rect 5036 636 5047 670
rect 4991 602 5047 636
rect 4991 568 5002 602
rect 5036 568 5047 602
rect 4991 534 5047 568
rect 4991 500 5002 534
rect 5036 500 5047 534
rect 4991 466 5047 500
rect 4991 432 5002 466
rect 5036 432 5047 466
rect 4991 398 5047 432
rect 4991 364 5002 398
rect 5036 364 5047 398
rect 4991 330 5047 364
rect 4991 296 5002 330
rect 5036 296 5047 330
rect 4991 262 5047 296
rect 4991 228 5002 262
rect 5036 228 5047 262
rect 4991 194 5047 228
rect 4991 160 5002 194
rect 5036 160 5047 194
rect 4991 148 5047 160
rect 5097 1078 5153 1148
rect 5097 1044 5108 1078
rect 5142 1044 5153 1078
rect 5097 1010 5153 1044
rect 5097 976 5108 1010
rect 5142 976 5153 1010
rect 5097 942 5153 976
rect 5097 908 5108 942
rect 5142 908 5153 942
rect 5097 874 5153 908
rect 5097 840 5108 874
rect 5142 840 5153 874
rect 5097 806 5153 840
rect 5097 772 5108 806
rect 5142 772 5153 806
rect 5097 738 5153 772
rect 5097 704 5108 738
rect 5142 704 5153 738
rect 5097 670 5153 704
rect 5097 636 5108 670
rect 5142 636 5153 670
rect 5097 602 5153 636
rect 5097 568 5108 602
rect 5142 568 5153 602
rect 5097 534 5153 568
rect 5097 500 5108 534
rect 5142 500 5153 534
rect 5097 466 5153 500
rect 5097 432 5108 466
rect 5142 432 5153 466
rect 5097 398 5153 432
rect 5097 364 5108 398
rect 5142 364 5153 398
rect 5097 330 5153 364
rect 5097 296 5108 330
rect 5142 296 5153 330
rect 5097 262 5153 296
rect 5097 228 5108 262
rect 5142 228 5153 262
rect 5097 194 5153 228
rect 5097 160 5108 194
rect 5142 160 5153 194
rect 5097 148 5153 160
rect 5203 1078 5259 1148
rect 5203 1044 5214 1078
rect 5248 1044 5259 1078
rect 5203 1010 5259 1044
rect 5203 976 5214 1010
rect 5248 976 5259 1010
rect 5203 942 5259 976
rect 5203 908 5214 942
rect 5248 908 5259 942
rect 5203 874 5259 908
rect 5203 840 5214 874
rect 5248 840 5259 874
rect 5203 806 5259 840
rect 5203 772 5214 806
rect 5248 772 5259 806
rect 5203 738 5259 772
rect 5203 704 5214 738
rect 5248 704 5259 738
rect 5203 670 5259 704
rect 5203 636 5214 670
rect 5248 636 5259 670
rect 5203 602 5259 636
rect 5203 568 5214 602
rect 5248 568 5259 602
rect 5203 534 5259 568
rect 5203 500 5214 534
rect 5248 500 5259 534
rect 5203 466 5259 500
rect 5203 432 5214 466
rect 5248 432 5259 466
rect 5203 398 5259 432
rect 5203 364 5214 398
rect 5248 364 5259 398
rect 5203 330 5259 364
rect 5203 296 5214 330
rect 5248 296 5259 330
rect 5203 262 5259 296
rect 5203 228 5214 262
rect 5248 228 5259 262
rect 5203 194 5259 228
rect 5203 160 5214 194
rect 5248 160 5259 194
rect 5203 148 5259 160
rect 5309 1078 5365 1148
rect 5309 1044 5320 1078
rect 5354 1044 5365 1078
rect 5309 1010 5365 1044
rect 5309 976 5320 1010
rect 5354 976 5365 1010
rect 5309 942 5365 976
rect 5309 908 5320 942
rect 5354 908 5365 942
rect 5309 874 5365 908
rect 5309 840 5320 874
rect 5354 840 5365 874
rect 5309 806 5365 840
rect 5309 772 5320 806
rect 5354 772 5365 806
rect 5309 738 5365 772
rect 5309 704 5320 738
rect 5354 704 5365 738
rect 5309 670 5365 704
rect 5309 636 5320 670
rect 5354 636 5365 670
rect 5309 602 5365 636
rect 5309 568 5320 602
rect 5354 568 5365 602
rect 5309 534 5365 568
rect 5309 500 5320 534
rect 5354 500 5365 534
rect 5309 466 5365 500
rect 5309 432 5320 466
rect 5354 432 5365 466
rect 5309 398 5365 432
rect 5309 364 5320 398
rect 5354 364 5365 398
rect 5309 330 5365 364
rect 5309 296 5320 330
rect 5354 296 5365 330
rect 5309 262 5365 296
rect 5309 228 5320 262
rect 5354 228 5365 262
rect 5309 194 5365 228
rect 5309 160 5320 194
rect 5354 160 5365 194
rect 5309 148 5365 160
rect 5415 1078 5471 1148
rect 5415 1044 5426 1078
rect 5460 1044 5471 1078
rect 5415 1010 5471 1044
rect 5415 976 5426 1010
rect 5460 976 5471 1010
rect 5415 942 5471 976
rect 5415 908 5426 942
rect 5460 908 5471 942
rect 5415 874 5471 908
rect 5415 840 5426 874
rect 5460 840 5471 874
rect 5415 806 5471 840
rect 5415 772 5426 806
rect 5460 772 5471 806
rect 5415 738 5471 772
rect 5415 704 5426 738
rect 5460 704 5471 738
rect 5415 670 5471 704
rect 5415 636 5426 670
rect 5460 636 5471 670
rect 5415 602 5471 636
rect 5415 568 5426 602
rect 5460 568 5471 602
rect 5415 534 5471 568
rect 5415 500 5426 534
rect 5460 500 5471 534
rect 5415 466 5471 500
rect 5415 432 5426 466
rect 5460 432 5471 466
rect 5415 398 5471 432
rect 5415 364 5426 398
rect 5460 364 5471 398
rect 5415 330 5471 364
rect 5415 296 5426 330
rect 5460 296 5471 330
rect 5415 262 5471 296
rect 5415 228 5426 262
rect 5460 228 5471 262
rect 5415 194 5471 228
rect 5415 160 5426 194
rect 5460 160 5471 194
rect 5415 148 5471 160
rect 5521 1078 5577 1148
rect 5521 1044 5532 1078
rect 5566 1044 5577 1078
rect 5521 1010 5577 1044
rect 5521 976 5532 1010
rect 5566 976 5577 1010
rect 5521 942 5577 976
rect 5521 908 5532 942
rect 5566 908 5577 942
rect 5521 874 5577 908
rect 5521 840 5532 874
rect 5566 840 5577 874
rect 5521 806 5577 840
rect 5521 772 5532 806
rect 5566 772 5577 806
rect 5521 738 5577 772
rect 5521 704 5532 738
rect 5566 704 5577 738
rect 5521 670 5577 704
rect 5521 636 5532 670
rect 5566 636 5577 670
rect 5521 602 5577 636
rect 5521 568 5532 602
rect 5566 568 5577 602
rect 5521 534 5577 568
rect 5521 500 5532 534
rect 5566 500 5577 534
rect 5521 466 5577 500
rect 5521 432 5532 466
rect 5566 432 5577 466
rect 5521 398 5577 432
rect 5521 364 5532 398
rect 5566 364 5577 398
rect 5521 330 5577 364
rect 5521 296 5532 330
rect 5566 296 5577 330
rect 5521 262 5577 296
rect 5521 228 5532 262
rect 5566 228 5577 262
rect 5521 194 5577 228
rect 5521 160 5532 194
rect 5566 160 5577 194
rect 5521 148 5577 160
rect 5627 1078 5680 1148
rect 5627 1044 5638 1078
rect 5672 1044 5680 1078
rect 5627 1010 5680 1044
rect 5627 976 5638 1010
rect 5672 976 5680 1010
rect 5627 942 5680 976
rect 5627 908 5638 942
rect 5672 908 5680 942
rect 5627 874 5680 908
rect 5627 840 5638 874
rect 5672 840 5680 874
rect 5627 806 5680 840
rect 5627 772 5638 806
rect 5672 772 5680 806
rect 5627 738 5680 772
rect 5627 704 5638 738
rect 5672 704 5680 738
rect 5627 670 5680 704
rect 5627 636 5638 670
rect 5672 636 5680 670
rect 5627 602 5680 636
rect 5627 568 5638 602
rect 5672 568 5680 602
rect 5627 534 5680 568
rect 5627 500 5638 534
rect 5672 500 5680 534
rect 5627 466 5680 500
rect 5627 432 5638 466
rect 5672 432 5680 466
rect 5627 398 5680 432
rect 5627 364 5638 398
rect 5672 364 5680 398
rect 5627 330 5680 364
rect 5627 296 5638 330
rect 5672 296 5680 330
rect 5627 262 5680 296
rect 5627 228 5638 262
rect 5672 228 5680 262
rect 5627 194 5680 228
rect 5627 160 5638 194
rect 5672 160 5680 194
rect 5627 148 5680 160
<< mvndiff >>
rect -109 2760 -56 2838
rect -109 2726 -101 2760
rect -67 2726 -56 2760
rect -109 2692 -56 2726
rect -109 2658 -101 2692
rect -67 2658 -56 2692
rect -109 2624 -56 2658
rect -109 2590 -101 2624
rect -67 2590 -56 2624
rect -109 2556 -56 2590
rect -109 2522 -101 2556
rect -67 2522 -56 2556
rect -109 2488 -56 2522
rect -109 2454 -101 2488
rect -67 2454 -56 2488
rect -109 2420 -56 2454
rect -109 2386 -101 2420
rect -67 2386 -56 2420
rect -109 2352 -56 2386
rect -109 2318 -101 2352
rect -67 2318 -56 2352
rect -109 2284 -56 2318
rect -109 2250 -101 2284
rect -67 2250 -56 2284
rect -109 2238 -56 2250
rect 44 2760 97 2838
rect 44 2726 55 2760
rect 89 2726 97 2760
rect 44 2692 97 2726
rect 44 2658 55 2692
rect 89 2658 97 2692
rect 44 2624 97 2658
rect 44 2590 55 2624
rect 89 2590 97 2624
rect 44 2556 97 2590
rect 44 2522 55 2556
rect 89 2522 97 2556
rect 44 2488 97 2522
rect 44 2454 55 2488
rect 89 2454 97 2488
rect 44 2420 97 2454
rect 44 2386 55 2420
rect 89 2386 97 2420
rect 44 2352 97 2386
rect 44 2318 55 2352
rect 89 2318 97 2352
rect 44 2284 97 2318
rect 44 2250 55 2284
rect 89 2250 97 2284
rect 44 2238 97 2250
rect 12218 2660 14218 2668
rect 12218 2626 12268 2660
rect 12302 2626 12336 2660
rect 12370 2626 12404 2660
rect 12438 2626 12472 2660
rect 12506 2626 12540 2660
rect 12574 2626 12608 2660
rect 12642 2626 12676 2660
rect 12710 2626 12744 2660
rect 12778 2626 12812 2660
rect 12846 2626 12880 2660
rect 12914 2626 12948 2660
rect 12982 2626 13016 2660
rect 13050 2626 13084 2660
rect 13118 2626 13152 2660
rect 13186 2626 13220 2660
rect 13254 2626 13288 2660
rect 13322 2626 13356 2660
rect 13390 2626 13424 2660
rect 13458 2626 13492 2660
rect 13526 2626 13560 2660
rect 13594 2626 13628 2660
rect 13662 2626 13696 2660
rect 13730 2626 13764 2660
rect 13798 2626 13832 2660
rect 13866 2626 13900 2660
rect 13934 2626 13968 2660
rect 14002 2626 14036 2660
rect 14070 2626 14104 2660
rect 14138 2626 14172 2660
rect 14206 2626 14218 2660
rect 12218 2615 14218 2626
rect 14862 2660 16862 2668
rect 14862 2626 14912 2660
rect 14946 2626 14980 2660
rect 15014 2626 15048 2660
rect 15082 2626 15116 2660
rect 15150 2626 15184 2660
rect 15218 2626 15252 2660
rect 15286 2626 15320 2660
rect 15354 2626 15388 2660
rect 15422 2626 15456 2660
rect 15490 2626 15524 2660
rect 15558 2626 15592 2660
rect 15626 2626 15660 2660
rect 15694 2626 15728 2660
rect 15762 2626 15796 2660
rect 15830 2626 15864 2660
rect 15898 2626 15932 2660
rect 15966 2626 16000 2660
rect 16034 2626 16068 2660
rect 16102 2626 16136 2660
rect 16170 2626 16204 2660
rect 16238 2626 16272 2660
rect 16306 2626 16340 2660
rect 16374 2626 16408 2660
rect 16442 2626 16476 2660
rect 16510 2626 16544 2660
rect 16578 2626 16612 2660
rect 16646 2626 16680 2660
rect 16714 2626 16748 2660
rect 16782 2626 16816 2660
rect 16850 2626 16862 2660
rect 14862 2615 16862 2626
rect 12218 2424 14218 2435
rect 12218 2390 12268 2424
rect 12302 2390 12336 2424
rect 12370 2390 12404 2424
rect 12438 2390 12472 2424
rect 12506 2390 12540 2424
rect 12574 2390 12608 2424
rect 12642 2390 12676 2424
rect 12710 2390 12744 2424
rect 12778 2390 12812 2424
rect 12846 2390 12880 2424
rect 12914 2390 12948 2424
rect 12982 2390 13016 2424
rect 13050 2390 13084 2424
rect 13118 2390 13152 2424
rect 13186 2390 13220 2424
rect 13254 2390 13288 2424
rect 13322 2390 13356 2424
rect 13390 2390 13424 2424
rect 13458 2390 13492 2424
rect 13526 2390 13560 2424
rect 13594 2390 13628 2424
rect 13662 2390 13696 2424
rect 13730 2390 13764 2424
rect 13798 2390 13832 2424
rect 13866 2390 13900 2424
rect 13934 2390 13968 2424
rect 14002 2390 14036 2424
rect 14070 2390 14104 2424
rect 14138 2390 14172 2424
rect 14206 2390 14218 2424
rect 12218 2379 14218 2390
rect 12218 2188 14218 2199
rect 12218 2154 12268 2188
rect 12302 2154 12336 2188
rect 12370 2154 12404 2188
rect 12438 2154 12472 2188
rect 12506 2154 12540 2188
rect 12574 2154 12608 2188
rect 12642 2154 12676 2188
rect 12710 2154 12744 2188
rect 12778 2154 12812 2188
rect 12846 2154 12880 2188
rect 12914 2154 12948 2188
rect 12982 2154 13016 2188
rect 13050 2154 13084 2188
rect 13118 2154 13152 2188
rect 13186 2154 13220 2188
rect 13254 2154 13288 2188
rect 13322 2154 13356 2188
rect 13390 2154 13424 2188
rect 13458 2154 13492 2188
rect 13526 2154 13560 2188
rect 13594 2154 13628 2188
rect 13662 2154 13696 2188
rect 13730 2154 13764 2188
rect 13798 2154 13832 2188
rect 13866 2154 13900 2188
rect 13934 2154 13968 2188
rect 14002 2154 14036 2188
rect 14070 2154 14104 2188
rect 14138 2154 14172 2188
rect 14206 2154 14218 2188
rect 12218 2143 14218 2154
rect 12218 1952 14218 1963
rect 12218 1918 12268 1952
rect 12302 1918 12336 1952
rect 12370 1918 12404 1952
rect 12438 1918 12472 1952
rect 12506 1918 12540 1952
rect 12574 1918 12608 1952
rect 12642 1918 12676 1952
rect 12710 1918 12744 1952
rect 12778 1918 12812 1952
rect 12846 1918 12880 1952
rect 12914 1918 12948 1952
rect 12982 1918 13016 1952
rect 13050 1918 13084 1952
rect 13118 1918 13152 1952
rect 13186 1918 13220 1952
rect 13254 1918 13288 1952
rect 13322 1918 13356 1952
rect 13390 1918 13424 1952
rect 13458 1918 13492 1952
rect 13526 1918 13560 1952
rect 13594 1918 13628 1952
rect 13662 1918 13696 1952
rect 13730 1918 13764 1952
rect 13798 1918 13832 1952
rect 13866 1918 13900 1952
rect 13934 1918 13968 1952
rect 14002 1918 14036 1952
rect 14070 1918 14104 1952
rect 14138 1918 14172 1952
rect 14206 1918 14218 1952
rect 12218 1910 14218 1918
rect 14862 2424 16862 2435
rect 14862 2390 14912 2424
rect 14946 2390 14980 2424
rect 15014 2390 15048 2424
rect 15082 2390 15116 2424
rect 15150 2390 15184 2424
rect 15218 2390 15252 2424
rect 15286 2390 15320 2424
rect 15354 2390 15388 2424
rect 15422 2390 15456 2424
rect 15490 2390 15524 2424
rect 15558 2390 15592 2424
rect 15626 2390 15660 2424
rect 15694 2390 15728 2424
rect 15762 2390 15796 2424
rect 15830 2390 15864 2424
rect 15898 2390 15932 2424
rect 15966 2390 16000 2424
rect 16034 2390 16068 2424
rect 16102 2390 16136 2424
rect 16170 2390 16204 2424
rect 16238 2390 16272 2424
rect 16306 2390 16340 2424
rect 16374 2390 16408 2424
rect 16442 2390 16476 2424
rect 16510 2390 16544 2424
rect 16578 2390 16612 2424
rect 16646 2390 16680 2424
rect 16714 2390 16748 2424
rect 16782 2390 16816 2424
rect 16850 2390 16862 2424
rect 14862 2379 16862 2390
rect 14862 2188 16862 2199
rect 14862 2154 14912 2188
rect 14946 2154 14980 2188
rect 15014 2154 15048 2188
rect 15082 2154 15116 2188
rect 15150 2154 15184 2188
rect 15218 2154 15252 2188
rect 15286 2154 15320 2188
rect 15354 2154 15388 2188
rect 15422 2154 15456 2188
rect 15490 2154 15524 2188
rect 15558 2154 15592 2188
rect 15626 2154 15660 2188
rect 15694 2154 15728 2188
rect 15762 2154 15796 2188
rect 15830 2154 15864 2188
rect 15898 2154 15932 2188
rect 15966 2154 16000 2188
rect 16034 2154 16068 2188
rect 16102 2154 16136 2188
rect 16170 2154 16204 2188
rect 16238 2154 16272 2188
rect 16306 2154 16340 2188
rect 16374 2154 16408 2188
rect 16442 2154 16476 2188
rect 16510 2154 16544 2188
rect 16578 2154 16612 2188
rect 16646 2154 16680 2188
rect 16714 2154 16748 2188
rect 16782 2154 16816 2188
rect 16850 2154 16862 2188
rect 14862 2143 16862 2154
rect 14862 1952 16862 1963
rect 14862 1918 14912 1952
rect 14946 1918 14980 1952
rect 15014 1918 15048 1952
rect 15082 1918 15116 1952
rect 15150 1918 15184 1952
rect 15218 1918 15252 1952
rect 15286 1918 15320 1952
rect 15354 1918 15388 1952
rect 15422 1918 15456 1952
rect 15490 1918 15524 1952
rect 15558 1918 15592 1952
rect 15626 1918 15660 1952
rect 15694 1918 15728 1952
rect 15762 1918 15796 1952
rect 15830 1918 15864 1952
rect 15898 1918 15932 1952
rect 15966 1918 16000 1952
rect 16034 1918 16068 1952
rect 16102 1918 16136 1952
rect 16170 1918 16204 1952
rect 16238 1918 16272 1952
rect 16306 1918 16340 1952
rect 16374 1918 16408 1952
rect 16442 1918 16476 1952
rect 16510 1918 16544 1952
rect 16578 1918 16612 1952
rect 16646 1918 16680 1952
rect 16714 1918 16748 1952
rect 16782 1918 16816 1952
rect 16850 1918 16862 1952
rect 14862 1910 16862 1918
rect 5892 1130 5945 1148
rect 5892 1096 5900 1130
rect 5934 1096 5945 1130
rect 5892 1062 5945 1096
rect 5892 1028 5900 1062
rect 5934 1028 5945 1062
rect 5892 994 5945 1028
rect 5892 960 5900 994
rect 5934 960 5945 994
rect 5892 948 5945 960
rect 6105 1130 6161 1148
rect 6105 1096 6116 1130
rect 6150 1096 6161 1130
rect 6105 1062 6161 1096
rect 6105 1028 6116 1062
rect 6150 1028 6161 1062
rect 6105 994 6161 1028
rect 6105 960 6116 994
rect 6150 960 6161 994
rect 6105 948 6161 960
rect 6321 1130 6377 1148
rect 6321 1096 6332 1130
rect 6366 1096 6377 1130
rect 6321 1062 6377 1096
rect 6321 1028 6332 1062
rect 6366 1028 6377 1062
rect 6321 994 6377 1028
rect 6321 960 6332 994
rect 6366 960 6377 994
rect 6321 948 6377 960
rect 6537 1130 6590 1148
rect 6537 1096 6548 1130
rect 6582 1096 6590 1130
rect 6537 1062 6590 1096
rect 6537 1028 6548 1062
rect 6582 1028 6590 1062
rect 6537 994 6590 1028
rect 6537 960 6548 994
rect 6582 960 6590 994
rect 6537 948 6590 960
rect 6650 1070 6703 1148
rect 6650 1036 6658 1070
rect 6692 1036 6703 1070
rect 6650 1002 6703 1036
rect 6650 968 6658 1002
rect 6692 968 6703 1002
rect 6650 934 6703 968
rect 6650 900 6658 934
rect 6692 900 6703 934
rect 6650 866 6703 900
rect 6650 832 6658 866
rect 6692 832 6703 866
rect 5892 800 5945 818
rect 5892 766 5900 800
rect 5934 766 5945 800
rect 5892 732 5945 766
rect 5892 698 5900 732
rect 5934 698 5945 732
rect 5892 664 5945 698
rect 5892 630 5900 664
rect 5934 630 5945 664
rect 5892 618 5945 630
rect 6105 800 6161 818
rect 6105 766 6116 800
rect 6150 766 6161 800
rect 6105 732 6161 766
rect 6105 698 6116 732
rect 6150 698 6161 732
rect 6105 664 6161 698
rect 6105 630 6116 664
rect 6150 630 6161 664
rect 6105 618 6161 630
rect 6321 800 6377 818
rect 6321 766 6332 800
rect 6366 766 6377 800
rect 6321 732 6377 766
rect 6321 698 6332 732
rect 6366 698 6377 732
rect 6321 664 6377 698
rect 6321 630 6332 664
rect 6366 630 6377 664
rect 6321 618 6377 630
rect 6537 800 6590 818
rect 6537 766 6548 800
rect 6582 766 6590 800
rect 6537 732 6590 766
rect 6537 698 6548 732
rect 6582 698 6590 732
rect 6537 664 6590 698
rect 6537 630 6548 664
rect 6582 630 6590 664
rect 6537 618 6590 630
rect 6650 798 6703 832
rect 6650 764 6658 798
rect 6692 764 6703 798
rect 6650 730 6703 764
rect 6650 696 6658 730
rect 6692 696 6703 730
rect 6650 662 6703 696
rect 6650 628 6658 662
rect 6692 628 6703 662
rect 6650 594 6703 628
rect 6650 560 6658 594
rect 6692 560 6703 594
rect 6650 548 6703 560
rect 6803 1070 6859 1148
rect 6803 1036 6814 1070
rect 6848 1036 6859 1070
rect 6803 1002 6859 1036
rect 6803 968 6814 1002
rect 6848 968 6859 1002
rect 6803 934 6859 968
rect 6803 900 6814 934
rect 6848 900 6859 934
rect 6803 866 6859 900
rect 6803 832 6814 866
rect 6848 832 6859 866
rect 6803 798 6859 832
rect 6803 764 6814 798
rect 6848 764 6859 798
rect 6803 730 6859 764
rect 6803 696 6814 730
rect 6848 696 6859 730
rect 6803 662 6859 696
rect 6803 628 6814 662
rect 6848 628 6859 662
rect 6803 594 6859 628
rect 6803 560 6814 594
rect 6848 560 6859 594
rect 6803 548 6859 560
rect 6959 1070 7015 1148
rect 6959 1036 6970 1070
rect 7004 1036 7015 1070
rect 6959 1002 7015 1036
rect 6959 968 6970 1002
rect 7004 968 7015 1002
rect 6959 934 7015 968
rect 6959 900 6970 934
rect 7004 900 7015 934
rect 6959 866 7015 900
rect 6959 832 6970 866
rect 7004 832 7015 866
rect 6959 798 7015 832
rect 6959 764 6970 798
rect 7004 764 7015 798
rect 6959 730 7015 764
rect 6959 696 6970 730
rect 7004 696 7015 730
rect 6959 662 7015 696
rect 6959 628 6970 662
rect 7004 628 7015 662
rect 6959 594 7015 628
rect 6959 560 6970 594
rect 7004 560 7015 594
rect 6959 548 7015 560
rect 7115 1070 7168 1148
rect 7115 1036 7126 1070
rect 7160 1036 7168 1070
rect 7115 1002 7168 1036
rect 7115 968 7126 1002
rect 7160 968 7168 1002
rect 7115 934 7168 968
rect 7115 900 7126 934
rect 7160 900 7168 934
rect 7115 866 7168 900
rect 7115 832 7126 866
rect 7160 832 7168 866
rect 7115 798 7168 832
rect 7115 764 7126 798
rect 7160 764 7168 798
rect 7115 730 7168 764
rect 7115 696 7126 730
rect 7160 696 7168 730
rect 7115 662 7168 696
rect 7115 628 7126 662
rect 7160 628 7168 662
rect 7115 594 7168 628
rect 7115 560 7126 594
rect 7160 560 7168 594
rect 7115 548 7168 560
rect 7228 1078 7281 1148
rect 7228 1044 7236 1078
rect 7270 1044 7281 1078
rect 7228 1010 7281 1044
rect 7228 976 7236 1010
rect 7270 976 7281 1010
rect 7228 942 7281 976
rect 7228 908 7236 942
rect 7270 908 7281 942
rect 7228 874 7281 908
rect 7228 840 7236 874
rect 7270 840 7281 874
rect 7228 806 7281 840
rect 7228 772 7236 806
rect 7270 772 7281 806
rect 7228 738 7281 772
rect 7228 704 7236 738
rect 7270 704 7281 738
rect 7228 670 7281 704
rect 7228 636 7236 670
rect 7270 636 7281 670
rect 7228 602 7281 636
rect 7228 568 7236 602
rect 7270 568 7281 602
rect 7228 534 7281 568
rect 7228 500 7236 534
rect 7270 500 7281 534
rect 7228 466 7281 500
rect 5892 434 5945 446
rect 5892 400 5900 434
rect 5934 400 5945 434
rect 5892 366 5945 400
rect 5892 332 5900 366
rect 5934 332 5945 366
rect 5892 298 5945 332
rect 5892 264 5900 298
rect 5934 264 5945 298
rect 5892 246 5945 264
rect 6105 434 6161 446
rect 6105 400 6116 434
rect 6150 400 6161 434
rect 6105 366 6161 400
rect 6105 332 6116 366
rect 6150 332 6161 366
rect 6105 298 6161 332
rect 6105 264 6116 298
rect 6150 264 6161 298
rect 6105 246 6161 264
rect 6321 434 6377 446
rect 6321 400 6332 434
rect 6366 400 6377 434
rect 6321 366 6377 400
rect 6321 332 6332 366
rect 6366 332 6377 366
rect 6321 298 6377 332
rect 6321 264 6332 298
rect 6366 264 6377 298
rect 6321 246 6377 264
rect 6537 434 6590 446
rect 6537 400 6548 434
rect 6582 400 6590 434
rect 6537 366 6590 400
rect 6537 332 6548 366
rect 6582 332 6590 366
rect 6537 298 6590 332
rect 6537 264 6548 298
rect 6582 264 6590 298
rect 6537 246 6590 264
rect 7228 432 7236 466
rect 7270 432 7281 466
rect 7228 398 7281 432
rect 7228 364 7236 398
rect 7270 364 7281 398
rect 7228 330 7281 364
rect 7228 296 7236 330
rect 7270 296 7281 330
rect 7228 262 7281 296
rect 7228 228 7236 262
rect 7270 228 7281 262
rect 7228 194 7281 228
rect 7228 160 7236 194
rect 7270 160 7281 194
rect 7228 148 7281 160
rect 7381 1078 7434 1148
rect 7381 1044 7392 1078
rect 7426 1044 7434 1078
rect 7381 1010 7434 1044
rect 7381 976 7392 1010
rect 7426 976 7434 1010
rect 7381 942 7434 976
rect 7381 908 7392 942
rect 7426 908 7434 942
rect 7381 874 7434 908
rect 7381 840 7392 874
rect 7426 840 7434 874
rect 7381 806 7434 840
rect 7381 772 7392 806
rect 7426 772 7434 806
rect 7381 738 7434 772
rect 7381 704 7392 738
rect 7426 704 7434 738
rect 7381 670 7434 704
rect 7381 636 7392 670
rect 7426 636 7434 670
rect 7381 602 7434 636
rect 7381 568 7392 602
rect 7426 568 7434 602
rect 7381 534 7434 568
rect 7381 500 7392 534
rect 7426 500 7434 534
rect 7381 466 7434 500
rect 7381 432 7392 466
rect 7426 432 7434 466
rect 7381 398 7434 432
rect 7381 364 7392 398
rect 7426 364 7434 398
rect 7381 330 7434 364
rect 7381 296 7392 330
rect 7426 296 7434 330
rect 7381 262 7434 296
rect 7381 228 7392 262
rect 7426 228 7434 262
rect 7381 194 7434 228
rect 7381 160 7392 194
rect 7426 160 7434 194
rect 7381 148 7434 160
rect 7494 1078 7547 1148
rect 7494 1044 7502 1078
rect 7536 1044 7547 1078
rect 7494 1010 7547 1044
rect 7494 976 7502 1010
rect 7536 976 7547 1010
rect 7494 942 7547 976
rect 7494 908 7502 942
rect 7536 908 7547 942
rect 7494 874 7547 908
rect 7494 840 7502 874
rect 7536 840 7547 874
rect 7494 806 7547 840
rect 7494 772 7502 806
rect 7536 772 7547 806
rect 7494 738 7547 772
rect 7494 704 7502 738
rect 7536 704 7547 738
rect 7494 670 7547 704
rect 7494 636 7502 670
rect 7536 636 7547 670
rect 7494 602 7547 636
rect 7494 568 7502 602
rect 7536 568 7547 602
rect 7494 534 7547 568
rect 7494 500 7502 534
rect 7536 500 7547 534
rect 7494 466 7547 500
rect 7494 432 7502 466
rect 7536 432 7547 466
rect 7494 398 7547 432
rect 7494 364 7502 398
rect 7536 364 7547 398
rect 7494 330 7547 364
rect 7494 296 7502 330
rect 7536 296 7547 330
rect 7494 262 7547 296
rect 7494 228 7502 262
rect 7536 228 7547 262
rect 7494 194 7547 228
rect 7494 160 7502 194
rect 7536 160 7547 194
rect 7494 148 7547 160
rect 7707 1078 7763 1148
rect 7707 1044 7718 1078
rect 7752 1044 7763 1078
rect 7707 1010 7763 1044
rect 7707 976 7718 1010
rect 7752 976 7763 1010
rect 7707 942 7763 976
rect 7707 908 7718 942
rect 7752 908 7763 942
rect 7707 874 7763 908
rect 7707 840 7718 874
rect 7752 840 7763 874
rect 7707 806 7763 840
rect 7707 772 7718 806
rect 7752 772 7763 806
rect 7707 738 7763 772
rect 7707 704 7718 738
rect 7752 704 7763 738
rect 7707 670 7763 704
rect 7707 636 7718 670
rect 7752 636 7763 670
rect 7707 602 7763 636
rect 7707 568 7718 602
rect 7752 568 7763 602
rect 7707 534 7763 568
rect 7707 500 7718 534
rect 7752 500 7763 534
rect 7707 466 7763 500
rect 7707 432 7718 466
rect 7752 432 7763 466
rect 7707 398 7763 432
rect 7707 364 7718 398
rect 7752 364 7763 398
rect 7707 330 7763 364
rect 7707 296 7718 330
rect 7752 296 7763 330
rect 7707 262 7763 296
rect 7707 228 7718 262
rect 7752 228 7763 262
rect 7707 194 7763 228
rect 7707 160 7718 194
rect 7752 160 7763 194
rect 7707 148 7763 160
rect 7923 1078 7979 1148
rect 7923 1044 7934 1078
rect 7968 1044 7979 1078
rect 7923 1010 7979 1044
rect 7923 976 7934 1010
rect 7968 976 7979 1010
rect 7923 942 7979 976
rect 7923 908 7934 942
rect 7968 908 7979 942
rect 7923 874 7979 908
rect 7923 840 7934 874
rect 7968 840 7979 874
rect 7923 806 7979 840
rect 7923 772 7934 806
rect 7968 772 7979 806
rect 7923 738 7979 772
rect 7923 704 7934 738
rect 7968 704 7979 738
rect 7923 670 7979 704
rect 7923 636 7934 670
rect 7968 636 7979 670
rect 7923 602 7979 636
rect 7923 568 7934 602
rect 7968 568 7979 602
rect 7923 534 7979 568
rect 7923 500 7934 534
rect 7968 500 7979 534
rect 7923 466 7979 500
rect 7923 432 7934 466
rect 7968 432 7979 466
rect 7923 398 7979 432
rect 7923 364 7934 398
rect 7968 364 7979 398
rect 7923 330 7979 364
rect 7923 296 7934 330
rect 7968 296 7979 330
rect 7923 262 7979 296
rect 7923 228 7934 262
rect 7968 228 7979 262
rect 7923 194 7979 228
rect 7923 160 7934 194
rect 7968 160 7979 194
rect 7923 148 7979 160
rect 8139 1078 8195 1148
rect 8139 1044 8150 1078
rect 8184 1044 8195 1078
rect 8139 1010 8195 1044
rect 8139 976 8150 1010
rect 8184 976 8195 1010
rect 8139 942 8195 976
rect 8139 908 8150 942
rect 8184 908 8195 942
rect 8139 874 8195 908
rect 8139 840 8150 874
rect 8184 840 8195 874
rect 8139 806 8195 840
rect 8139 772 8150 806
rect 8184 772 8195 806
rect 8139 738 8195 772
rect 8139 704 8150 738
rect 8184 704 8195 738
rect 8139 670 8195 704
rect 8139 636 8150 670
rect 8184 636 8195 670
rect 8139 602 8195 636
rect 8139 568 8150 602
rect 8184 568 8195 602
rect 8139 534 8195 568
rect 8139 500 8150 534
rect 8184 500 8195 534
rect 8139 466 8195 500
rect 8139 432 8150 466
rect 8184 432 8195 466
rect 8139 398 8195 432
rect 8139 364 8150 398
rect 8184 364 8195 398
rect 8139 330 8195 364
rect 8139 296 8150 330
rect 8184 296 8195 330
rect 8139 262 8195 296
rect 8139 228 8150 262
rect 8184 228 8195 262
rect 8139 194 8195 228
rect 8139 160 8150 194
rect 8184 160 8195 194
rect 8139 148 8195 160
rect 8355 1078 8411 1148
rect 8355 1044 8366 1078
rect 8400 1044 8411 1078
rect 8355 1010 8411 1044
rect 8355 976 8366 1010
rect 8400 976 8411 1010
rect 8355 942 8411 976
rect 8355 908 8366 942
rect 8400 908 8411 942
rect 8355 874 8411 908
rect 8355 840 8366 874
rect 8400 840 8411 874
rect 8355 806 8411 840
rect 8355 772 8366 806
rect 8400 772 8411 806
rect 8355 738 8411 772
rect 8355 704 8366 738
rect 8400 704 8411 738
rect 8355 670 8411 704
rect 8355 636 8366 670
rect 8400 636 8411 670
rect 8355 602 8411 636
rect 8355 568 8366 602
rect 8400 568 8411 602
rect 8355 534 8411 568
rect 8355 500 8366 534
rect 8400 500 8411 534
rect 8355 466 8411 500
rect 8355 432 8366 466
rect 8400 432 8411 466
rect 8355 398 8411 432
rect 8355 364 8366 398
rect 8400 364 8411 398
rect 8355 330 8411 364
rect 8355 296 8366 330
rect 8400 296 8411 330
rect 8355 262 8411 296
rect 8355 228 8366 262
rect 8400 228 8411 262
rect 8355 194 8411 228
rect 8355 160 8366 194
rect 8400 160 8411 194
rect 8355 148 8411 160
rect 8571 1078 8627 1148
rect 8571 1044 8582 1078
rect 8616 1044 8627 1078
rect 8571 1010 8627 1044
rect 8571 976 8582 1010
rect 8616 976 8627 1010
rect 8571 942 8627 976
rect 8571 908 8582 942
rect 8616 908 8627 942
rect 8571 874 8627 908
rect 8571 840 8582 874
rect 8616 840 8627 874
rect 8571 806 8627 840
rect 8571 772 8582 806
rect 8616 772 8627 806
rect 8571 738 8627 772
rect 8571 704 8582 738
rect 8616 704 8627 738
rect 8571 670 8627 704
rect 8571 636 8582 670
rect 8616 636 8627 670
rect 8571 602 8627 636
rect 8571 568 8582 602
rect 8616 568 8627 602
rect 8571 534 8627 568
rect 8571 500 8582 534
rect 8616 500 8627 534
rect 8571 466 8627 500
rect 8571 432 8582 466
rect 8616 432 8627 466
rect 8571 398 8627 432
rect 8571 364 8582 398
rect 8616 364 8627 398
rect 8571 330 8627 364
rect 8571 296 8582 330
rect 8616 296 8627 330
rect 8571 262 8627 296
rect 8571 228 8582 262
rect 8616 228 8627 262
rect 8571 194 8627 228
rect 8571 160 8582 194
rect 8616 160 8627 194
rect 8571 148 8627 160
rect 8787 1078 8843 1148
rect 8787 1044 8798 1078
rect 8832 1044 8843 1078
rect 8787 1010 8843 1044
rect 8787 976 8798 1010
rect 8832 976 8843 1010
rect 8787 942 8843 976
rect 8787 908 8798 942
rect 8832 908 8843 942
rect 8787 874 8843 908
rect 8787 840 8798 874
rect 8832 840 8843 874
rect 8787 806 8843 840
rect 8787 772 8798 806
rect 8832 772 8843 806
rect 8787 738 8843 772
rect 8787 704 8798 738
rect 8832 704 8843 738
rect 8787 670 8843 704
rect 8787 636 8798 670
rect 8832 636 8843 670
rect 8787 602 8843 636
rect 8787 568 8798 602
rect 8832 568 8843 602
rect 8787 534 8843 568
rect 8787 500 8798 534
rect 8832 500 8843 534
rect 8787 466 8843 500
rect 8787 432 8798 466
rect 8832 432 8843 466
rect 8787 398 8843 432
rect 8787 364 8798 398
rect 8832 364 8843 398
rect 8787 330 8843 364
rect 8787 296 8798 330
rect 8832 296 8843 330
rect 8787 262 8843 296
rect 8787 228 8798 262
rect 8832 228 8843 262
rect 8787 194 8843 228
rect 8787 160 8798 194
rect 8832 160 8843 194
rect 8787 148 8843 160
rect 9003 1078 9059 1148
rect 9003 1044 9014 1078
rect 9048 1044 9059 1078
rect 9003 1010 9059 1044
rect 9003 976 9014 1010
rect 9048 976 9059 1010
rect 9003 942 9059 976
rect 9003 908 9014 942
rect 9048 908 9059 942
rect 9003 874 9059 908
rect 9003 840 9014 874
rect 9048 840 9059 874
rect 9003 806 9059 840
rect 9003 772 9014 806
rect 9048 772 9059 806
rect 9003 738 9059 772
rect 9003 704 9014 738
rect 9048 704 9059 738
rect 9003 670 9059 704
rect 9003 636 9014 670
rect 9048 636 9059 670
rect 9003 602 9059 636
rect 9003 568 9014 602
rect 9048 568 9059 602
rect 9003 534 9059 568
rect 9003 500 9014 534
rect 9048 500 9059 534
rect 9003 466 9059 500
rect 9003 432 9014 466
rect 9048 432 9059 466
rect 9003 398 9059 432
rect 9003 364 9014 398
rect 9048 364 9059 398
rect 9003 330 9059 364
rect 9003 296 9014 330
rect 9048 296 9059 330
rect 9003 262 9059 296
rect 9003 228 9014 262
rect 9048 228 9059 262
rect 9003 194 9059 228
rect 9003 160 9014 194
rect 9048 160 9059 194
rect 9003 148 9059 160
rect 9219 1078 9275 1148
rect 9219 1044 9230 1078
rect 9264 1044 9275 1078
rect 9219 1010 9275 1044
rect 9219 976 9230 1010
rect 9264 976 9275 1010
rect 9219 942 9275 976
rect 9219 908 9230 942
rect 9264 908 9275 942
rect 9219 874 9275 908
rect 9219 840 9230 874
rect 9264 840 9275 874
rect 9219 806 9275 840
rect 9219 772 9230 806
rect 9264 772 9275 806
rect 9219 738 9275 772
rect 9219 704 9230 738
rect 9264 704 9275 738
rect 9219 670 9275 704
rect 9219 636 9230 670
rect 9264 636 9275 670
rect 9219 602 9275 636
rect 9219 568 9230 602
rect 9264 568 9275 602
rect 9219 534 9275 568
rect 9219 500 9230 534
rect 9264 500 9275 534
rect 9219 466 9275 500
rect 9219 432 9230 466
rect 9264 432 9275 466
rect 9219 398 9275 432
rect 9219 364 9230 398
rect 9264 364 9275 398
rect 9219 330 9275 364
rect 9219 296 9230 330
rect 9264 296 9275 330
rect 9219 262 9275 296
rect 9219 228 9230 262
rect 9264 228 9275 262
rect 9219 194 9275 228
rect 9219 160 9230 194
rect 9264 160 9275 194
rect 9219 148 9275 160
rect 9435 1078 9491 1148
rect 9435 1044 9446 1078
rect 9480 1044 9491 1078
rect 9435 1010 9491 1044
rect 9435 976 9446 1010
rect 9480 976 9491 1010
rect 9435 942 9491 976
rect 9435 908 9446 942
rect 9480 908 9491 942
rect 9435 874 9491 908
rect 9435 840 9446 874
rect 9480 840 9491 874
rect 9435 806 9491 840
rect 9435 772 9446 806
rect 9480 772 9491 806
rect 9435 738 9491 772
rect 9435 704 9446 738
rect 9480 704 9491 738
rect 9435 670 9491 704
rect 9435 636 9446 670
rect 9480 636 9491 670
rect 9435 602 9491 636
rect 9435 568 9446 602
rect 9480 568 9491 602
rect 9435 534 9491 568
rect 9435 500 9446 534
rect 9480 500 9491 534
rect 9435 466 9491 500
rect 9435 432 9446 466
rect 9480 432 9491 466
rect 9435 398 9491 432
rect 9435 364 9446 398
rect 9480 364 9491 398
rect 9435 330 9491 364
rect 9435 296 9446 330
rect 9480 296 9491 330
rect 9435 262 9491 296
rect 9435 228 9446 262
rect 9480 228 9491 262
rect 9435 194 9491 228
rect 9435 160 9446 194
rect 9480 160 9491 194
rect 9435 148 9491 160
rect 9651 1078 9707 1148
rect 9651 1044 9662 1078
rect 9696 1044 9707 1078
rect 9651 1010 9707 1044
rect 9651 976 9662 1010
rect 9696 976 9707 1010
rect 9651 942 9707 976
rect 9651 908 9662 942
rect 9696 908 9707 942
rect 9651 874 9707 908
rect 9651 840 9662 874
rect 9696 840 9707 874
rect 9651 806 9707 840
rect 9651 772 9662 806
rect 9696 772 9707 806
rect 9651 738 9707 772
rect 9651 704 9662 738
rect 9696 704 9707 738
rect 9651 670 9707 704
rect 9651 636 9662 670
rect 9696 636 9707 670
rect 9651 602 9707 636
rect 9651 568 9662 602
rect 9696 568 9707 602
rect 9651 534 9707 568
rect 9651 500 9662 534
rect 9696 500 9707 534
rect 9651 466 9707 500
rect 9651 432 9662 466
rect 9696 432 9707 466
rect 9651 398 9707 432
rect 9651 364 9662 398
rect 9696 364 9707 398
rect 9651 330 9707 364
rect 9651 296 9662 330
rect 9696 296 9707 330
rect 9651 262 9707 296
rect 9651 228 9662 262
rect 9696 228 9707 262
rect 9651 194 9707 228
rect 9651 160 9662 194
rect 9696 160 9707 194
rect 9651 148 9707 160
rect 9867 1078 9923 1148
rect 9867 1044 9878 1078
rect 9912 1044 9923 1078
rect 9867 1010 9923 1044
rect 9867 976 9878 1010
rect 9912 976 9923 1010
rect 9867 942 9923 976
rect 9867 908 9878 942
rect 9912 908 9923 942
rect 9867 874 9923 908
rect 9867 840 9878 874
rect 9912 840 9923 874
rect 9867 806 9923 840
rect 9867 772 9878 806
rect 9912 772 9923 806
rect 9867 738 9923 772
rect 9867 704 9878 738
rect 9912 704 9923 738
rect 9867 670 9923 704
rect 9867 636 9878 670
rect 9912 636 9923 670
rect 9867 602 9923 636
rect 9867 568 9878 602
rect 9912 568 9923 602
rect 9867 534 9923 568
rect 9867 500 9878 534
rect 9912 500 9923 534
rect 9867 466 9923 500
rect 9867 432 9878 466
rect 9912 432 9923 466
rect 9867 398 9923 432
rect 9867 364 9878 398
rect 9912 364 9923 398
rect 9867 330 9923 364
rect 9867 296 9878 330
rect 9912 296 9923 330
rect 9867 262 9923 296
rect 9867 228 9878 262
rect 9912 228 9923 262
rect 9867 194 9923 228
rect 9867 160 9878 194
rect 9912 160 9923 194
rect 9867 148 9923 160
rect 10083 1078 10139 1148
rect 10083 1044 10094 1078
rect 10128 1044 10139 1078
rect 10083 1010 10139 1044
rect 10083 976 10094 1010
rect 10128 976 10139 1010
rect 10083 942 10139 976
rect 10083 908 10094 942
rect 10128 908 10139 942
rect 10083 874 10139 908
rect 10083 840 10094 874
rect 10128 840 10139 874
rect 10083 806 10139 840
rect 10083 772 10094 806
rect 10128 772 10139 806
rect 10083 738 10139 772
rect 10083 704 10094 738
rect 10128 704 10139 738
rect 10083 670 10139 704
rect 10083 636 10094 670
rect 10128 636 10139 670
rect 10083 602 10139 636
rect 10083 568 10094 602
rect 10128 568 10139 602
rect 10083 534 10139 568
rect 10083 500 10094 534
rect 10128 500 10139 534
rect 10083 466 10139 500
rect 10083 432 10094 466
rect 10128 432 10139 466
rect 10083 398 10139 432
rect 10083 364 10094 398
rect 10128 364 10139 398
rect 10083 330 10139 364
rect 10083 296 10094 330
rect 10128 296 10139 330
rect 10083 262 10139 296
rect 10083 228 10094 262
rect 10128 228 10139 262
rect 10083 194 10139 228
rect 10083 160 10094 194
rect 10128 160 10139 194
rect 10083 148 10139 160
rect 10299 1078 10355 1148
rect 10299 1044 10310 1078
rect 10344 1044 10355 1078
rect 10299 1010 10355 1044
rect 10299 976 10310 1010
rect 10344 976 10355 1010
rect 10299 942 10355 976
rect 10299 908 10310 942
rect 10344 908 10355 942
rect 10299 874 10355 908
rect 10299 840 10310 874
rect 10344 840 10355 874
rect 10299 806 10355 840
rect 10299 772 10310 806
rect 10344 772 10355 806
rect 10299 738 10355 772
rect 10299 704 10310 738
rect 10344 704 10355 738
rect 10299 670 10355 704
rect 10299 636 10310 670
rect 10344 636 10355 670
rect 10299 602 10355 636
rect 10299 568 10310 602
rect 10344 568 10355 602
rect 10299 534 10355 568
rect 10299 500 10310 534
rect 10344 500 10355 534
rect 10299 466 10355 500
rect 10299 432 10310 466
rect 10344 432 10355 466
rect 10299 398 10355 432
rect 10299 364 10310 398
rect 10344 364 10355 398
rect 10299 330 10355 364
rect 10299 296 10310 330
rect 10344 296 10355 330
rect 10299 262 10355 296
rect 10299 228 10310 262
rect 10344 228 10355 262
rect 10299 194 10355 228
rect 10299 160 10310 194
rect 10344 160 10355 194
rect 10299 148 10355 160
rect 10515 1078 10571 1148
rect 10515 1044 10526 1078
rect 10560 1044 10571 1078
rect 10515 1010 10571 1044
rect 10515 976 10526 1010
rect 10560 976 10571 1010
rect 10515 942 10571 976
rect 10515 908 10526 942
rect 10560 908 10571 942
rect 10515 874 10571 908
rect 10515 840 10526 874
rect 10560 840 10571 874
rect 10515 806 10571 840
rect 10515 772 10526 806
rect 10560 772 10571 806
rect 10515 738 10571 772
rect 10515 704 10526 738
rect 10560 704 10571 738
rect 10515 670 10571 704
rect 10515 636 10526 670
rect 10560 636 10571 670
rect 10515 602 10571 636
rect 10515 568 10526 602
rect 10560 568 10571 602
rect 10515 534 10571 568
rect 10515 500 10526 534
rect 10560 500 10571 534
rect 10515 466 10571 500
rect 10515 432 10526 466
rect 10560 432 10571 466
rect 10515 398 10571 432
rect 10515 364 10526 398
rect 10560 364 10571 398
rect 10515 330 10571 364
rect 10515 296 10526 330
rect 10560 296 10571 330
rect 10515 262 10571 296
rect 10515 228 10526 262
rect 10560 228 10571 262
rect 10515 194 10571 228
rect 10515 160 10526 194
rect 10560 160 10571 194
rect 10515 148 10571 160
rect 10731 1078 10787 1148
rect 10731 1044 10742 1078
rect 10776 1044 10787 1078
rect 10731 1010 10787 1044
rect 10731 976 10742 1010
rect 10776 976 10787 1010
rect 10731 942 10787 976
rect 10731 908 10742 942
rect 10776 908 10787 942
rect 10731 874 10787 908
rect 10731 840 10742 874
rect 10776 840 10787 874
rect 10731 806 10787 840
rect 10731 772 10742 806
rect 10776 772 10787 806
rect 10731 738 10787 772
rect 10731 704 10742 738
rect 10776 704 10787 738
rect 10731 670 10787 704
rect 10731 636 10742 670
rect 10776 636 10787 670
rect 10731 602 10787 636
rect 10731 568 10742 602
rect 10776 568 10787 602
rect 10731 534 10787 568
rect 10731 500 10742 534
rect 10776 500 10787 534
rect 10731 466 10787 500
rect 10731 432 10742 466
rect 10776 432 10787 466
rect 10731 398 10787 432
rect 10731 364 10742 398
rect 10776 364 10787 398
rect 10731 330 10787 364
rect 10731 296 10742 330
rect 10776 296 10787 330
rect 10731 262 10787 296
rect 10731 228 10742 262
rect 10776 228 10787 262
rect 10731 194 10787 228
rect 10731 160 10742 194
rect 10776 160 10787 194
rect 10731 148 10787 160
rect 10947 1078 11003 1148
rect 10947 1044 10958 1078
rect 10992 1044 11003 1078
rect 10947 1010 11003 1044
rect 10947 976 10958 1010
rect 10992 976 11003 1010
rect 10947 942 11003 976
rect 10947 908 10958 942
rect 10992 908 11003 942
rect 10947 874 11003 908
rect 10947 840 10958 874
rect 10992 840 11003 874
rect 10947 806 11003 840
rect 10947 772 10958 806
rect 10992 772 11003 806
rect 10947 738 11003 772
rect 10947 704 10958 738
rect 10992 704 11003 738
rect 10947 670 11003 704
rect 10947 636 10958 670
rect 10992 636 11003 670
rect 10947 602 11003 636
rect 10947 568 10958 602
rect 10992 568 11003 602
rect 10947 534 11003 568
rect 10947 500 10958 534
rect 10992 500 11003 534
rect 10947 466 11003 500
rect 10947 432 10958 466
rect 10992 432 11003 466
rect 10947 398 11003 432
rect 10947 364 10958 398
rect 10992 364 11003 398
rect 10947 330 11003 364
rect 10947 296 10958 330
rect 10992 296 11003 330
rect 10947 262 11003 296
rect 10947 228 10958 262
rect 10992 228 11003 262
rect 10947 194 11003 228
rect 10947 160 10958 194
rect 10992 160 11003 194
rect 10947 148 11003 160
rect 11163 1078 11219 1148
rect 11163 1044 11174 1078
rect 11208 1044 11219 1078
rect 11163 1010 11219 1044
rect 11163 976 11174 1010
rect 11208 976 11219 1010
rect 11163 942 11219 976
rect 11163 908 11174 942
rect 11208 908 11219 942
rect 11163 874 11219 908
rect 11163 840 11174 874
rect 11208 840 11219 874
rect 11163 806 11219 840
rect 11163 772 11174 806
rect 11208 772 11219 806
rect 11163 738 11219 772
rect 11163 704 11174 738
rect 11208 704 11219 738
rect 11163 670 11219 704
rect 11163 636 11174 670
rect 11208 636 11219 670
rect 11163 602 11219 636
rect 11163 568 11174 602
rect 11208 568 11219 602
rect 11163 534 11219 568
rect 11163 500 11174 534
rect 11208 500 11219 534
rect 11163 466 11219 500
rect 11163 432 11174 466
rect 11208 432 11219 466
rect 11163 398 11219 432
rect 11163 364 11174 398
rect 11208 364 11219 398
rect 11163 330 11219 364
rect 11163 296 11174 330
rect 11208 296 11219 330
rect 11163 262 11219 296
rect 11163 228 11174 262
rect 11208 228 11219 262
rect 11163 194 11219 228
rect 11163 160 11174 194
rect 11208 160 11219 194
rect 11163 148 11219 160
rect 11379 1078 11435 1148
rect 11379 1044 11390 1078
rect 11424 1044 11435 1078
rect 11379 1010 11435 1044
rect 11379 976 11390 1010
rect 11424 976 11435 1010
rect 11379 942 11435 976
rect 11379 908 11390 942
rect 11424 908 11435 942
rect 11379 874 11435 908
rect 11379 840 11390 874
rect 11424 840 11435 874
rect 11379 806 11435 840
rect 11379 772 11390 806
rect 11424 772 11435 806
rect 11379 738 11435 772
rect 11379 704 11390 738
rect 11424 704 11435 738
rect 11379 670 11435 704
rect 11379 636 11390 670
rect 11424 636 11435 670
rect 11379 602 11435 636
rect 11379 568 11390 602
rect 11424 568 11435 602
rect 11379 534 11435 568
rect 11379 500 11390 534
rect 11424 500 11435 534
rect 11379 466 11435 500
rect 11379 432 11390 466
rect 11424 432 11435 466
rect 11379 398 11435 432
rect 11379 364 11390 398
rect 11424 364 11435 398
rect 11379 330 11435 364
rect 11379 296 11390 330
rect 11424 296 11435 330
rect 11379 262 11435 296
rect 11379 228 11390 262
rect 11424 228 11435 262
rect 11379 194 11435 228
rect 11379 160 11390 194
rect 11424 160 11435 194
rect 11379 148 11435 160
rect 11595 1078 11651 1148
rect 11595 1044 11606 1078
rect 11640 1044 11651 1078
rect 11595 1010 11651 1044
rect 11595 976 11606 1010
rect 11640 976 11651 1010
rect 11595 942 11651 976
rect 11595 908 11606 942
rect 11640 908 11651 942
rect 11595 874 11651 908
rect 11595 840 11606 874
rect 11640 840 11651 874
rect 11595 806 11651 840
rect 11595 772 11606 806
rect 11640 772 11651 806
rect 11595 738 11651 772
rect 11595 704 11606 738
rect 11640 704 11651 738
rect 11595 670 11651 704
rect 11595 636 11606 670
rect 11640 636 11651 670
rect 11595 602 11651 636
rect 11595 568 11606 602
rect 11640 568 11651 602
rect 11595 534 11651 568
rect 11595 500 11606 534
rect 11640 500 11651 534
rect 11595 466 11651 500
rect 11595 432 11606 466
rect 11640 432 11651 466
rect 11595 398 11651 432
rect 11595 364 11606 398
rect 11640 364 11651 398
rect 11595 330 11651 364
rect 11595 296 11606 330
rect 11640 296 11651 330
rect 11595 262 11651 296
rect 11595 228 11606 262
rect 11640 228 11651 262
rect 11595 194 11651 228
rect 11595 160 11606 194
rect 11640 160 11651 194
rect 11595 148 11651 160
rect 11811 1078 11867 1148
rect 11811 1044 11822 1078
rect 11856 1044 11867 1078
rect 11811 1010 11867 1044
rect 11811 976 11822 1010
rect 11856 976 11867 1010
rect 11811 942 11867 976
rect 11811 908 11822 942
rect 11856 908 11867 942
rect 11811 874 11867 908
rect 11811 840 11822 874
rect 11856 840 11867 874
rect 11811 806 11867 840
rect 11811 772 11822 806
rect 11856 772 11867 806
rect 11811 738 11867 772
rect 11811 704 11822 738
rect 11856 704 11867 738
rect 11811 670 11867 704
rect 11811 636 11822 670
rect 11856 636 11867 670
rect 11811 602 11867 636
rect 11811 568 11822 602
rect 11856 568 11867 602
rect 11811 534 11867 568
rect 11811 500 11822 534
rect 11856 500 11867 534
rect 11811 466 11867 500
rect 11811 432 11822 466
rect 11856 432 11867 466
rect 11811 398 11867 432
rect 11811 364 11822 398
rect 11856 364 11867 398
rect 11811 330 11867 364
rect 11811 296 11822 330
rect 11856 296 11867 330
rect 11811 262 11867 296
rect 11811 228 11822 262
rect 11856 228 11867 262
rect 11811 194 11867 228
rect 11811 160 11822 194
rect 11856 160 11867 194
rect 11811 148 11867 160
rect 12027 1078 12083 1148
rect 12027 1044 12038 1078
rect 12072 1044 12083 1078
rect 12027 1010 12083 1044
rect 12027 976 12038 1010
rect 12072 976 12083 1010
rect 12027 942 12083 976
rect 12027 908 12038 942
rect 12072 908 12083 942
rect 12027 874 12083 908
rect 12027 840 12038 874
rect 12072 840 12083 874
rect 12027 806 12083 840
rect 12027 772 12038 806
rect 12072 772 12083 806
rect 12027 738 12083 772
rect 12027 704 12038 738
rect 12072 704 12083 738
rect 12027 670 12083 704
rect 12027 636 12038 670
rect 12072 636 12083 670
rect 12027 602 12083 636
rect 12027 568 12038 602
rect 12072 568 12083 602
rect 12027 534 12083 568
rect 12027 500 12038 534
rect 12072 500 12083 534
rect 12027 466 12083 500
rect 12027 432 12038 466
rect 12072 432 12083 466
rect 12027 398 12083 432
rect 12027 364 12038 398
rect 12072 364 12083 398
rect 12027 330 12083 364
rect 12027 296 12038 330
rect 12072 296 12083 330
rect 12027 262 12083 296
rect 12027 228 12038 262
rect 12072 228 12083 262
rect 12027 194 12083 228
rect 12027 160 12038 194
rect 12072 160 12083 194
rect 12027 148 12083 160
rect 12243 1078 12299 1148
rect 12243 1044 12254 1078
rect 12288 1044 12299 1078
rect 12243 1010 12299 1044
rect 12243 976 12254 1010
rect 12288 976 12299 1010
rect 12243 942 12299 976
rect 12243 908 12254 942
rect 12288 908 12299 942
rect 12243 874 12299 908
rect 12243 840 12254 874
rect 12288 840 12299 874
rect 12243 806 12299 840
rect 12243 772 12254 806
rect 12288 772 12299 806
rect 12243 738 12299 772
rect 12243 704 12254 738
rect 12288 704 12299 738
rect 12243 670 12299 704
rect 12243 636 12254 670
rect 12288 636 12299 670
rect 12243 602 12299 636
rect 12243 568 12254 602
rect 12288 568 12299 602
rect 12243 534 12299 568
rect 12243 500 12254 534
rect 12288 500 12299 534
rect 12243 466 12299 500
rect 12243 432 12254 466
rect 12288 432 12299 466
rect 12243 398 12299 432
rect 12243 364 12254 398
rect 12288 364 12299 398
rect 12243 330 12299 364
rect 12243 296 12254 330
rect 12288 296 12299 330
rect 12243 262 12299 296
rect 12243 228 12254 262
rect 12288 228 12299 262
rect 12243 194 12299 228
rect 12243 160 12254 194
rect 12288 160 12299 194
rect 12243 148 12299 160
rect 12459 1078 12515 1148
rect 12459 1044 12470 1078
rect 12504 1044 12515 1078
rect 12459 1010 12515 1044
rect 12459 976 12470 1010
rect 12504 976 12515 1010
rect 12459 942 12515 976
rect 12459 908 12470 942
rect 12504 908 12515 942
rect 12459 874 12515 908
rect 12459 840 12470 874
rect 12504 840 12515 874
rect 12459 806 12515 840
rect 12459 772 12470 806
rect 12504 772 12515 806
rect 12459 738 12515 772
rect 12459 704 12470 738
rect 12504 704 12515 738
rect 12459 670 12515 704
rect 12459 636 12470 670
rect 12504 636 12515 670
rect 12459 602 12515 636
rect 12459 568 12470 602
rect 12504 568 12515 602
rect 12459 534 12515 568
rect 12459 500 12470 534
rect 12504 500 12515 534
rect 12459 466 12515 500
rect 12459 432 12470 466
rect 12504 432 12515 466
rect 12459 398 12515 432
rect 12459 364 12470 398
rect 12504 364 12515 398
rect 12459 330 12515 364
rect 12459 296 12470 330
rect 12504 296 12515 330
rect 12459 262 12515 296
rect 12459 228 12470 262
rect 12504 228 12515 262
rect 12459 194 12515 228
rect 12459 160 12470 194
rect 12504 160 12515 194
rect 12459 148 12515 160
rect 12675 1078 12731 1148
rect 12675 1044 12686 1078
rect 12720 1044 12731 1078
rect 12675 1010 12731 1044
rect 12675 976 12686 1010
rect 12720 976 12731 1010
rect 12675 942 12731 976
rect 12675 908 12686 942
rect 12720 908 12731 942
rect 12675 874 12731 908
rect 12675 840 12686 874
rect 12720 840 12731 874
rect 12675 806 12731 840
rect 12675 772 12686 806
rect 12720 772 12731 806
rect 12675 738 12731 772
rect 12675 704 12686 738
rect 12720 704 12731 738
rect 12675 670 12731 704
rect 12675 636 12686 670
rect 12720 636 12731 670
rect 12675 602 12731 636
rect 12675 568 12686 602
rect 12720 568 12731 602
rect 12675 534 12731 568
rect 12675 500 12686 534
rect 12720 500 12731 534
rect 12675 466 12731 500
rect 12675 432 12686 466
rect 12720 432 12731 466
rect 12675 398 12731 432
rect 12675 364 12686 398
rect 12720 364 12731 398
rect 12675 330 12731 364
rect 12675 296 12686 330
rect 12720 296 12731 330
rect 12675 262 12731 296
rect 12675 228 12686 262
rect 12720 228 12731 262
rect 12675 194 12731 228
rect 12675 160 12686 194
rect 12720 160 12731 194
rect 12675 148 12731 160
rect 12891 1078 12947 1148
rect 12891 1044 12902 1078
rect 12936 1044 12947 1078
rect 12891 1010 12947 1044
rect 12891 976 12902 1010
rect 12936 976 12947 1010
rect 12891 942 12947 976
rect 12891 908 12902 942
rect 12936 908 12947 942
rect 12891 874 12947 908
rect 12891 840 12902 874
rect 12936 840 12947 874
rect 12891 806 12947 840
rect 12891 772 12902 806
rect 12936 772 12947 806
rect 12891 738 12947 772
rect 12891 704 12902 738
rect 12936 704 12947 738
rect 12891 670 12947 704
rect 12891 636 12902 670
rect 12936 636 12947 670
rect 12891 602 12947 636
rect 12891 568 12902 602
rect 12936 568 12947 602
rect 12891 534 12947 568
rect 12891 500 12902 534
rect 12936 500 12947 534
rect 12891 466 12947 500
rect 12891 432 12902 466
rect 12936 432 12947 466
rect 12891 398 12947 432
rect 12891 364 12902 398
rect 12936 364 12947 398
rect 12891 330 12947 364
rect 12891 296 12902 330
rect 12936 296 12947 330
rect 12891 262 12947 296
rect 12891 228 12902 262
rect 12936 228 12947 262
rect 12891 194 12947 228
rect 12891 160 12902 194
rect 12936 160 12947 194
rect 12891 148 12947 160
rect 13107 1078 13163 1148
rect 13107 1044 13118 1078
rect 13152 1044 13163 1078
rect 13107 1010 13163 1044
rect 13107 976 13118 1010
rect 13152 976 13163 1010
rect 13107 942 13163 976
rect 13107 908 13118 942
rect 13152 908 13163 942
rect 13107 874 13163 908
rect 13107 840 13118 874
rect 13152 840 13163 874
rect 13107 806 13163 840
rect 13107 772 13118 806
rect 13152 772 13163 806
rect 13107 738 13163 772
rect 13107 704 13118 738
rect 13152 704 13163 738
rect 13107 670 13163 704
rect 13107 636 13118 670
rect 13152 636 13163 670
rect 13107 602 13163 636
rect 13107 568 13118 602
rect 13152 568 13163 602
rect 13107 534 13163 568
rect 13107 500 13118 534
rect 13152 500 13163 534
rect 13107 466 13163 500
rect 13107 432 13118 466
rect 13152 432 13163 466
rect 13107 398 13163 432
rect 13107 364 13118 398
rect 13152 364 13163 398
rect 13107 330 13163 364
rect 13107 296 13118 330
rect 13152 296 13163 330
rect 13107 262 13163 296
rect 13107 228 13118 262
rect 13152 228 13163 262
rect 13107 194 13163 228
rect 13107 160 13118 194
rect 13152 160 13163 194
rect 13107 148 13163 160
rect 13323 1078 13379 1148
rect 13323 1044 13334 1078
rect 13368 1044 13379 1078
rect 13323 1010 13379 1044
rect 13323 976 13334 1010
rect 13368 976 13379 1010
rect 13323 942 13379 976
rect 13323 908 13334 942
rect 13368 908 13379 942
rect 13323 874 13379 908
rect 13323 840 13334 874
rect 13368 840 13379 874
rect 13323 806 13379 840
rect 13323 772 13334 806
rect 13368 772 13379 806
rect 13323 738 13379 772
rect 13323 704 13334 738
rect 13368 704 13379 738
rect 13323 670 13379 704
rect 13323 636 13334 670
rect 13368 636 13379 670
rect 13323 602 13379 636
rect 13323 568 13334 602
rect 13368 568 13379 602
rect 13323 534 13379 568
rect 13323 500 13334 534
rect 13368 500 13379 534
rect 13323 466 13379 500
rect 13323 432 13334 466
rect 13368 432 13379 466
rect 13323 398 13379 432
rect 13323 364 13334 398
rect 13368 364 13379 398
rect 13323 330 13379 364
rect 13323 296 13334 330
rect 13368 296 13379 330
rect 13323 262 13379 296
rect 13323 228 13334 262
rect 13368 228 13379 262
rect 13323 194 13379 228
rect 13323 160 13334 194
rect 13368 160 13379 194
rect 13323 148 13379 160
rect 13539 1078 13595 1148
rect 13539 1044 13550 1078
rect 13584 1044 13595 1078
rect 13539 1010 13595 1044
rect 13539 976 13550 1010
rect 13584 976 13595 1010
rect 13539 942 13595 976
rect 13539 908 13550 942
rect 13584 908 13595 942
rect 13539 874 13595 908
rect 13539 840 13550 874
rect 13584 840 13595 874
rect 13539 806 13595 840
rect 13539 772 13550 806
rect 13584 772 13595 806
rect 13539 738 13595 772
rect 13539 704 13550 738
rect 13584 704 13595 738
rect 13539 670 13595 704
rect 13539 636 13550 670
rect 13584 636 13595 670
rect 13539 602 13595 636
rect 13539 568 13550 602
rect 13584 568 13595 602
rect 13539 534 13595 568
rect 13539 500 13550 534
rect 13584 500 13595 534
rect 13539 466 13595 500
rect 13539 432 13550 466
rect 13584 432 13595 466
rect 13539 398 13595 432
rect 13539 364 13550 398
rect 13584 364 13595 398
rect 13539 330 13595 364
rect 13539 296 13550 330
rect 13584 296 13595 330
rect 13539 262 13595 296
rect 13539 228 13550 262
rect 13584 228 13595 262
rect 13539 194 13595 228
rect 13539 160 13550 194
rect 13584 160 13595 194
rect 13539 148 13595 160
rect 13755 1078 13811 1148
rect 13755 1044 13766 1078
rect 13800 1044 13811 1078
rect 13755 1010 13811 1044
rect 13755 976 13766 1010
rect 13800 976 13811 1010
rect 13755 942 13811 976
rect 13755 908 13766 942
rect 13800 908 13811 942
rect 13755 874 13811 908
rect 13755 840 13766 874
rect 13800 840 13811 874
rect 13755 806 13811 840
rect 13755 772 13766 806
rect 13800 772 13811 806
rect 13755 738 13811 772
rect 13755 704 13766 738
rect 13800 704 13811 738
rect 13755 670 13811 704
rect 13755 636 13766 670
rect 13800 636 13811 670
rect 13755 602 13811 636
rect 13755 568 13766 602
rect 13800 568 13811 602
rect 13755 534 13811 568
rect 13755 500 13766 534
rect 13800 500 13811 534
rect 13755 466 13811 500
rect 13755 432 13766 466
rect 13800 432 13811 466
rect 13755 398 13811 432
rect 13755 364 13766 398
rect 13800 364 13811 398
rect 13755 330 13811 364
rect 13755 296 13766 330
rect 13800 296 13811 330
rect 13755 262 13811 296
rect 13755 228 13766 262
rect 13800 228 13811 262
rect 13755 194 13811 228
rect 13755 160 13766 194
rect 13800 160 13811 194
rect 13755 148 13811 160
rect 13971 1078 14027 1148
rect 13971 1044 13982 1078
rect 14016 1044 14027 1078
rect 13971 1010 14027 1044
rect 13971 976 13982 1010
rect 14016 976 14027 1010
rect 13971 942 14027 976
rect 13971 908 13982 942
rect 14016 908 14027 942
rect 13971 874 14027 908
rect 13971 840 13982 874
rect 14016 840 14027 874
rect 13971 806 14027 840
rect 13971 772 13982 806
rect 14016 772 14027 806
rect 13971 738 14027 772
rect 13971 704 13982 738
rect 14016 704 14027 738
rect 13971 670 14027 704
rect 13971 636 13982 670
rect 14016 636 14027 670
rect 13971 602 14027 636
rect 13971 568 13982 602
rect 14016 568 14027 602
rect 13971 534 14027 568
rect 13971 500 13982 534
rect 14016 500 14027 534
rect 13971 466 14027 500
rect 13971 432 13982 466
rect 14016 432 14027 466
rect 13971 398 14027 432
rect 13971 364 13982 398
rect 14016 364 14027 398
rect 13971 330 14027 364
rect 13971 296 13982 330
rect 14016 296 14027 330
rect 13971 262 14027 296
rect 13971 228 13982 262
rect 14016 228 14027 262
rect 13971 194 14027 228
rect 13971 160 13982 194
rect 14016 160 14027 194
rect 13971 148 14027 160
rect 14187 1078 14243 1148
rect 14187 1044 14198 1078
rect 14232 1044 14243 1078
rect 14187 1010 14243 1044
rect 14187 976 14198 1010
rect 14232 976 14243 1010
rect 14187 942 14243 976
rect 14187 908 14198 942
rect 14232 908 14243 942
rect 14187 874 14243 908
rect 14187 840 14198 874
rect 14232 840 14243 874
rect 14187 806 14243 840
rect 14187 772 14198 806
rect 14232 772 14243 806
rect 14187 738 14243 772
rect 14187 704 14198 738
rect 14232 704 14243 738
rect 14187 670 14243 704
rect 14187 636 14198 670
rect 14232 636 14243 670
rect 14187 602 14243 636
rect 14187 568 14198 602
rect 14232 568 14243 602
rect 14187 534 14243 568
rect 14187 500 14198 534
rect 14232 500 14243 534
rect 14187 466 14243 500
rect 14187 432 14198 466
rect 14232 432 14243 466
rect 14187 398 14243 432
rect 14187 364 14198 398
rect 14232 364 14243 398
rect 14187 330 14243 364
rect 14187 296 14198 330
rect 14232 296 14243 330
rect 14187 262 14243 296
rect 14187 228 14198 262
rect 14232 228 14243 262
rect 14187 194 14243 228
rect 14187 160 14198 194
rect 14232 160 14243 194
rect 14187 148 14243 160
rect 14403 1078 14459 1148
rect 14403 1044 14414 1078
rect 14448 1044 14459 1078
rect 14403 1010 14459 1044
rect 14403 976 14414 1010
rect 14448 976 14459 1010
rect 14403 942 14459 976
rect 14403 908 14414 942
rect 14448 908 14459 942
rect 14403 874 14459 908
rect 14403 840 14414 874
rect 14448 840 14459 874
rect 14403 806 14459 840
rect 14403 772 14414 806
rect 14448 772 14459 806
rect 14403 738 14459 772
rect 14403 704 14414 738
rect 14448 704 14459 738
rect 14403 670 14459 704
rect 14403 636 14414 670
rect 14448 636 14459 670
rect 14403 602 14459 636
rect 14403 568 14414 602
rect 14448 568 14459 602
rect 14403 534 14459 568
rect 14403 500 14414 534
rect 14448 500 14459 534
rect 14403 466 14459 500
rect 14403 432 14414 466
rect 14448 432 14459 466
rect 14403 398 14459 432
rect 14403 364 14414 398
rect 14448 364 14459 398
rect 14403 330 14459 364
rect 14403 296 14414 330
rect 14448 296 14459 330
rect 14403 262 14459 296
rect 14403 228 14414 262
rect 14448 228 14459 262
rect 14403 194 14459 228
rect 14403 160 14414 194
rect 14448 160 14459 194
rect 14403 148 14459 160
rect 14619 1078 14675 1148
rect 14619 1044 14630 1078
rect 14664 1044 14675 1078
rect 14619 1010 14675 1044
rect 14619 976 14630 1010
rect 14664 976 14675 1010
rect 14619 942 14675 976
rect 14619 908 14630 942
rect 14664 908 14675 942
rect 14619 874 14675 908
rect 14619 840 14630 874
rect 14664 840 14675 874
rect 14619 806 14675 840
rect 14619 772 14630 806
rect 14664 772 14675 806
rect 14619 738 14675 772
rect 14619 704 14630 738
rect 14664 704 14675 738
rect 14619 670 14675 704
rect 14619 636 14630 670
rect 14664 636 14675 670
rect 14619 602 14675 636
rect 14619 568 14630 602
rect 14664 568 14675 602
rect 14619 534 14675 568
rect 14619 500 14630 534
rect 14664 500 14675 534
rect 14619 466 14675 500
rect 14619 432 14630 466
rect 14664 432 14675 466
rect 14619 398 14675 432
rect 14619 364 14630 398
rect 14664 364 14675 398
rect 14619 330 14675 364
rect 14619 296 14630 330
rect 14664 296 14675 330
rect 14619 262 14675 296
rect 14619 228 14630 262
rect 14664 228 14675 262
rect 14619 194 14675 228
rect 14619 160 14630 194
rect 14664 160 14675 194
rect 14619 148 14675 160
rect 14835 1078 14891 1148
rect 14835 1044 14846 1078
rect 14880 1044 14891 1078
rect 14835 1010 14891 1044
rect 14835 976 14846 1010
rect 14880 976 14891 1010
rect 14835 942 14891 976
rect 14835 908 14846 942
rect 14880 908 14891 942
rect 14835 874 14891 908
rect 14835 840 14846 874
rect 14880 840 14891 874
rect 14835 806 14891 840
rect 14835 772 14846 806
rect 14880 772 14891 806
rect 14835 738 14891 772
rect 14835 704 14846 738
rect 14880 704 14891 738
rect 14835 670 14891 704
rect 14835 636 14846 670
rect 14880 636 14891 670
rect 14835 602 14891 636
rect 14835 568 14846 602
rect 14880 568 14891 602
rect 14835 534 14891 568
rect 14835 500 14846 534
rect 14880 500 14891 534
rect 14835 466 14891 500
rect 14835 432 14846 466
rect 14880 432 14891 466
rect 14835 398 14891 432
rect 14835 364 14846 398
rect 14880 364 14891 398
rect 14835 330 14891 364
rect 14835 296 14846 330
rect 14880 296 14891 330
rect 14835 262 14891 296
rect 14835 228 14846 262
rect 14880 228 14891 262
rect 14835 194 14891 228
rect 14835 160 14846 194
rect 14880 160 14891 194
rect 14835 148 14891 160
rect 15051 1078 15104 1148
rect 15051 1044 15062 1078
rect 15096 1044 15104 1078
rect 15051 1010 15104 1044
rect 15051 976 15062 1010
rect 15096 976 15104 1010
rect 15051 942 15104 976
rect 15051 908 15062 942
rect 15096 908 15104 942
rect 15051 874 15104 908
rect 15051 840 15062 874
rect 15096 840 15104 874
rect 15051 806 15104 840
rect 15051 772 15062 806
rect 15096 772 15104 806
rect 15051 738 15104 772
rect 15051 704 15062 738
rect 15096 704 15104 738
rect 15051 670 15104 704
rect 15051 636 15062 670
rect 15096 636 15104 670
rect 15051 602 15104 636
rect 15051 568 15062 602
rect 15096 568 15104 602
rect 15051 534 15104 568
rect 15164 1070 15217 1148
rect 15164 1036 15172 1070
rect 15206 1036 15217 1070
rect 15164 1002 15217 1036
rect 15164 968 15172 1002
rect 15206 968 15217 1002
rect 15164 934 15217 968
rect 15164 900 15172 934
rect 15206 900 15217 934
rect 15164 866 15217 900
rect 15164 832 15172 866
rect 15206 832 15217 866
rect 15164 798 15217 832
rect 15164 764 15172 798
rect 15206 764 15217 798
rect 15164 730 15217 764
rect 15164 696 15172 730
rect 15206 696 15217 730
rect 15164 662 15217 696
rect 15164 628 15172 662
rect 15206 628 15217 662
rect 15164 594 15217 628
rect 15164 560 15172 594
rect 15206 560 15217 594
rect 15164 548 15217 560
rect 15417 1070 15470 1148
rect 15417 1036 15428 1070
rect 15462 1036 15470 1070
rect 15417 1002 15470 1036
rect 15417 968 15428 1002
rect 15462 968 15470 1002
rect 15417 934 15470 968
rect 15417 900 15428 934
rect 15462 900 15470 934
rect 15417 866 15470 900
rect 15417 832 15428 866
rect 15462 832 15470 866
rect 15417 798 15470 832
rect 15417 764 15428 798
rect 15462 764 15470 798
rect 15417 730 15470 764
rect 15417 696 15428 730
rect 15462 696 15470 730
rect 15417 662 15470 696
rect 15417 628 15428 662
rect 15462 628 15470 662
rect 15417 594 15470 628
rect 15417 560 15428 594
rect 15462 560 15470 594
rect 15417 548 15470 560
rect 15530 1078 15583 1148
rect 15530 1044 15538 1078
rect 15572 1044 15583 1078
rect 15530 1010 15583 1044
rect 15530 976 15538 1010
rect 15572 976 15583 1010
rect 15530 942 15583 976
rect 15530 908 15538 942
rect 15572 908 15583 942
rect 15530 874 15583 908
rect 15530 840 15538 874
rect 15572 840 15583 874
rect 15530 806 15583 840
rect 15530 772 15538 806
rect 15572 772 15583 806
rect 15530 738 15583 772
rect 15530 704 15538 738
rect 15572 704 15583 738
rect 15530 670 15583 704
rect 15530 636 15538 670
rect 15572 636 15583 670
rect 15530 602 15583 636
rect 15530 568 15538 602
rect 15572 568 15583 602
rect 15051 500 15062 534
rect 15096 500 15104 534
rect 15530 534 15583 568
rect 15051 466 15104 500
rect 15051 432 15062 466
rect 15096 432 15104 466
rect 15051 398 15104 432
rect 15051 364 15062 398
rect 15096 364 15104 398
rect 15051 330 15104 364
rect 15051 296 15062 330
rect 15096 296 15104 330
rect 15051 262 15104 296
rect 15051 228 15062 262
rect 15096 228 15104 262
rect 15051 194 15104 228
rect 15051 160 15062 194
rect 15096 160 15104 194
rect 15051 148 15104 160
rect 15530 500 15538 534
rect 15572 500 15583 534
rect 15530 466 15583 500
rect 15530 432 15538 466
rect 15572 432 15583 466
rect 15530 398 15583 432
rect 15530 364 15538 398
rect 15572 364 15583 398
rect 15530 330 15583 364
rect 15530 296 15538 330
rect 15572 296 15583 330
rect 15530 262 15583 296
rect 15530 228 15538 262
rect 15572 228 15583 262
rect 15530 194 15583 228
rect 15530 160 15538 194
rect 15572 160 15583 194
rect 15530 148 15583 160
rect 15743 1078 15799 1148
rect 15743 1044 15754 1078
rect 15788 1044 15799 1078
rect 15743 1010 15799 1044
rect 15743 976 15754 1010
rect 15788 976 15799 1010
rect 15743 942 15799 976
rect 15743 908 15754 942
rect 15788 908 15799 942
rect 15743 874 15799 908
rect 15743 840 15754 874
rect 15788 840 15799 874
rect 15743 806 15799 840
rect 15743 772 15754 806
rect 15788 772 15799 806
rect 15743 738 15799 772
rect 15743 704 15754 738
rect 15788 704 15799 738
rect 15743 670 15799 704
rect 15743 636 15754 670
rect 15788 636 15799 670
rect 15743 602 15799 636
rect 15743 568 15754 602
rect 15788 568 15799 602
rect 15743 534 15799 568
rect 15743 500 15754 534
rect 15788 500 15799 534
rect 15743 466 15799 500
rect 15743 432 15754 466
rect 15788 432 15799 466
rect 15743 398 15799 432
rect 15743 364 15754 398
rect 15788 364 15799 398
rect 15743 330 15799 364
rect 15743 296 15754 330
rect 15788 296 15799 330
rect 15743 262 15799 296
rect 15743 228 15754 262
rect 15788 228 15799 262
rect 15743 194 15799 228
rect 15743 160 15754 194
rect 15788 160 15799 194
rect 15743 148 15799 160
rect 15959 1078 16012 1148
rect 15959 1044 15970 1078
rect 16004 1044 16012 1078
rect 15959 1010 16012 1044
rect 15959 976 15970 1010
rect 16004 976 16012 1010
rect 15959 942 16012 976
rect 15959 908 15970 942
rect 16004 908 16012 942
rect 15959 874 16012 908
rect 15959 840 15970 874
rect 16004 840 16012 874
rect 15959 806 16012 840
rect 15959 772 15970 806
rect 16004 772 16012 806
rect 15959 738 16012 772
rect 15959 704 15970 738
rect 16004 704 16012 738
rect 15959 670 16012 704
rect 15959 636 15970 670
rect 16004 636 16012 670
rect 15959 602 16012 636
rect 15959 568 15970 602
rect 16004 568 16012 602
rect 15959 534 16012 568
rect 15959 500 15970 534
rect 16004 500 16012 534
rect 15959 466 16012 500
rect 15959 432 15970 466
rect 16004 432 16012 466
rect 15959 398 16012 432
rect 15959 364 15970 398
rect 16004 364 16012 398
rect 15959 330 16012 364
rect 15959 296 15970 330
rect 16004 296 16012 330
rect 15959 262 16012 296
rect 15959 228 15970 262
rect 16004 228 16012 262
rect 15959 194 16012 228
rect 15959 160 15970 194
rect 16004 160 16012 194
rect 15959 148 16012 160
<< mvpdiff >>
rect 712 2851 765 2921
rect 712 2817 720 2851
rect 754 2817 765 2851
rect 712 2783 765 2817
rect 712 2749 720 2783
rect 754 2749 765 2783
rect 712 2715 765 2749
rect 712 2681 720 2715
rect 754 2681 765 2715
rect 712 2647 765 2681
rect 712 2613 720 2647
rect 754 2613 765 2647
rect 712 2579 765 2613
rect 712 2545 720 2579
rect 754 2545 765 2579
rect 712 2511 765 2545
rect 712 2477 720 2511
rect 754 2477 765 2511
rect 712 2443 765 2477
rect 712 2409 720 2443
rect 754 2409 765 2443
rect 712 2375 765 2409
rect 712 2341 720 2375
rect 754 2341 765 2375
rect 712 2307 765 2341
rect 712 2273 720 2307
rect 754 2273 765 2307
rect 712 2239 765 2273
rect 712 2205 720 2239
rect 754 2205 765 2239
rect 712 2171 765 2205
rect 712 2137 720 2171
rect 754 2137 765 2171
rect 712 2103 765 2137
rect 712 2069 720 2103
rect 754 2069 765 2103
rect 712 2035 765 2069
rect 712 2001 720 2035
rect 754 2001 765 2035
rect 712 1967 765 2001
rect 712 1933 720 1967
rect 754 1933 765 1967
rect 712 1921 765 1933
rect 865 2851 921 2921
rect 865 2817 876 2851
rect 910 2817 921 2851
rect 865 2783 921 2817
rect 865 2749 876 2783
rect 910 2749 921 2783
rect 865 2715 921 2749
rect 865 2681 876 2715
rect 910 2681 921 2715
rect 865 2647 921 2681
rect 865 2613 876 2647
rect 910 2613 921 2647
rect 865 2579 921 2613
rect 865 2545 876 2579
rect 910 2545 921 2579
rect 865 2511 921 2545
rect 865 2477 876 2511
rect 910 2477 921 2511
rect 865 2443 921 2477
rect 865 2409 876 2443
rect 910 2409 921 2443
rect 865 2375 921 2409
rect 865 2341 876 2375
rect 910 2341 921 2375
rect 865 2307 921 2341
rect 865 2273 876 2307
rect 910 2273 921 2307
rect 865 2239 921 2273
rect 865 2205 876 2239
rect 910 2205 921 2239
rect 865 2171 921 2205
rect 865 2137 876 2171
rect 910 2137 921 2171
rect 865 2103 921 2137
rect 865 2069 876 2103
rect 910 2069 921 2103
rect 865 2035 921 2069
rect 865 2001 876 2035
rect 910 2001 921 2035
rect 865 1967 921 2001
rect 865 1933 876 1967
rect 910 1933 921 1967
rect 865 1921 921 1933
rect 1021 2851 1074 2921
rect 1021 2817 1032 2851
rect 1066 2817 1074 2851
rect 1021 2783 1074 2817
rect 1021 2749 1032 2783
rect 1066 2749 1074 2783
rect 1021 2715 1074 2749
rect 1021 2681 1032 2715
rect 1066 2681 1074 2715
rect 1021 2647 1074 2681
rect 1021 2613 1032 2647
rect 1066 2613 1074 2647
rect 1021 2579 1074 2613
rect 1021 2545 1032 2579
rect 1066 2545 1074 2579
rect 1021 2511 1074 2545
rect 1021 2477 1032 2511
rect 1066 2477 1074 2511
rect 1021 2443 1074 2477
rect 1021 2409 1032 2443
rect 1066 2409 1074 2443
rect 1021 2375 1074 2409
rect 1021 2341 1032 2375
rect 1066 2341 1074 2375
rect 1021 2307 1074 2341
rect 1021 2273 1032 2307
rect 1066 2273 1074 2307
rect 1021 2239 1074 2273
rect 1021 2205 1032 2239
rect 1066 2205 1074 2239
rect 1021 2171 1074 2205
rect 1021 2137 1032 2171
rect 1066 2137 1074 2171
rect 1021 2103 1074 2137
rect 1021 2069 1032 2103
rect 1066 2069 1074 2103
rect 1021 2035 1074 2069
rect 1021 2001 1032 2035
rect 1066 2001 1074 2035
rect 1021 1967 1074 2001
rect 1021 1933 1032 1967
rect 1066 1933 1074 1967
rect 1021 1921 1074 1933
rect 1134 2851 1187 2921
rect 1134 2817 1142 2851
rect 1176 2817 1187 2851
rect 1134 2783 1187 2817
rect 1134 2749 1142 2783
rect 1176 2749 1187 2783
rect 1134 2715 1187 2749
rect 1134 2681 1142 2715
rect 1176 2681 1187 2715
rect 1134 2647 1187 2681
rect 1134 2613 1142 2647
rect 1176 2613 1187 2647
rect 1134 2579 1187 2613
rect 1134 2545 1142 2579
rect 1176 2545 1187 2579
rect 1134 2511 1187 2545
rect 1134 2477 1142 2511
rect 1176 2477 1187 2511
rect 1134 2443 1187 2477
rect 1134 2409 1142 2443
rect 1176 2409 1187 2443
rect 1134 2375 1187 2409
rect 1134 2341 1142 2375
rect 1176 2341 1187 2375
rect 1134 2307 1187 2341
rect 1134 2273 1142 2307
rect 1176 2273 1187 2307
rect 1134 2239 1187 2273
rect 1134 2205 1142 2239
rect 1176 2205 1187 2239
rect 1134 2171 1187 2205
rect 1134 2137 1142 2171
rect 1176 2137 1187 2171
rect 1134 2103 1187 2137
rect 1134 2069 1142 2103
rect 1176 2069 1187 2103
rect 1134 2035 1187 2069
rect 1134 2001 1142 2035
rect 1176 2001 1187 2035
rect 1134 1967 1187 2001
rect 1134 1933 1142 1967
rect 1176 1933 1187 1967
rect 1134 1921 1187 1933
rect 1287 2851 1343 2921
rect 1287 2817 1298 2851
rect 1332 2817 1343 2851
rect 1287 2783 1343 2817
rect 1287 2749 1298 2783
rect 1332 2749 1343 2783
rect 1287 2715 1343 2749
rect 1287 2681 1298 2715
rect 1332 2681 1343 2715
rect 1287 2647 1343 2681
rect 1287 2613 1298 2647
rect 1332 2613 1343 2647
rect 1287 2579 1343 2613
rect 1287 2545 1298 2579
rect 1332 2545 1343 2579
rect 1287 2511 1343 2545
rect 1287 2477 1298 2511
rect 1332 2477 1343 2511
rect 1287 2443 1343 2477
rect 1287 2409 1298 2443
rect 1332 2409 1343 2443
rect 1287 2375 1343 2409
rect 1287 2341 1298 2375
rect 1332 2341 1343 2375
rect 1287 2307 1343 2341
rect 1287 2273 1298 2307
rect 1332 2273 1343 2307
rect 1287 2239 1343 2273
rect 1287 2205 1298 2239
rect 1332 2205 1343 2239
rect 1287 2171 1343 2205
rect 1287 2137 1298 2171
rect 1332 2137 1343 2171
rect 1287 2103 1343 2137
rect 1287 2069 1298 2103
rect 1332 2069 1343 2103
rect 1287 2035 1343 2069
rect 1287 2001 1298 2035
rect 1332 2001 1343 2035
rect 1287 1967 1343 2001
rect 1287 1933 1298 1967
rect 1332 1933 1343 1967
rect 1287 1921 1343 1933
rect 1443 2851 1499 2921
rect 1443 2817 1454 2851
rect 1488 2817 1499 2851
rect 1443 2783 1499 2817
rect 1443 2749 1454 2783
rect 1488 2749 1499 2783
rect 1443 2715 1499 2749
rect 1443 2681 1454 2715
rect 1488 2681 1499 2715
rect 1443 2647 1499 2681
rect 1443 2613 1454 2647
rect 1488 2613 1499 2647
rect 1443 2579 1499 2613
rect 1443 2545 1454 2579
rect 1488 2545 1499 2579
rect 1443 2511 1499 2545
rect 1443 2477 1454 2511
rect 1488 2477 1499 2511
rect 1443 2443 1499 2477
rect 1443 2409 1454 2443
rect 1488 2409 1499 2443
rect 1443 2375 1499 2409
rect 1443 2341 1454 2375
rect 1488 2341 1499 2375
rect 1443 2307 1499 2341
rect 1443 2273 1454 2307
rect 1488 2273 1499 2307
rect 1443 2239 1499 2273
rect 1443 2205 1454 2239
rect 1488 2205 1499 2239
rect 1443 2171 1499 2205
rect 1443 2137 1454 2171
rect 1488 2137 1499 2171
rect 1443 2103 1499 2137
rect 1443 2069 1454 2103
rect 1488 2069 1499 2103
rect 1443 2035 1499 2069
rect 1443 2001 1454 2035
rect 1488 2001 1499 2035
rect 1443 1967 1499 2001
rect 1443 1933 1454 1967
rect 1488 1933 1499 1967
rect 1443 1921 1499 1933
rect 1599 2851 1655 2921
rect 1599 2817 1610 2851
rect 1644 2817 1655 2851
rect 1599 2783 1655 2817
rect 1599 2749 1610 2783
rect 1644 2749 1655 2783
rect 1599 2715 1655 2749
rect 1599 2681 1610 2715
rect 1644 2681 1655 2715
rect 1599 2647 1655 2681
rect 1599 2613 1610 2647
rect 1644 2613 1655 2647
rect 1599 2579 1655 2613
rect 1599 2545 1610 2579
rect 1644 2545 1655 2579
rect 1599 2511 1655 2545
rect 1599 2477 1610 2511
rect 1644 2477 1655 2511
rect 1599 2443 1655 2477
rect 1599 2409 1610 2443
rect 1644 2409 1655 2443
rect 1599 2375 1655 2409
rect 1599 2341 1610 2375
rect 1644 2341 1655 2375
rect 1599 2307 1655 2341
rect 1599 2273 1610 2307
rect 1644 2273 1655 2307
rect 1599 2239 1655 2273
rect 1599 2205 1610 2239
rect 1644 2205 1655 2239
rect 1599 2171 1655 2205
rect 1599 2137 1610 2171
rect 1644 2137 1655 2171
rect 1599 2103 1655 2137
rect 1599 2069 1610 2103
rect 1644 2069 1655 2103
rect 1599 2035 1655 2069
rect 1599 2001 1610 2035
rect 1644 2001 1655 2035
rect 1599 1967 1655 2001
rect 1599 1933 1610 1967
rect 1644 1933 1655 1967
rect 1599 1921 1655 1933
rect 1755 2851 1811 2921
rect 1755 2817 1766 2851
rect 1800 2817 1811 2851
rect 1755 2783 1811 2817
rect 1755 2749 1766 2783
rect 1800 2749 1811 2783
rect 1755 2715 1811 2749
rect 1755 2681 1766 2715
rect 1800 2681 1811 2715
rect 1755 2647 1811 2681
rect 1755 2613 1766 2647
rect 1800 2613 1811 2647
rect 1755 2579 1811 2613
rect 1755 2545 1766 2579
rect 1800 2545 1811 2579
rect 1755 2511 1811 2545
rect 1755 2477 1766 2511
rect 1800 2477 1811 2511
rect 1755 2443 1811 2477
rect 1755 2409 1766 2443
rect 1800 2409 1811 2443
rect 1755 2375 1811 2409
rect 1755 2341 1766 2375
rect 1800 2341 1811 2375
rect 1755 2307 1811 2341
rect 1755 2273 1766 2307
rect 1800 2273 1811 2307
rect 1755 2239 1811 2273
rect 1755 2205 1766 2239
rect 1800 2205 1811 2239
rect 1755 2171 1811 2205
rect 1755 2137 1766 2171
rect 1800 2137 1811 2171
rect 1755 2103 1811 2137
rect 1755 2069 1766 2103
rect 1800 2069 1811 2103
rect 1755 2035 1811 2069
rect 1755 2001 1766 2035
rect 1800 2001 1811 2035
rect 1755 1967 1811 2001
rect 1755 1933 1766 1967
rect 1800 1933 1811 1967
rect 1755 1921 1811 1933
rect 1911 2851 1967 2921
rect 1911 2817 1922 2851
rect 1956 2817 1967 2851
rect 1911 2783 1967 2817
rect 1911 2749 1922 2783
rect 1956 2749 1967 2783
rect 1911 2715 1967 2749
rect 1911 2681 1922 2715
rect 1956 2681 1967 2715
rect 1911 2647 1967 2681
rect 1911 2613 1922 2647
rect 1956 2613 1967 2647
rect 1911 2579 1967 2613
rect 1911 2545 1922 2579
rect 1956 2545 1967 2579
rect 1911 2511 1967 2545
rect 1911 2477 1922 2511
rect 1956 2477 1967 2511
rect 1911 2443 1967 2477
rect 1911 2409 1922 2443
rect 1956 2409 1967 2443
rect 1911 2375 1967 2409
rect 1911 2341 1922 2375
rect 1956 2341 1967 2375
rect 1911 2307 1967 2341
rect 1911 2273 1922 2307
rect 1956 2273 1967 2307
rect 1911 2239 1967 2273
rect 1911 2205 1922 2239
rect 1956 2205 1967 2239
rect 1911 2171 1967 2205
rect 1911 2137 1922 2171
rect 1956 2137 1967 2171
rect 1911 2103 1967 2137
rect 1911 2069 1922 2103
rect 1956 2069 1967 2103
rect 1911 2035 1967 2069
rect 1911 2001 1922 2035
rect 1956 2001 1967 2035
rect 1911 1967 1967 2001
rect 1911 1933 1922 1967
rect 1956 1933 1967 1967
rect 1911 1921 1967 1933
rect 2067 2851 2123 2921
rect 2067 2817 2078 2851
rect 2112 2817 2123 2851
rect 2067 2783 2123 2817
rect 2067 2749 2078 2783
rect 2112 2749 2123 2783
rect 2067 2715 2123 2749
rect 2067 2681 2078 2715
rect 2112 2681 2123 2715
rect 2067 2647 2123 2681
rect 2067 2613 2078 2647
rect 2112 2613 2123 2647
rect 2067 2579 2123 2613
rect 2067 2545 2078 2579
rect 2112 2545 2123 2579
rect 2067 2511 2123 2545
rect 2067 2477 2078 2511
rect 2112 2477 2123 2511
rect 2067 2443 2123 2477
rect 2067 2409 2078 2443
rect 2112 2409 2123 2443
rect 2067 2375 2123 2409
rect 2067 2341 2078 2375
rect 2112 2341 2123 2375
rect 2067 2307 2123 2341
rect 2067 2273 2078 2307
rect 2112 2273 2123 2307
rect 2067 2239 2123 2273
rect 2067 2205 2078 2239
rect 2112 2205 2123 2239
rect 2067 2171 2123 2205
rect 2067 2137 2078 2171
rect 2112 2137 2123 2171
rect 2067 2103 2123 2137
rect 2067 2069 2078 2103
rect 2112 2069 2123 2103
rect 2067 2035 2123 2069
rect 2067 2001 2078 2035
rect 2112 2001 2123 2035
rect 2067 1967 2123 2001
rect 2067 1933 2078 1967
rect 2112 1933 2123 1967
rect 2067 1921 2123 1933
rect 2223 2851 2279 2921
rect 2223 2817 2234 2851
rect 2268 2817 2279 2851
rect 2223 2783 2279 2817
rect 2223 2749 2234 2783
rect 2268 2749 2279 2783
rect 2223 2715 2279 2749
rect 2223 2681 2234 2715
rect 2268 2681 2279 2715
rect 2223 2647 2279 2681
rect 2223 2613 2234 2647
rect 2268 2613 2279 2647
rect 2223 2579 2279 2613
rect 2223 2545 2234 2579
rect 2268 2545 2279 2579
rect 2223 2511 2279 2545
rect 2223 2477 2234 2511
rect 2268 2477 2279 2511
rect 2223 2443 2279 2477
rect 2223 2409 2234 2443
rect 2268 2409 2279 2443
rect 2223 2375 2279 2409
rect 2223 2341 2234 2375
rect 2268 2341 2279 2375
rect 2223 2307 2279 2341
rect 2223 2273 2234 2307
rect 2268 2273 2279 2307
rect 2223 2239 2279 2273
rect 2223 2205 2234 2239
rect 2268 2205 2279 2239
rect 2223 2171 2279 2205
rect 2223 2137 2234 2171
rect 2268 2137 2279 2171
rect 2223 2103 2279 2137
rect 2223 2069 2234 2103
rect 2268 2069 2279 2103
rect 2223 2035 2279 2069
rect 2223 2001 2234 2035
rect 2268 2001 2279 2035
rect 2223 1967 2279 2001
rect 2223 1933 2234 1967
rect 2268 1933 2279 1967
rect 2223 1921 2279 1933
rect 2379 2851 2435 2921
rect 2379 2817 2390 2851
rect 2424 2817 2435 2851
rect 2379 2783 2435 2817
rect 2379 2749 2390 2783
rect 2424 2749 2435 2783
rect 2379 2715 2435 2749
rect 2379 2681 2390 2715
rect 2424 2681 2435 2715
rect 2379 2647 2435 2681
rect 2379 2613 2390 2647
rect 2424 2613 2435 2647
rect 2379 2579 2435 2613
rect 2379 2545 2390 2579
rect 2424 2545 2435 2579
rect 2379 2511 2435 2545
rect 2379 2477 2390 2511
rect 2424 2477 2435 2511
rect 2379 2443 2435 2477
rect 2379 2409 2390 2443
rect 2424 2409 2435 2443
rect 2379 2375 2435 2409
rect 2379 2341 2390 2375
rect 2424 2341 2435 2375
rect 2379 2307 2435 2341
rect 2379 2273 2390 2307
rect 2424 2273 2435 2307
rect 2379 2239 2435 2273
rect 2379 2205 2390 2239
rect 2424 2205 2435 2239
rect 2379 2171 2435 2205
rect 2379 2137 2390 2171
rect 2424 2137 2435 2171
rect 2379 2103 2435 2137
rect 2379 2069 2390 2103
rect 2424 2069 2435 2103
rect 2379 2035 2435 2069
rect 2379 2001 2390 2035
rect 2424 2001 2435 2035
rect 2379 1967 2435 2001
rect 2379 1933 2390 1967
rect 2424 1933 2435 1967
rect 2379 1921 2435 1933
rect 2535 2851 2591 2921
rect 2535 2817 2546 2851
rect 2580 2817 2591 2851
rect 2535 2783 2591 2817
rect 2535 2749 2546 2783
rect 2580 2749 2591 2783
rect 2535 2715 2591 2749
rect 2535 2681 2546 2715
rect 2580 2681 2591 2715
rect 2535 2647 2591 2681
rect 2535 2613 2546 2647
rect 2580 2613 2591 2647
rect 2535 2579 2591 2613
rect 2535 2545 2546 2579
rect 2580 2545 2591 2579
rect 2535 2511 2591 2545
rect 2535 2477 2546 2511
rect 2580 2477 2591 2511
rect 2535 2443 2591 2477
rect 2535 2409 2546 2443
rect 2580 2409 2591 2443
rect 2535 2375 2591 2409
rect 2535 2341 2546 2375
rect 2580 2341 2591 2375
rect 2535 2307 2591 2341
rect 2535 2273 2546 2307
rect 2580 2273 2591 2307
rect 2535 2239 2591 2273
rect 2535 2205 2546 2239
rect 2580 2205 2591 2239
rect 2535 2171 2591 2205
rect 2535 2137 2546 2171
rect 2580 2137 2591 2171
rect 2535 2103 2591 2137
rect 2535 2069 2546 2103
rect 2580 2069 2591 2103
rect 2535 2035 2591 2069
rect 2535 2001 2546 2035
rect 2580 2001 2591 2035
rect 2535 1967 2591 2001
rect 2535 1933 2546 1967
rect 2580 1933 2591 1967
rect 2535 1921 2591 1933
rect 2691 2851 2747 2921
rect 2691 2817 2702 2851
rect 2736 2817 2747 2851
rect 2691 2783 2747 2817
rect 2691 2749 2702 2783
rect 2736 2749 2747 2783
rect 2691 2715 2747 2749
rect 2691 2681 2702 2715
rect 2736 2681 2747 2715
rect 2691 2647 2747 2681
rect 2691 2613 2702 2647
rect 2736 2613 2747 2647
rect 2691 2579 2747 2613
rect 2691 2545 2702 2579
rect 2736 2545 2747 2579
rect 2691 2511 2747 2545
rect 2691 2477 2702 2511
rect 2736 2477 2747 2511
rect 2691 2443 2747 2477
rect 2691 2409 2702 2443
rect 2736 2409 2747 2443
rect 2691 2375 2747 2409
rect 2691 2341 2702 2375
rect 2736 2341 2747 2375
rect 2691 2307 2747 2341
rect 2691 2273 2702 2307
rect 2736 2273 2747 2307
rect 2691 2239 2747 2273
rect 2691 2205 2702 2239
rect 2736 2205 2747 2239
rect 2691 2171 2747 2205
rect 2691 2137 2702 2171
rect 2736 2137 2747 2171
rect 2691 2103 2747 2137
rect 2691 2069 2702 2103
rect 2736 2069 2747 2103
rect 2691 2035 2747 2069
rect 2691 2001 2702 2035
rect 2736 2001 2747 2035
rect 2691 1967 2747 2001
rect 2691 1933 2702 1967
rect 2736 1933 2747 1967
rect 2691 1921 2747 1933
rect 2847 2851 2903 2921
rect 2847 2817 2858 2851
rect 2892 2817 2903 2851
rect 2847 2783 2903 2817
rect 2847 2749 2858 2783
rect 2892 2749 2903 2783
rect 2847 2715 2903 2749
rect 2847 2681 2858 2715
rect 2892 2681 2903 2715
rect 2847 2647 2903 2681
rect 2847 2613 2858 2647
rect 2892 2613 2903 2647
rect 2847 2579 2903 2613
rect 2847 2545 2858 2579
rect 2892 2545 2903 2579
rect 2847 2511 2903 2545
rect 2847 2477 2858 2511
rect 2892 2477 2903 2511
rect 2847 2443 2903 2477
rect 2847 2409 2858 2443
rect 2892 2409 2903 2443
rect 2847 2375 2903 2409
rect 2847 2341 2858 2375
rect 2892 2341 2903 2375
rect 2847 2307 2903 2341
rect 2847 2273 2858 2307
rect 2892 2273 2903 2307
rect 2847 2239 2903 2273
rect 2847 2205 2858 2239
rect 2892 2205 2903 2239
rect 2847 2171 2903 2205
rect 2847 2137 2858 2171
rect 2892 2137 2903 2171
rect 2847 2103 2903 2137
rect 2847 2069 2858 2103
rect 2892 2069 2903 2103
rect 2847 2035 2903 2069
rect 2847 2001 2858 2035
rect 2892 2001 2903 2035
rect 2847 1967 2903 2001
rect 2847 1933 2858 1967
rect 2892 1933 2903 1967
rect 2847 1921 2903 1933
rect 3003 2851 3059 2921
rect 3003 2817 3014 2851
rect 3048 2817 3059 2851
rect 3003 2783 3059 2817
rect 3003 2749 3014 2783
rect 3048 2749 3059 2783
rect 3003 2715 3059 2749
rect 3003 2681 3014 2715
rect 3048 2681 3059 2715
rect 3003 2647 3059 2681
rect 3003 2613 3014 2647
rect 3048 2613 3059 2647
rect 3003 2579 3059 2613
rect 3003 2545 3014 2579
rect 3048 2545 3059 2579
rect 3003 2511 3059 2545
rect 3003 2477 3014 2511
rect 3048 2477 3059 2511
rect 3003 2443 3059 2477
rect 3003 2409 3014 2443
rect 3048 2409 3059 2443
rect 3003 2375 3059 2409
rect 3003 2341 3014 2375
rect 3048 2341 3059 2375
rect 3003 2307 3059 2341
rect 3003 2273 3014 2307
rect 3048 2273 3059 2307
rect 3003 2239 3059 2273
rect 3003 2205 3014 2239
rect 3048 2205 3059 2239
rect 3003 2171 3059 2205
rect 3003 2137 3014 2171
rect 3048 2137 3059 2171
rect 3003 2103 3059 2137
rect 3003 2069 3014 2103
rect 3048 2069 3059 2103
rect 3003 2035 3059 2069
rect 3003 2001 3014 2035
rect 3048 2001 3059 2035
rect 3003 1967 3059 2001
rect 3003 1933 3014 1967
rect 3048 1933 3059 1967
rect 3003 1921 3059 1933
rect 3159 2851 3215 2921
rect 3159 2817 3170 2851
rect 3204 2817 3215 2851
rect 3159 2783 3215 2817
rect 3159 2749 3170 2783
rect 3204 2749 3215 2783
rect 3159 2715 3215 2749
rect 3159 2681 3170 2715
rect 3204 2681 3215 2715
rect 3159 2647 3215 2681
rect 3159 2613 3170 2647
rect 3204 2613 3215 2647
rect 3159 2579 3215 2613
rect 3159 2545 3170 2579
rect 3204 2545 3215 2579
rect 3159 2511 3215 2545
rect 3159 2477 3170 2511
rect 3204 2477 3215 2511
rect 3159 2443 3215 2477
rect 3159 2409 3170 2443
rect 3204 2409 3215 2443
rect 3159 2375 3215 2409
rect 3159 2341 3170 2375
rect 3204 2341 3215 2375
rect 3159 2307 3215 2341
rect 3159 2273 3170 2307
rect 3204 2273 3215 2307
rect 3159 2239 3215 2273
rect 3159 2205 3170 2239
rect 3204 2205 3215 2239
rect 3159 2171 3215 2205
rect 3159 2137 3170 2171
rect 3204 2137 3215 2171
rect 3159 2103 3215 2137
rect 3159 2069 3170 2103
rect 3204 2069 3215 2103
rect 3159 2035 3215 2069
rect 3159 2001 3170 2035
rect 3204 2001 3215 2035
rect 3159 1967 3215 2001
rect 3159 1933 3170 1967
rect 3204 1933 3215 1967
rect 3159 1921 3215 1933
rect 3315 2851 3371 2921
rect 3315 2817 3326 2851
rect 3360 2817 3371 2851
rect 3315 2783 3371 2817
rect 3315 2749 3326 2783
rect 3360 2749 3371 2783
rect 3315 2715 3371 2749
rect 3315 2681 3326 2715
rect 3360 2681 3371 2715
rect 3315 2647 3371 2681
rect 3315 2613 3326 2647
rect 3360 2613 3371 2647
rect 3315 2579 3371 2613
rect 3315 2545 3326 2579
rect 3360 2545 3371 2579
rect 3315 2511 3371 2545
rect 3315 2477 3326 2511
rect 3360 2477 3371 2511
rect 3315 2443 3371 2477
rect 3315 2409 3326 2443
rect 3360 2409 3371 2443
rect 3315 2375 3371 2409
rect 3315 2341 3326 2375
rect 3360 2341 3371 2375
rect 3315 2307 3371 2341
rect 3315 2273 3326 2307
rect 3360 2273 3371 2307
rect 3315 2239 3371 2273
rect 3315 2205 3326 2239
rect 3360 2205 3371 2239
rect 3315 2171 3371 2205
rect 3315 2137 3326 2171
rect 3360 2137 3371 2171
rect 3315 2103 3371 2137
rect 3315 2069 3326 2103
rect 3360 2069 3371 2103
rect 3315 2035 3371 2069
rect 3315 2001 3326 2035
rect 3360 2001 3371 2035
rect 3315 1967 3371 2001
rect 3315 1933 3326 1967
rect 3360 1933 3371 1967
rect 3315 1921 3371 1933
rect 3471 2851 3527 2921
rect 3471 2817 3482 2851
rect 3516 2817 3527 2851
rect 3471 2783 3527 2817
rect 3471 2749 3482 2783
rect 3516 2749 3527 2783
rect 3471 2715 3527 2749
rect 3471 2681 3482 2715
rect 3516 2681 3527 2715
rect 3471 2647 3527 2681
rect 3471 2613 3482 2647
rect 3516 2613 3527 2647
rect 3471 2579 3527 2613
rect 3471 2545 3482 2579
rect 3516 2545 3527 2579
rect 3471 2511 3527 2545
rect 3471 2477 3482 2511
rect 3516 2477 3527 2511
rect 3471 2443 3527 2477
rect 3471 2409 3482 2443
rect 3516 2409 3527 2443
rect 3471 2375 3527 2409
rect 3471 2341 3482 2375
rect 3516 2341 3527 2375
rect 3471 2307 3527 2341
rect 3471 2273 3482 2307
rect 3516 2273 3527 2307
rect 3471 2239 3527 2273
rect 3471 2205 3482 2239
rect 3516 2205 3527 2239
rect 3471 2171 3527 2205
rect 3471 2137 3482 2171
rect 3516 2137 3527 2171
rect 3471 2103 3527 2137
rect 3471 2069 3482 2103
rect 3516 2069 3527 2103
rect 3471 2035 3527 2069
rect 3471 2001 3482 2035
rect 3516 2001 3527 2035
rect 3471 1967 3527 2001
rect 3471 1933 3482 1967
rect 3516 1933 3527 1967
rect 3471 1921 3527 1933
rect 3627 2851 3683 2921
rect 3627 2817 3638 2851
rect 3672 2817 3683 2851
rect 3627 2783 3683 2817
rect 3627 2749 3638 2783
rect 3672 2749 3683 2783
rect 3627 2715 3683 2749
rect 3627 2681 3638 2715
rect 3672 2681 3683 2715
rect 3627 2647 3683 2681
rect 3627 2613 3638 2647
rect 3672 2613 3683 2647
rect 3627 2579 3683 2613
rect 3627 2545 3638 2579
rect 3672 2545 3683 2579
rect 3627 2511 3683 2545
rect 3627 2477 3638 2511
rect 3672 2477 3683 2511
rect 3627 2443 3683 2477
rect 3627 2409 3638 2443
rect 3672 2409 3683 2443
rect 3627 2375 3683 2409
rect 3627 2341 3638 2375
rect 3672 2341 3683 2375
rect 3627 2307 3683 2341
rect 3627 2273 3638 2307
rect 3672 2273 3683 2307
rect 3627 2239 3683 2273
rect 3627 2205 3638 2239
rect 3672 2205 3683 2239
rect 3627 2171 3683 2205
rect 3627 2137 3638 2171
rect 3672 2137 3683 2171
rect 3627 2103 3683 2137
rect 3627 2069 3638 2103
rect 3672 2069 3683 2103
rect 3627 2035 3683 2069
rect 3627 2001 3638 2035
rect 3672 2001 3683 2035
rect 3627 1967 3683 2001
rect 3627 1933 3638 1967
rect 3672 1933 3683 1967
rect 3627 1921 3683 1933
rect 3783 2851 3839 2921
rect 3783 2817 3794 2851
rect 3828 2817 3839 2851
rect 3783 2783 3839 2817
rect 3783 2749 3794 2783
rect 3828 2749 3839 2783
rect 3783 2715 3839 2749
rect 3783 2681 3794 2715
rect 3828 2681 3839 2715
rect 3783 2647 3839 2681
rect 3783 2613 3794 2647
rect 3828 2613 3839 2647
rect 3783 2579 3839 2613
rect 3783 2545 3794 2579
rect 3828 2545 3839 2579
rect 3783 2511 3839 2545
rect 3783 2477 3794 2511
rect 3828 2477 3839 2511
rect 3783 2443 3839 2477
rect 3783 2409 3794 2443
rect 3828 2409 3839 2443
rect 3783 2375 3839 2409
rect 3783 2341 3794 2375
rect 3828 2341 3839 2375
rect 3783 2307 3839 2341
rect 3783 2273 3794 2307
rect 3828 2273 3839 2307
rect 3783 2239 3839 2273
rect 3783 2205 3794 2239
rect 3828 2205 3839 2239
rect 3783 2171 3839 2205
rect 3783 2137 3794 2171
rect 3828 2137 3839 2171
rect 3783 2103 3839 2137
rect 3783 2069 3794 2103
rect 3828 2069 3839 2103
rect 3783 2035 3839 2069
rect 3783 2001 3794 2035
rect 3828 2001 3839 2035
rect 3783 1967 3839 2001
rect 3783 1933 3794 1967
rect 3828 1933 3839 1967
rect 3783 1921 3839 1933
rect 3939 2851 3995 2921
rect 3939 2817 3950 2851
rect 3984 2817 3995 2851
rect 3939 2783 3995 2817
rect 3939 2749 3950 2783
rect 3984 2749 3995 2783
rect 3939 2715 3995 2749
rect 3939 2681 3950 2715
rect 3984 2681 3995 2715
rect 3939 2647 3995 2681
rect 3939 2613 3950 2647
rect 3984 2613 3995 2647
rect 3939 2579 3995 2613
rect 3939 2545 3950 2579
rect 3984 2545 3995 2579
rect 3939 2511 3995 2545
rect 3939 2477 3950 2511
rect 3984 2477 3995 2511
rect 3939 2443 3995 2477
rect 3939 2409 3950 2443
rect 3984 2409 3995 2443
rect 3939 2375 3995 2409
rect 3939 2341 3950 2375
rect 3984 2341 3995 2375
rect 3939 2307 3995 2341
rect 3939 2273 3950 2307
rect 3984 2273 3995 2307
rect 3939 2239 3995 2273
rect 3939 2205 3950 2239
rect 3984 2205 3995 2239
rect 3939 2171 3995 2205
rect 3939 2137 3950 2171
rect 3984 2137 3995 2171
rect 3939 2103 3995 2137
rect 3939 2069 3950 2103
rect 3984 2069 3995 2103
rect 3939 2035 3995 2069
rect 3939 2001 3950 2035
rect 3984 2001 3995 2035
rect 3939 1967 3995 2001
rect 3939 1933 3950 1967
rect 3984 1933 3995 1967
rect 3939 1921 3995 1933
rect 4095 2851 4148 2921
rect 4095 2817 4106 2851
rect 4140 2817 4148 2851
rect 4095 2783 4148 2817
rect 4095 2749 4106 2783
rect 4140 2749 4148 2783
rect 4095 2715 4148 2749
rect 4095 2681 4106 2715
rect 4140 2681 4148 2715
rect 4095 2647 4148 2681
rect 4095 2613 4106 2647
rect 4140 2613 4148 2647
rect 4095 2579 4148 2613
rect 4095 2545 4106 2579
rect 4140 2545 4148 2579
rect 4095 2511 4148 2545
rect 4095 2477 4106 2511
rect 4140 2477 4148 2511
rect 4095 2443 4148 2477
rect 4095 2409 4106 2443
rect 4140 2409 4148 2443
rect 4095 2375 4148 2409
rect 4095 2341 4106 2375
rect 4140 2341 4148 2375
rect 4095 2307 4148 2341
rect 4095 2273 4106 2307
rect 4140 2273 4148 2307
rect 4095 2239 4148 2273
rect 4095 2205 4106 2239
rect 4140 2205 4148 2239
rect 4095 2171 4148 2205
rect 4095 2137 4106 2171
rect 4140 2137 4148 2171
rect 4095 2103 4148 2137
rect 4095 2069 4106 2103
rect 4140 2069 4148 2103
rect 4095 2035 4148 2069
rect 4095 2001 4106 2035
rect 4140 2001 4148 2035
rect 4095 1967 4148 2001
rect 4095 1933 4106 1967
rect 4140 1933 4148 1967
rect 4095 1921 4148 1933
rect 4208 2443 4261 2521
rect 4208 2409 4216 2443
rect 4250 2409 4261 2443
rect 4208 2375 4261 2409
rect 4208 2341 4216 2375
rect 4250 2341 4261 2375
rect 4208 2307 4261 2341
rect 4208 2273 4216 2307
rect 4250 2273 4261 2307
rect 4208 2239 4261 2273
rect 4208 2205 4216 2239
rect 4250 2205 4261 2239
rect 4208 2171 4261 2205
rect 4208 2137 4216 2171
rect 4250 2137 4261 2171
rect 4208 2103 4261 2137
rect 4208 2069 4216 2103
rect 4250 2069 4261 2103
rect 4208 2035 4261 2069
rect 4208 2001 4216 2035
rect 4250 2001 4261 2035
rect 4208 1967 4261 2001
rect 4208 1933 4216 1967
rect 4250 1933 4261 1967
rect 4208 1921 4261 1933
rect 4361 2443 4417 2521
rect 4361 2409 4372 2443
rect 4406 2409 4417 2443
rect 4361 2375 4417 2409
rect 4361 2341 4372 2375
rect 4406 2341 4417 2375
rect 4361 2307 4417 2341
rect 4361 2273 4372 2307
rect 4406 2273 4417 2307
rect 4361 2239 4417 2273
rect 4361 2205 4372 2239
rect 4406 2205 4417 2239
rect 4361 2171 4417 2205
rect 4361 2137 4372 2171
rect 4406 2137 4417 2171
rect 4361 2103 4417 2137
rect 4361 2069 4372 2103
rect 4406 2069 4417 2103
rect 4361 2035 4417 2069
rect 4361 2001 4372 2035
rect 4406 2001 4417 2035
rect 4361 1967 4417 2001
rect 4361 1933 4372 1967
rect 4406 1933 4417 1967
rect 4361 1921 4417 1933
rect 4517 2443 4570 2521
rect 4517 2409 4528 2443
rect 4562 2409 4570 2443
rect 4517 2375 4570 2409
rect 4517 2341 4528 2375
rect 4562 2341 4570 2375
rect 4517 2307 4570 2341
rect 4517 2273 4528 2307
rect 4562 2273 4570 2307
rect 4517 2239 4570 2273
rect 4517 2205 4528 2239
rect 4562 2205 4570 2239
rect 4517 2171 4570 2205
rect 4517 2137 4528 2171
rect 4562 2137 4570 2171
rect 4517 2103 4570 2137
rect 4517 2069 4528 2103
rect 4562 2069 4570 2103
rect 4517 2035 4570 2069
rect 4517 2001 4528 2035
rect 4562 2001 4570 2035
rect 4517 1967 4570 2001
rect 4517 1933 4528 1967
rect 4562 1933 4570 1967
rect 4517 1921 4570 1933
rect 5494 2851 5547 2921
rect 5494 2817 5502 2851
rect 5536 2817 5547 2851
rect 5494 2783 5547 2817
rect 5494 2749 5502 2783
rect 5536 2749 5547 2783
rect 5494 2715 5547 2749
rect 5494 2681 5502 2715
rect 5536 2681 5547 2715
rect 5494 2647 5547 2681
rect 5494 2613 5502 2647
rect 5536 2613 5547 2647
rect 5494 2579 5547 2613
rect 5494 2545 5502 2579
rect 5536 2545 5547 2579
rect 5494 2511 5547 2545
rect 5494 2477 5502 2511
rect 5536 2477 5547 2511
rect 5494 2443 5547 2477
rect 5494 2409 5502 2443
rect 5536 2409 5547 2443
rect 5494 2375 5547 2409
rect 5494 2341 5502 2375
rect 5536 2341 5547 2375
rect 5494 2307 5547 2341
rect 5494 2273 5502 2307
rect 5536 2273 5547 2307
rect 5494 2239 5547 2273
rect 5494 2205 5502 2239
rect 5536 2205 5547 2239
rect 5494 2171 5547 2205
rect 5494 2137 5502 2171
rect 5536 2137 5547 2171
rect 5494 2103 5547 2137
rect 5494 2069 5502 2103
rect 5536 2069 5547 2103
rect 5494 2035 5547 2069
rect 5494 2001 5502 2035
rect 5536 2001 5547 2035
rect 5494 1967 5547 2001
rect 5494 1933 5502 1967
rect 5536 1933 5547 1967
rect 5494 1921 5547 1933
rect 5647 2851 5703 2921
rect 5647 2817 5658 2851
rect 5692 2817 5703 2851
rect 5647 2783 5703 2817
rect 5647 2749 5658 2783
rect 5692 2749 5703 2783
rect 5647 2715 5703 2749
rect 5647 2681 5658 2715
rect 5692 2681 5703 2715
rect 5647 2647 5703 2681
rect 5647 2613 5658 2647
rect 5692 2613 5703 2647
rect 5647 2579 5703 2613
rect 5647 2545 5658 2579
rect 5692 2545 5703 2579
rect 5647 2511 5703 2545
rect 5647 2477 5658 2511
rect 5692 2477 5703 2511
rect 5647 2443 5703 2477
rect 5647 2409 5658 2443
rect 5692 2409 5703 2443
rect 5647 2375 5703 2409
rect 5647 2341 5658 2375
rect 5692 2341 5703 2375
rect 5647 2307 5703 2341
rect 5647 2273 5658 2307
rect 5692 2273 5703 2307
rect 5647 2239 5703 2273
rect 5647 2205 5658 2239
rect 5692 2205 5703 2239
rect 5647 2171 5703 2205
rect 5647 2137 5658 2171
rect 5692 2137 5703 2171
rect 5647 2103 5703 2137
rect 5647 2069 5658 2103
rect 5692 2069 5703 2103
rect 5647 2035 5703 2069
rect 5647 2001 5658 2035
rect 5692 2001 5703 2035
rect 5647 1967 5703 2001
rect 5647 1933 5658 1967
rect 5692 1933 5703 1967
rect 5647 1921 5703 1933
rect 5803 2851 5859 2921
rect 5803 2817 5814 2851
rect 5848 2817 5859 2851
rect 5803 2783 5859 2817
rect 5803 2749 5814 2783
rect 5848 2749 5859 2783
rect 5803 2715 5859 2749
rect 5803 2681 5814 2715
rect 5848 2681 5859 2715
rect 5803 2647 5859 2681
rect 5803 2613 5814 2647
rect 5848 2613 5859 2647
rect 5803 2579 5859 2613
rect 5803 2545 5814 2579
rect 5848 2545 5859 2579
rect 5803 2511 5859 2545
rect 5803 2477 5814 2511
rect 5848 2477 5859 2511
rect 5803 2443 5859 2477
rect 5803 2409 5814 2443
rect 5848 2409 5859 2443
rect 5803 2375 5859 2409
rect 5803 2341 5814 2375
rect 5848 2341 5859 2375
rect 5803 2307 5859 2341
rect 5803 2273 5814 2307
rect 5848 2273 5859 2307
rect 5803 2239 5859 2273
rect 5803 2205 5814 2239
rect 5848 2205 5859 2239
rect 5803 2171 5859 2205
rect 5803 2137 5814 2171
rect 5848 2137 5859 2171
rect 5803 2103 5859 2137
rect 5803 2069 5814 2103
rect 5848 2069 5859 2103
rect 5803 2035 5859 2069
rect 5803 2001 5814 2035
rect 5848 2001 5859 2035
rect 5803 1967 5859 2001
rect 5803 1933 5814 1967
rect 5848 1933 5859 1967
rect 5803 1921 5859 1933
rect 6019 2851 6075 2921
rect 6019 2817 6030 2851
rect 6064 2817 6075 2851
rect 6019 2783 6075 2817
rect 6019 2749 6030 2783
rect 6064 2749 6075 2783
rect 6019 2715 6075 2749
rect 6019 2681 6030 2715
rect 6064 2681 6075 2715
rect 6019 2647 6075 2681
rect 6019 2613 6030 2647
rect 6064 2613 6075 2647
rect 6019 2579 6075 2613
rect 6019 2545 6030 2579
rect 6064 2545 6075 2579
rect 6019 2511 6075 2545
rect 6019 2477 6030 2511
rect 6064 2477 6075 2511
rect 6019 2443 6075 2477
rect 6019 2409 6030 2443
rect 6064 2409 6075 2443
rect 6019 2375 6075 2409
rect 6019 2341 6030 2375
rect 6064 2341 6075 2375
rect 6019 2307 6075 2341
rect 6019 2273 6030 2307
rect 6064 2273 6075 2307
rect 6019 2239 6075 2273
rect 6019 2205 6030 2239
rect 6064 2205 6075 2239
rect 6019 2171 6075 2205
rect 6019 2137 6030 2171
rect 6064 2137 6075 2171
rect 6019 2103 6075 2137
rect 6019 2069 6030 2103
rect 6064 2069 6075 2103
rect 6019 2035 6075 2069
rect 6019 2001 6030 2035
rect 6064 2001 6075 2035
rect 6019 1967 6075 2001
rect 6019 1933 6030 1967
rect 6064 1933 6075 1967
rect 6019 1921 6075 1933
rect 6235 2851 6288 2921
rect 6235 2817 6246 2851
rect 6280 2817 6288 2851
rect 6235 2783 6288 2817
rect 6235 2749 6246 2783
rect 6280 2749 6288 2783
rect 6235 2715 6288 2749
rect 6235 2681 6246 2715
rect 6280 2681 6288 2715
rect 6235 2647 6288 2681
rect 6235 2613 6246 2647
rect 6280 2613 6288 2647
rect 6235 2579 6288 2613
rect 6235 2545 6246 2579
rect 6280 2545 6288 2579
rect 6235 2511 6288 2545
rect 6235 2477 6246 2511
rect 6280 2477 6288 2511
rect 6235 2443 6288 2477
rect 6235 2409 6246 2443
rect 6280 2409 6288 2443
rect 6235 2375 6288 2409
rect 6235 2341 6246 2375
rect 6280 2341 6288 2375
rect 6235 2307 6288 2341
rect 6348 2503 6401 2521
rect 6348 2469 6356 2503
rect 6390 2469 6401 2503
rect 6348 2435 6401 2469
rect 6348 2401 6356 2435
rect 6390 2401 6401 2435
rect 6348 2367 6401 2401
rect 6348 2333 6356 2367
rect 6390 2333 6401 2367
rect 6348 2321 6401 2333
rect 6501 2503 6554 2521
rect 6501 2469 6512 2503
rect 6546 2469 6554 2503
rect 6501 2435 6554 2469
rect 6501 2401 6512 2435
rect 6546 2401 6554 2435
rect 6501 2367 6554 2401
rect 6501 2333 6512 2367
rect 6546 2333 6554 2367
rect 6501 2321 6554 2333
rect 6235 2273 6246 2307
rect 6280 2273 6288 2307
rect 6235 2239 6288 2273
rect 6235 2205 6246 2239
rect 6280 2205 6288 2239
rect 6235 2171 6288 2205
rect 6235 2137 6246 2171
rect 6280 2137 6288 2171
rect 6235 2103 6288 2137
rect 6235 2069 6246 2103
rect 6280 2069 6288 2103
rect 6235 2035 6288 2069
rect 6235 2001 6246 2035
rect 6280 2001 6288 2035
rect 6235 1967 6288 2001
rect 6235 1933 6246 1967
rect 6280 1933 6288 1967
rect 6235 1921 6288 1933
rect 7362 2851 7415 2921
rect 7362 2817 7370 2851
rect 7404 2817 7415 2851
rect 7362 2783 7415 2817
rect 7362 2749 7370 2783
rect 7404 2749 7415 2783
rect 7362 2715 7415 2749
rect 7362 2681 7370 2715
rect 7404 2681 7415 2715
rect 7362 2647 7415 2681
rect 7362 2613 7370 2647
rect 7404 2613 7415 2647
rect 7362 2579 7415 2613
rect 7362 2545 7370 2579
rect 7404 2545 7415 2579
rect 7362 2511 7415 2545
rect 7362 2477 7370 2511
rect 7404 2477 7415 2511
rect 7362 2443 7415 2477
rect 7362 2409 7370 2443
rect 7404 2409 7415 2443
rect 7362 2375 7415 2409
rect 7362 2341 7370 2375
rect 7404 2341 7415 2375
rect 7362 2307 7415 2341
rect 7362 2273 7370 2307
rect 7404 2273 7415 2307
rect 7362 2239 7415 2273
rect 7362 2205 7370 2239
rect 7404 2205 7415 2239
rect 7362 2171 7415 2205
rect 7362 2137 7370 2171
rect 7404 2137 7415 2171
rect 7362 2103 7415 2137
rect 7362 2069 7370 2103
rect 7404 2069 7415 2103
rect 7362 2035 7415 2069
rect 7362 2001 7370 2035
rect 7404 2001 7415 2035
rect 7362 1967 7415 2001
rect 7362 1933 7370 1967
rect 7404 1933 7415 1967
rect 7362 1921 7415 1933
rect 7575 2851 7631 2921
rect 7575 2817 7586 2851
rect 7620 2817 7631 2851
rect 7575 2783 7631 2817
rect 7575 2749 7586 2783
rect 7620 2749 7631 2783
rect 7575 2715 7631 2749
rect 7575 2681 7586 2715
rect 7620 2681 7631 2715
rect 7575 2647 7631 2681
rect 7575 2613 7586 2647
rect 7620 2613 7631 2647
rect 7575 2579 7631 2613
rect 7575 2545 7586 2579
rect 7620 2545 7631 2579
rect 7575 2511 7631 2545
rect 7575 2477 7586 2511
rect 7620 2477 7631 2511
rect 7575 2443 7631 2477
rect 7575 2409 7586 2443
rect 7620 2409 7631 2443
rect 7575 2375 7631 2409
rect 7575 2341 7586 2375
rect 7620 2341 7631 2375
rect 7575 2307 7631 2341
rect 7575 2273 7586 2307
rect 7620 2273 7631 2307
rect 7575 2239 7631 2273
rect 7575 2205 7586 2239
rect 7620 2205 7631 2239
rect 7575 2171 7631 2205
rect 7575 2137 7586 2171
rect 7620 2137 7631 2171
rect 7575 2103 7631 2137
rect 7575 2069 7586 2103
rect 7620 2069 7631 2103
rect 7575 2035 7631 2069
rect 7575 2001 7586 2035
rect 7620 2001 7631 2035
rect 7575 1967 7631 2001
rect 7575 1933 7586 1967
rect 7620 1933 7631 1967
rect 7575 1921 7631 1933
rect 7791 2851 7847 2921
rect 7791 2817 7802 2851
rect 7836 2817 7847 2851
rect 7791 2783 7847 2817
rect 7791 2749 7802 2783
rect 7836 2749 7847 2783
rect 7791 2715 7847 2749
rect 7791 2681 7802 2715
rect 7836 2681 7847 2715
rect 7791 2647 7847 2681
rect 7791 2613 7802 2647
rect 7836 2613 7847 2647
rect 7791 2579 7847 2613
rect 7791 2545 7802 2579
rect 7836 2545 7847 2579
rect 7791 2511 7847 2545
rect 7791 2477 7802 2511
rect 7836 2477 7847 2511
rect 7791 2443 7847 2477
rect 7791 2409 7802 2443
rect 7836 2409 7847 2443
rect 7791 2375 7847 2409
rect 7791 2341 7802 2375
rect 7836 2341 7847 2375
rect 7791 2307 7847 2341
rect 7791 2273 7802 2307
rect 7836 2273 7847 2307
rect 7791 2239 7847 2273
rect 7791 2205 7802 2239
rect 7836 2205 7847 2239
rect 7791 2171 7847 2205
rect 7791 2137 7802 2171
rect 7836 2137 7847 2171
rect 7791 2103 7847 2137
rect 7791 2069 7802 2103
rect 7836 2069 7847 2103
rect 7791 2035 7847 2069
rect 7791 2001 7802 2035
rect 7836 2001 7847 2035
rect 7791 1967 7847 2001
rect 7791 1933 7802 1967
rect 7836 1933 7847 1967
rect 7791 1921 7847 1933
rect 8007 2851 8063 2921
rect 8007 2817 8018 2851
rect 8052 2817 8063 2851
rect 8007 2783 8063 2817
rect 8007 2749 8018 2783
rect 8052 2749 8063 2783
rect 8007 2715 8063 2749
rect 8007 2681 8018 2715
rect 8052 2681 8063 2715
rect 8007 2647 8063 2681
rect 8007 2613 8018 2647
rect 8052 2613 8063 2647
rect 8007 2579 8063 2613
rect 8007 2545 8018 2579
rect 8052 2545 8063 2579
rect 8007 2511 8063 2545
rect 8007 2477 8018 2511
rect 8052 2477 8063 2511
rect 8007 2443 8063 2477
rect 8007 2409 8018 2443
rect 8052 2409 8063 2443
rect 8007 2375 8063 2409
rect 8007 2341 8018 2375
rect 8052 2341 8063 2375
rect 8007 2307 8063 2341
rect 8007 2273 8018 2307
rect 8052 2273 8063 2307
rect 8007 2239 8063 2273
rect 8007 2205 8018 2239
rect 8052 2205 8063 2239
rect 8007 2171 8063 2205
rect 8007 2137 8018 2171
rect 8052 2137 8063 2171
rect 8007 2103 8063 2137
rect 8007 2069 8018 2103
rect 8052 2069 8063 2103
rect 8007 2035 8063 2069
rect 8007 2001 8018 2035
rect 8052 2001 8063 2035
rect 8007 1967 8063 2001
rect 8007 1933 8018 1967
rect 8052 1933 8063 1967
rect 8007 1921 8063 1933
rect 8163 2851 8219 2921
rect 8163 2817 8174 2851
rect 8208 2817 8219 2851
rect 8163 2783 8219 2817
rect 8163 2749 8174 2783
rect 8208 2749 8219 2783
rect 8163 2715 8219 2749
rect 8163 2681 8174 2715
rect 8208 2681 8219 2715
rect 8163 2647 8219 2681
rect 8163 2613 8174 2647
rect 8208 2613 8219 2647
rect 8163 2579 8219 2613
rect 8163 2545 8174 2579
rect 8208 2545 8219 2579
rect 8163 2511 8219 2545
rect 8163 2477 8174 2511
rect 8208 2477 8219 2511
rect 8163 2443 8219 2477
rect 8163 2409 8174 2443
rect 8208 2409 8219 2443
rect 8163 2375 8219 2409
rect 8163 2341 8174 2375
rect 8208 2341 8219 2375
rect 8163 2307 8219 2341
rect 8163 2273 8174 2307
rect 8208 2273 8219 2307
rect 8163 2239 8219 2273
rect 8163 2205 8174 2239
rect 8208 2205 8219 2239
rect 8163 2171 8219 2205
rect 8163 2137 8174 2171
rect 8208 2137 8219 2171
rect 8163 2103 8219 2137
rect 8163 2069 8174 2103
rect 8208 2069 8219 2103
rect 8163 2035 8219 2069
rect 8163 2001 8174 2035
rect 8208 2001 8219 2035
rect 8163 1967 8219 2001
rect 8163 1933 8174 1967
rect 8208 1933 8219 1967
rect 8163 1921 8219 1933
rect 8319 2851 8375 2921
rect 8319 2817 8330 2851
rect 8364 2817 8375 2851
rect 8319 2783 8375 2817
rect 8319 2749 8330 2783
rect 8364 2749 8375 2783
rect 8319 2715 8375 2749
rect 8319 2681 8330 2715
rect 8364 2681 8375 2715
rect 8319 2647 8375 2681
rect 8319 2613 8330 2647
rect 8364 2613 8375 2647
rect 8319 2579 8375 2613
rect 8319 2545 8330 2579
rect 8364 2545 8375 2579
rect 8319 2511 8375 2545
rect 8319 2477 8330 2511
rect 8364 2477 8375 2511
rect 8319 2443 8375 2477
rect 8319 2409 8330 2443
rect 8364 2409 8375 2443
rect 8319 2375 8375 2409
rect 8319 2341 8330 2375
rect 8364 2341 8375 2375
rect 8319 2307 8375 2341
rect 8319 2273 8330 2307
rect 8364 2273 8375 2307
rect 8319 2239 8375 2273
rect 8319 2205 8330 2239
rect 8364 2205 8375 2239
rect 8319 2171 8375 2205
rect 8319 2137 8330 2171
rect 8364 2137 8375 2171
rect 8319 2103 8375 2137
rect 8319 2069 8330 2103
rect 8364 2069 8375 2103
rect 8319 2035 8375 2069
rect 8319 2001 8330 2035
rect 8364 2001 8375 2035
rect 8319 1967 8375 2001
rect 8319 1933 8330 1967
rect 8364 1933 8375 1967
rect 8319 1921 8375 1933
rect 8475 2851 8531 2921
rect 8475 2817 8486 2851
rect 8520 2817 8531 2851
rect 8475 2783 8531 2817
rect 8475 2749 8486 2783
rect 8520 2749 8531 2783
rect 8475 2715 8531 2749
rect 8475 2681 8486 2715
rect 8520 2681 8531 2715
rect 8475 2647 8531 2681
rect 8475 2613 8486 2647
rect 8520 2613 8531 2647
rect 8475 2579 8531 2613
rect 8475 2545 8486 2579
rect 8520 2545 8531 2579
rect 8475 2511 8531 2545
rect 8475 2477 8486 2511
rect 8520 2477 8531 2511
rect 8475 2443 8531 2477
rect 8475 2409 8486 2443
rect 8520 2409 8531 2443
rect 8475 2375 8531 2409
rect 8475 2341 8486 2375
rect 8520 2341 8531 2375
rect 8475 2307 8531 2341
rect 8475 2273 8486 2307
rect 8520 2273 8531 2307
rect 8475 2239 8531 2273
rect 8475 2205 8486 2239
rect 8520 2205 8531 2239
rect 8475 2171 8531 2205
rect 8475 2137 8486 2171
rect 8520 2137 8531 2171
rect 8475 2103 8531 2137
rect 8475 2069 8486 2103
rect 8520 2069 8531 2103
rect 8475 2035 8531 2069
rect 8475 2001 8486 2035
rect 8520 2001 8531 2035
rect 8475 1967 8531 2001
rect 8475 1933 8486 1967
rect 8520 1933 8531 1967
rect 8475 1921 8531 1933
rect 8631 2851 8684 2921
rect 8631 2817 8642 2851
rect 8676 2817 8684 2851
rect 8631 2783 8684 2817
rect 8631 2749 8642 2783
rect 8676 2749 8684 2783
rect 8631 2715 8684 2749
rect 8631 2681 8642 2715
rect 8676 2681 8684 2715
rect 8631 2647 8684 2681
rect 8631 2613 8642 2647
rect 8676 2613 8684 2647
rect 8631 2579 8684 2613
rect 8631 2545 8642 2579
rect 8676 2545 8684 2579
rect 8631 2511 8684 2545
rect 8631 2477 8642 2511
rect 8676 2477 8684 2511
rect 8631 2443 8684 2477
rect 8631 2409 8642 2443
rect 8676 2409 8684 2443
rect 8631 2375 8684 2409
rect 8631 2341 8642 2375
rect 8676 2341 8684 2375
rect 8631 2307 8684 2341
rect 8631 2273 8642 2307
rect 8676 2273 8684 2307
rect 8631 2239 8684 2273
rect 8631 2205 8642 2239
rect 8676 2205 8684 2239
rect 8631 2171 8684 2205
rect 8631 2137 8642 2171
rect 8676 2137 8684 2171
rect 8631 2103 8684 2137
rect 8631 2069 8642 2103
rect 8676 2069 8684 2103
rect 8631 2035 8684 2069
rect 8631 2001 8642 2035
rect 8676 2001 8684 2035
rect 8631 1967 8684 2001
rect 8631 1933 8642 1967
rect 8676 1933 8684 1967
rect 8631 1921 8684 1933
rect 9640 2851 9693 2921
rect 9640 2817 9648 2851
rect 9682 2817 9693 2851
rect 9640 2783 9693 2817
rect 9640 2749 9648 2783
rect 9682 2749 9693 2783
rect 9640 2715 9693 2749
rect 9640 2681 9648 2715
rect 9682 2681 9693 2715
rect 9640 2647 9693 2681
rect 9640 2613 9648 2647
rect 9682 2613 9693 2647
rect 9640 2579 9693 2613
rect 9640 2545 9648 2579
rect 9682 2545 9693 2579
rect 9640 2511 9693 2545
rect 9640 2477 9648 2511
rect 9682 2477 9693 2511
rect 9640 2443 9693 2477
rect 9640 2409 9648 2443
rect 9682 2409 9693 2443
rect 9640 2375 9693 2409
rect 9640 2341 9648 2375
rect 9682 2341 9693 2375
rect 9640 2307 9693 2341
rect 9640 2273 9648 2307
rect 9682 2273 9693 2307
rect 9640 2239 9693 2273
rect 9640 2205 9648 2239
rect 9682 2205 9693 2239
rect 9640 2171 9693 2205
rect 9640 2137 9648 2171
rect 9682 2137 9693 2171
rect 9640 2103 9693 2137
rect 9640 2069 9648 2103
rect 9682 2069 9693 2103
rect 9640 2035 9693 2069
rect 9640 2001 9648 2035
rect 9682 2001 9693 2035
rect 9640 1967 9693 2001
rect 9640 1933 9648 1967
rect 9682 1933 9693 1967
rect 9640 1921 9693 1933
rect 9793 2851 9849 2921
rect 9793 2817 9804 2851
rect 9838 2817 9849 2851
rect 9793 2783 9849 2817
rect 9793 2749 9804 2783
rect 9838 2749 9849 2783
rect 9793 2715 9849 2749
rect 9793 2681 9804 2715
rect 9838 2681 9849 2715
rect 9793 2647 9849 2681
rect 9793 2613 9804 2647
rect 9838 2613 9849 2647
rect 9793 2579 9849 2613
rect 9793 2545 9804 2579
rect 9838 2545 9849 2579
rect 9793 2511 9849 2545
rect 9793 2477 9804 2511
rect 9838 2477 9849 2511
rect 9793 2443 9849 2477
rect 9793 2409 9804 2443
rect 9838 2409 9849 2443
rect 9793 2375 9849 2409
rect 9793 2341 9804 2375
rect 9838 2341 9849 2375
rect 9793 2307 9849 2341
rect 9793 2273 9804 2307
rect 9838 2273 9849 2307
rect 9793 2239 9849 2273
rect 9793 2205 9804 2239
rect 9838 2205 9849 2239
rect 9793 2171 9849 2205
rect 9793 2137 9804 2171
rect 9838 2137 9849 2171
rect 9793 2103 9849 2137
rect 9793 2069 9804 2103
rect 9838 2069 9849 2103
rect 9793 2035 9849 2069
rect 9793 2001 9804 2035
rect 9838 2001 9849 2035
rect 9793 1967 9849 2001
rect 9793 1933 9804 1967
rect 9838 1933 9849 1967
rect 9793 1921 9849 1933
rect 9949 2851 10005 2921
rect 9949 2817 9960 2851
rect 9994 2817 10005 2851
rect 9949 2783 10005 2817
rect 9949 2749 9960 2783
rect 9994 2749 10005 2783
rect 9949 2715 10005 2749
rect 9949 2681 9960 2715
rect 9994 2681 10005 2715
rect 9949 2647 10005 2681
rect 9949 2613 9960 2647
rect 9994 2613 10005 2647
rect 9949 2579 10005 2613
rect 9949 2545 9960 2579
rect 9994 2545 10005 2579
rect 9949 2511 10005 2545
rect 9949 2477 9960 2511
rect 9994 2477 10005 2511
rect 9949 2443 10005 2477
rect 9949 2409 9960 2443
rect 9994 2409 10005 2443
rect 9949 2375 10005 2409
rect 9949 2341 9960 2375
rect 9994 2341 10005 2375
rect 9949 2307 10005 2341
rect 9949 2273 9960 2307
rect 9994 2273 10005 2307
rect 9949 2239 10005 2273
rect 9949 2205 9960 2239
rect 9994 2205 10005 2239
rect 9949 2171 10005 2205
rect 9949 2137 9960 2171
rect 9994 2137 10005 2171
rect 9949 2103 10005 2137
rect 9949 2069 9960 2103
rect 9994 2069 10005 2103
rect 9949 2035 10005 2069
rect 9949 2001 9960 2035
rect 9994 2001 10005 2035
rect 9949 1967 10005 2001
rect 9949 1933 9960 1967
rect 9994 1933 10005 1967
rect 9949 1921 10005 1933
rect 10105 2851 10161 2921
rect 10105 2817 10116 2851
rect 10150 2817 10161 2851
rect 10105 2783 10161 2817
rect 10105 2749 10116 2783
rect 10150 2749 10161 2783
rect 10105 2715 10161 2749
rect 10105 2681 10116 2715
rect 10150 2681 10161 2715
rect 10105 2647 10161 2681
rect 10105 2613 10116 2647
rect 10150 2613 10161 2647
rect 10105 2579 10161 2613
rect 10105 2545 10116 2579
rect 10150 2545 10161 2579
rect 10105 2511 10161 2545
rect 10105 2477 10116 2511
rect 10150 2477 10161 2511
rect 10105 2443 10161 2477
rect 10105 2409 10116 2443
rect 10150 2409 10161 2443
rect 10105 2375 10161 2409
rect 10105 2341 10116 2375
rect 10150 2341 10161 2375
rect 10105 2307 10161 2341
rect 10105 2273 10116 2307
rect 10150 2273 10161 2307
rect 10105 2239 10161 2273
rect 10105 2205 10116 2239
rect 10150 2205 10161 2239
rect 10105 2171 10161 2205
rect 10105 2137 10116 2171
rect 10150 2137 10161 2171
rect 10105 2103 10161 2137
rect 10105 2069 10116 2103
rect 10150 2069 10161 2103
rect 10105 2035 10161 2069
rect 10105 2001 10116 2035
rect 10150 2001 10161 2035
rect 10105 1967 10161 2001
rect 10105 1933 10116 1967
rect 10150 1933 10161 1967
rect 10105 1921 10161 1933
rect 10261 2851 10317 2921
rect 10261 2817 10272 2851
rect 10306 2817 10317 2851
rect 10261 2783 10317 2817
rect 10261 2749 10272 2783
rect 10306 2749 10317 2783
rect 10261 2715 10317 2749
rect 10261 2681 10272 2715
rect 10306 2681 10317 2715
rect 10261 2647 10317 2681
rect 10261 2613 10272 2647
rect 10306 2613 10317 2647
rect 10261 2579 10317 2613
rect 10261 2545 10272 2579
rect 10306 2545 10317 2579
rect 10261 2511 10317 2545
rect 10261 2477 10272 2511
rect 10306 2477 10317 2511
rect 10261 2443 10317 2477
rect 10261 2409 10272 2443
rect 10306 2409 10317 2443
rect 10261 2375 10317 2409
rect 10261 2341 10272 2375
rect 10306 2341 10317 2375
rect 10261 2307 10317 2341
rect 10261 2273 10272 2307
rect 10306 2273 10317 2307
rect 10261 2239 10317 2273
rect 10261 2205 10272 2239
rect 10306 2205 10317 2239
rect 10261 2171 10317 2205
rect 10261 2137 10272 2171
rect 10306 2137 10317 2171
rect 10261 2103 10317 2137
rect 10261 2069 10272 2103
rect 10306 2069 10317 2103
rect 10261 2035 10317 2069
rect 10261 2001 10272 2035
rect 10306 2001 10317 2035
rect 10261 1967 10317 2001
rect 10261 1933 10272 1967
rect 10306 1933 10317 1967
rect 10261 1921 10317 1933
rect 10417 2851 10473 2921
rect 10417 2817 10428 2851
rect 10462 2817 10473 2851
rect 10417 2783 10473 2817
rect 10417 2749 10428 2783
rect 10462 2749 10473 2783
rect 10417 2715 10473 2749
rect 10417 2681 10428 2715
rect 10462 2681 10473 2715
rect 10417 2647 10473 2681
rect 10417 2613 10428 2647
rect 10462 2613 10473 2647
rect 10417 2579 10473 2613
rect 10417 2545 10428 2579
rect 10462 2545 10473 2579
rect 10417 2511 10473 2545
rect 10417 2477 10428 2511
rect 10462 2477 10473 2511
rect 10417 2443 10473 2477
rect 10417 2409 10428 2443
rect 10462 2409 10473 2443
rect 10417 2375 10473 2409
rect 10417 2341 10428 2375
rect 10462 2341 10473 2375
rect 10417 2307 10473 2341
rect 10417 2273 10428 2307
rect 10462 2273 10473 2307
rect 10417 2239 10473 2273
rect 10417 2205 10428 2239
rect 10462 2205 10473 2239
rect 10417 2171 10473 2205
rect 10417 2137 10428 2171
rect 10462 2137 10473 2171
rect 10417 2103 10473 2137
rect 10417 2069 10428 2103
rect 10462 2069 10473 2103
rect 10417 2035 10473 2069
rect 10417 2001 10428 2035
rect 10462 2001 10473 2035
rect 10417 1967 10473 2001
rect 10417 1933 10428 1967
rect 10462 1933 10473 1967
rect 10417 1921 10473 1933
rect 10573 2851 10629 2921
rect 10573 2817 10584 2851
rect 10618 2817 10629 2851
rect 10573 2783 10629 2817
rect 10573 2749 10584 2783
rect 10618 2749 10629 2783
rect 10573 2715 10629 2749
rect 10573 2681 10584 2715
rect 10618 2681 10629 2715
rect 10573 2647 10629 2681
rect 10573 2613 10584 2647
rect 10618 2613 10629 2647
rect 10573 2579 10629 2613
rect 10573 2545 10584 2579
rect 10618 2545 10629 2579
rect 10573 2511 10629 2545
rect 10573 2477 10584 2511
rect 10618 2477 10629 2511
rect 10573 2443 10629 2477
rect 10573 2409 10584 2443
rect 10618 2409 10629 2443
rect 10573 2375 10629 2409
rect 10573 2341 10584 2375
rect 10618 2341 10629 2375
rect 10573 2307 10629 2341
rect 10573 2273 10584 2307
rect 10618 2273 10629 2307
rect 10573 2239 10629 2273
rect 10573 2205 10584 2239
rect 10618 2205 10629 2239
rect 10573 2171 10629 2205
rect 10573 2137 10584 2171
rect 10618 2137 10629 2171
rect 10573 2103 10629 2137
rect 10573 2069 10584 2103
rect 10618 2069 10629 2103
rect 10573 2035 10629 2069
rect 10573 2001 10584 2035
rect 10618 2001 10629 2035
rect 10573 1967 10629 2001
rect 10573 1933 10584 1967
rect 10618 1933 10629 1967
rect 10573 1921 10629 1933
rect 10729 2851 10785 2921
rect 10729 2817 10740 2851
rect 10774 2817 10785 2851
rect 10729 2783 10785 2817
rect 10729 2749 10740 2783
rect 10774 2749 10785 2783
rect 10729 2715 10785 2749
rect 10729 2681 10740 2715
rect 10774 2681 10785 2715
rect 10729 2647 10785 2681
rect 10729 2613 10740 2647
rect 10774 2613 10785 2647
rect 10729 2579 10785 2613
rect 10729 2545 10740 2579
rect 10774 2545 10785 2579
rect 10729 2511 10785 2545
rect 10729 2477 10740 2511
rect 10774 2477 10785 2511
rect 10729 2443 10785 2477
rect 10729 2409 10740 2443
rect 10774 2409 10785 2443
rect 10729 2375 10785 2409
rect 10729 2341 10740 2375
rect 10774 2341 10785 2375
rect 10729 2307 10785 2341
rect 10729 2273 10740 2307
rect 10774 2273 10785 2307
rect 10729 2239 10785 2273
rect 10729 2205 10740 2239
rect 10774 2205 10785 2239
rect 10729 2171 10785 2205
rect 10729 2137 10740 2171
rect 10774 2137 10785 2171
rect 10729 2103 10785 2137
rect 10729 2069 10740 2103
rect 10774 2069 10785 2103
rect 10729 2035 10785 2069
rect 10729 2001 10740 2035
rect 10774 2001 10785 2035
rect 10729 1967 10785 2001
rect 10729 1933 10740 1967
rect 10774 1933 10785 1967
rect 10729 1921 10785 1933
rect 10885 2851 10941 2921
rect 10885 2817 10896 2851
rect 10930 2817 10941 2851
rect 10885 2783 10941 2817
rect 10885 2749 10896 2783
rect 10930 2749 10941 2783
rect 10885 2715 10941 2749
rect 10885 2681 10896 2715
rect 10930 2681 10941 2715
rect 10885 2647 10941 2681
rect 10885 2613 10896 2647
rect 10930 2613 10941 2647
rect 10885 2579 10941 2613
rect 10885 2545 10896 2579
rect 10930 2545 10941 2579
rect 10885 2511 10941 2545
rect 10885 2477 10896 2511
rect 10930 2477 10941 2511
rect 10885 2443 10941 2477
rect 10885 2409 10896 2443
rect 10930 2409 10941 2443
rect 10885 2375 10941 2409
rect 10885 2341 10896 2375
rect 10930 2341 10941 2375
rect 10885 2307 10941 2341
rect 10885 2273 10896 2307
rect 10930 2273 10941 2307
rect 10885 2239 10941 2273
rect 10885 2205 10896 2239
rect 10930 2205 10941 2239
rect 10885 2171 10941 2205
rect 10885 2137 10896 2171
rect 10930 2137 10941 2171
rect 10885 2103 10941 2137
rect 10885 2069 10896 2103
rect 10930 2069 10941 2103
rect 10885 2035 10941 2069
rect 10885 2001 10896 2035
rect 10930 2001 10941 2035
rect 10885 1967 10941 2001
rect 10885 1933 10896 1967
rect 10930 1933 10941 1967
rect 10885 1921 10941 1933
rect 11041 2851 11097 2921
rect 11041 2817 11052 2851
rect 11086 2817 11097 2851
rect 11041 2783 11097 2817
rect 11041 2749 11052 2783
rect 11086 2749 11097 2783
rect 11041 2715 11097 2749
rect 11041 2681 11052 2715
rect 11086 2681 11097 2715
rect 11041 2647 11097 2681
rect 11041 2613 11052 2647
rect 11086 2613 11097 2647
rect 11041 2579 11097 2613
rect 11041 2545 11052 2579
rect 11086 2545 11097 2579
rect 11041 2511 11097 2545
rect 11041 2477 11052 2511
rect 11086 2477 11097 2511
rect 11041 2443 11097 2477
rect 11041 2409 11052 2443
rect 11086 2409 11097 2443
rect 11041 2375 11097 2409
rect 11041 2341 11052 2375
rect 11086 2341 11097 2375
rect 11041 2307 11097 2341
rect 11041 2273 11052 2307
rect 11086 2273 11097 2307
rect 11041 2239 11097 2273
rect 11041 2205 11052 2239
rect 11086 2205 11097 2239
rect 11041 2171 11097 2205
rect 11041 2137 11052 2171
rect 11086 2137 11097 2171
rect 11041 2103 11097 2137
rect 11041 2069 11052 2103
rect 11086 2069 11097 2103
rect 11041 2035 11097 2069
rect 11041 2001 11052 2035
rect 11086 2001 11097 2035
rect 11041 1967 11097 2001
rect 11041 1933 11052 1967
rect 11086 1933 11097 1967
rect 11041 1921 11097 1933
rect 11197 2851 11253 2921
rect 11197 2817 11208 2851
rect 11242 2817 11253 2851
rect 11197 2783 11253 2817
rect 11197 2749 11208 2783
rect 11242 2749 11253 2783
rect 11197 2715 11253 2749
rect 11197 2681 11208 2715
rect 11242 2681 11253 2715
rect 11197 2647 11253 2681
rect 11197 2613 11208 2647
rect 11242 2613 11253 2647
rect 11197 2579 11253 2613
rect 11197 2545 11208 2579
rect 11242 2545 11253 2579
rect 11197 2511 11253 2545
rect 11197 2477 11208 2511
rect 11242 2477 11253 2511
rect 11197 2443 11253 2477
rect 11197 2409 11208 2443
rect 11242 2409 11253 2443
rect 11197 2375 11253 2409
rect 11197 2341 11208 2375
rect 11242 2341 11253 2375
rect 11197 2307 11253 2341
rect 11197 2273 11208 2307
rect 11242 2273 11253 2307
rect 11197 2239 11253 2273
rect 11197 2205 11208 2239
rect 11242 2205 11253 2239
rect 11197 2171 11253 2205
rect 11197 2137 11208 2171
rect 11242 2137 11253 2171
rect 11197 2103 11253 2137
rect 11197 2069 11208 2103
rect 11242 2069 11253 2103
rect 11197 2035 11253 2069
rect 11197 2001 11208 2035
rect 11242 2001 11253 2035
rect 11197 1967 11253 2001
rect 11197 1933 11208 1967
rect 11242 1933 11253 1967
rect 11197 1921 11253 1933
rect 11353 2851 11409 2921
rect 11353 2817 11364 2851
rect 11398 2817 11409 2851
rect 11353 2783 11409 2817
rect 11353 2749 11364 2783
rect 11398 2749 11409 2783
rect 11353 2715 11409 2749
rect 11353 2681 11364 2715
rect 11398 2681 11409 2715
rect 11353 2647 11409 2681
rect 11353 2613 11364 2647
rect 11398 2613 11409 2647
rect 11353 2579 11409 2613
rect 11353 2545 11364 2579
rect 11398 2545 11409 2579
rect 11353 2511 11409 2545
rect 11353 2477 11364 2511
rect 11398 2477 11409 2511
rect 11353 2443 11409 2477
rect 11353 2409 11364 2443
rect 11398 2409 11409 2443
rect 11353 2375 11409 2409
rect 11353 2341 11364 2375
rect 11398 2341 11409 2375
rect 11353 2307 11409 2341
rect 11353 2273 11364 2307
rect 11398 2273 11409 2307
rect 11353 2239 11409 2273
rect 11353 2205 11364 2239
rect 11398 2205 11409 2239
rect 11353 2171 11409 2205
rect 11353 2137 11364 2171
rect 11398 2137 11409 2171
rect 11353 2103 11409 2137
rect 11353 2069 11364 2103
rect 11398 2069 11409 2103
rect 11353 2035 11409 2069
rect 11353 2001 11364 2035
rect 11398 2001 11409 2035
rect 11353 1967 11409 2001
rect 11353 1933 11364 1967
rect 11398 1933 11409 1967
rect 11353 1921 11409 1933
rect 11509 2851 11562 2921
rect 11509 2817 11520 2851
rect 11554 2817 11562 2851
rect 11509 2783 11562 2817
rect 11509 2749 11520 2783
rect 11554 2749 11562 2783
rect 11509 2715 11562 2749
rect 11509 2681 11520 2715
rect 11554 2681 11562 2715
rect 11509 2647 11562 2681
rect 11509 2613 11520 2647
rect 11554 2613 11562 2647
rect 11509 2579 11562 2613
rect 11509 2545 11520 2579
rect 11554 2545 11562 2579
rect 11509 2511 11562 2545
rect 11509 2477 11520 2511
rect 11554 2477 11562 2511
rect 11509 2443 11562 2477
rect 11509 2409 11520 2443
rect 11554 2409 11562 2443
rect 11509 2375 11562 2409
rect 11509 2341 11520 2375
rect 11554 2341 11562 2375
rect 11509 2307 11562 2341
rect 11509 2273 11520 2307
rect 11554 2273 11562 2307
rect 11509 2239 11562 2273
rect 11509 2205 11520 2239
rect 11554 2205 11562 2239
rect 11509 2171 11562 2205
rect 11509 2137 11520 2171
rect 11554 2137 11562 2171
rect 11509 2103 11562 2137
rect 11509 2069 11520 2103
rect 11554 2069 11562 2103
rect 11509 2035 11562 2069
rect 11509 2001 11520 2035
rect 11554 2001 11562 2035
rect 11509 1967 11562 2001
rect 11509 1933 11520 1967
rect 11554 1933 11562 1967
rect 11509 1921 11562 1933
<< pdiffc >>
rect 3942 1044 3976 1078
rect 3942 976 3976 1010
rect 3942 908 3976 942
rect 3942 840 3976 874
rect 3942 772 3976 806
rect 3942 704 3976 738
rect 3942 636 3976 670
rect 3942 568 3976 602
rect 3942 500 3976 534
rect 3942 432 3976 466
rect 3942 364 3976 398
rect 3942 296 3976 330
rect 3942 228 3976 262
rect 3942 160 3976 194
rect 4048 1044 4082 1078
rect 4048 976 4082 1010
rect 4048 908 4082 942
rect 4048 840 4082 874
rect 4048 772 4082 806
rect 4048 704 4082 738
rect 4048 636 4082 670
rect 4048 568 4082 602
rect 4048 500 4082 534
rect 4048 432 4082 466
rect 4048 364 4082 398
rect 4048 296 4082 330
rect 4048 228 4082 262
rect 4048 160 4082 194
rect 4154 1044 4188 1078
rect 4154 976 4188 1010
rect 4154 908 4188 942
rect 4154 840 4188 874
rect 4154 772 4188 806
rect 4154 704 4188 738
rect 4154 636 4188 670
rect 4154 568 4188 602
rect 4154 500 4188 534
rect 4154 432 4188 466
rect 4154 364 4188 398
rect 4154 296 4188 330
rect 4154 228 4188 262
rect 4154 160 4188 194
rect 4260 1044 4294 1078
rect 4260 976 4294 1010
rect 4260 908 4294 942
rect 4260 840 4294 874
rect 4260 772 4294 806
rect 4260 704 4294 738
rect 4260 636 4294 670
rect 4260 568 4294 602
rect 4260 500 4294 534
rect 4260 432 4294 466
rect 4260 364 4294 398
rect 4260 296 4294 330
rect 4260 228 4294 262
rect 4260 160 4294 194
rect 4366 1044 4400 1078
rect 4366 976 4400 1010
rect 4366 908 4400 942
rect 4366 840 4400 874
rect 4366 772 4400 806
rect 4366 704 4400 738
rect 4366 636 4400 670
rect 4366 568 4400 602
rect 4366 500 4400 534
rect 4366 432 4400 466
rect 4366 364 4400 398
rect 4366 296 4400 330
rect 4366 228 4400 262
rect 4366 160 4400 194
rect 4472 1044 4506 1078
rect 4472 976 4506 1010
rect 4472 908 4506 942
rect 4472 840 4506 874
rect 4472 772 4506 806
rect 4472 704 4506 738
rect 4472 636 4506 670
rect 4472 568 4506 602
rect 4472 500 4506 534
rect 4472 432 4506 466
rect 4472 364 4506 398
rect 4472 296 4506 330
rect 4472 228 4506 262
rect 4472 160 4506 194
rect 4578 1044 4612 1078
rect 4578 976 4612 1010
rect 4578 908 4612 942
rect 4578 840 4612 874
rect 4578 772 4612 806
rect 4578 704 4612 738
rect 4578 636 4612 670
rect 4578 568 4612 602
rect 4578 500 4612 534
rect 4578 432 4612 466
rect 4578 364 4612 398
rect 4578 296 4612 330
rect 4578 228 4612 262
rect 4578 160 4612 194
rect 4684 1044 4718 1078
rect 4684 976 4718 1010
rect 4684 908 4718 942
rect 4684 840 4718 874
rect 4684 772 4718 806
rect 4684 704 4718 738
rect 4684 636 4718 670
rect 4684 568 4718 602
rect 4684 500 4718 534
rect 4684 432 4718 466
rect 4684 364 4718 398
rect 4684 296 4718 330
rect 4684 228 4718 262
rect 4684 160 4718 194
rect 4790 1044 4824 1078
rect 4790 976 4824 1010
rect 4790 908 4824 942
rect 4790 840 4824 874
rect 4790 772 4824 806
rect 4790 704 4824 738
rect 4790 636 4824 670
rect 4790 568 4824 602
rect 4790 500 4824 534
rect 4790 432 4824 466
rect 4790 364 4824 398
rect 4790 296 4824 330
rect 4790 228 4824 262
rect 4790 160 4824 194
rect 4896 1044 4930 1078
rect 4896 976 4930 1010
rect 4896 908 4930 942
rect 4896 840 4930 874
rect 4896 772 4930 806
rect 4896 704 4930 738
rect 4896 636 4930 670
rect 4896 568 4930 602
rect 4896 500 4930 534
rect 4896 432 4930 466
rect 4896 364 4930 398
rect 4896 296 4930 330
rect 4896 228 4930 262
rect 4896 160 4930 194
rect 5002 1044 5036 1078
rect 5002 976 5036 1010
rect 5002 908 5036 942
rect 5002 840 5036 874
rect 5002 772 5036 806
rect 5002 704 5036 738
rect 5002 636 5036 670
rect 5002 568 5036 602
rect 5002 500 5036 534
rect 5002 432 5036 466
rect 5002 364 5036 398
rect 5002 296 5036 330
rect 5002 228 5036 262
rect 5002 160 5036 194
rect 5108 1044 5142 1078
rect 5108 976 5142 1010
rect 5108 908 5142 942
rect 5108 840 5142 874
rect 5108 772 5142 806
rect 5108 704 5142 738
rect 5108 636 5142 670
rect 5108 568 5142 602
rect 5108 500 5142 534
rect 5108 432 5142 466
rect 5108 364 5142 398
rect 5108 296 5142 330
rect 5108 228 5142 262
rect 5108 160 5142 194
rect 5214 1044 5248 1078
rect 5214 976 5248 1010
rect 5214 908 5248 942
rect 5214 840 5248 874
rect 5214 772 5248 806
rect 5214 704 5248 738
rect 5214 636 5248 670
rect 5214 568 5248 602
rect 5214 500 5248 534
rect 5214 432 5248 466
rect 5214 364 5248 398
rect 5214 296 5248 330
rect 5214 228 5248 262
rect 5214 160 5248 194
rect 5320 1044 5354 1078
rect 5320 976 5354 1010
rect 5320 908 5354 942
rect 5320 840 5354 874
rect 5320 772 5354 806
rect 5320 704 5354 738
rect 5320 636 5354 670
rect 5320 568 5354 602
rect 5320 500 5354 534
rect 5320 432 5354 466
rect 5320 364 5354 398
rect 5320 296 5354 330
rect 5320 228 5354 262
rect 5320 160 5354 194
rect 5426 1044 5460 1078
rect 5426 976 5460 1010
rect 5426 908 5460 942
rect 5426 840 5460 874
rect 5426 772 5460 806
rect 5426 704 5460 738
rect 5426 636 5460 670
rect 5426 568 5460 602
rect 5426 500 5460 534
rect 5426 432 5460 466
rect 5426 364 5460 398
rect 5426 296 5460 330
rect 5426 228 5460 262
rect 5426 160 5460 194
rect 5532 1044 5566 1078
rect 5532 976 5566 1010
rect 5532 908 5566 942
rect 5532 840 5566 874
rect 5532 772 5566 806
rect 5532 704 5566 738
rect 5532 636 5566 670
rect 5532 568 5566 602
rect 5532 500 5566 534
rect 5532 432 5566 466
rect 5532 364 5566 398
rect 5532 296 5566 330
rect 5532 228 5566 262
rect 5532 160 5566 194
rect 5638 1044 5672 1078
rect 5638 976 5672 1010
rect 5638 908 5672 942
rect 5638 840 5672 874
rect 5638 772 5672 806
rect 5638 704 5672 738
rect 5638 636 5672 670
rect 5638 568 5672 602
rect 5638 500 5672 534
rect 5638 432 5672 466
rect 5638 364 5672 398
rect 5638 296 5672 330
rect 5638 228 5672 262
rect 5638 160 5672 194
<< mvndiffc >>
rect -101 2726 -67 2760
rect -101 2658 -67 2692
rect -101 2590 -67 2624
rect -101 2522 -67 2556
rect -101 2454 -67 2488
rect -101 2386 -67 2420
rect -101 2318 -67 2352
rect -101 2250 -67 2284
rect 55 2726 89 2760
rect 55 2658 89 2692
rect 55 2590 89 2624
rect 55 2522 89 2556
rect 55 2454 89 2488
rect 55 2386 89 2420
rect 55 2318 89 2352
rect 55 2250 89 2284
rect 12268 2626 12302 2660
rect 12336 2626 12370 2660
rect 12404 2626 12438 2660
rect 12472 2626 12506 2660
rect 12540 2626 12574 2660
rect 12608 2626 12642 2660
rect 12676 2626 12710 2660
rect 12744 2626 12778 2660
rect 12812 2626 12846 2660
rect 12880 2626 12914 2660
rect 12948 2626 12982 2660
rect 13016 2626 13050 2660
rect 13084 2626 13118 2660
rect 13152 2626 13186 2660
rect 13220 2626 13254 2660
rect 13288 2626 13322 2660
rect 13356 2626 13390 2660
rect 13424 2626 13458 2660
rect 13492 2626 13526 2660
rect 13560 2626 13594 2660
rect 13628 2626 13662 2660
rect 13696 2626 13730 2660
rect 13764 2626 13798 2660
rect 13832 2626 13866 2660
rect 13900 2626 13934 2660
rect 13968 2626 14002 2660
rect 14036 2626 14070 2660
rect 14104 2626 14138 2660
rect 14172 2626 14206 2660
rect 14912 2626 14946 2660
rect 14980 2626 15014 2660
rect 15048 2626 15082 2660
rect 15116 2626 15150 2660
rect 15184 2626 15218 2660
rect 15252 2626 15286 2660
rect 15320 2626 15354 2660
rect 15388 2626 15422 2660
rect 15456 2626 15490 2660
rect 15524 2626 15558 2660
rect 15592 2626 15626 2660
rect 15660 2626 15694 2660
rect 15728 2626 15762 2660
rect 15796 2626 15830 2660
rect 15864 2626 15898 2660
rect 15932 2626 15966 2660
rect 16000 2626 16034 2660
rect 16068 2626 16102 2660
rect 16136 2626 16170 2660
rect 16204 2626 16238 2660
rect 16272 2626 16306 2660
rect 16340 2626 16374 2660
rect 16408 2626 16442 2660
rect 16476 2626 16510 2660
rect 16544 2626 16578 2660
rect 16612 2626 16646 2660
rect 16680 2626 16714 2660
rect 16748 2626 16782 2660
rect 16816 2626 16850 2660
rect 12268 2390 12302 2424
rect 12336 2390 12370 2424
rect 12404 2390 12438 2424
rect 12472 2390 12506 2424
rect 12540 2390 12574 2424
rect 12608 2390 12642 2424
rect 12676 2390 12710 2424
rect 12744 2390 12778 2424
rect 12812 2390 12846 2424
rect 12880 2390 12914 2424
rect 12948 2390 12982 2424
rect 13016 2390 13050 2424
rect 13084 2390 13118 2424
rect 13152 2390 13186 2424
rect 13220 2390 13254 2424
rect 13288 2390 13322 2424
rect 13356 2390 13390 2424
rect 13424 2390 13458 2424
rect 13492 2390 13526 2424
rect 13560 2390 13594 2424
rect 13628 2390 13662 2424
rect 13696 2390 13730 2424
rect 13764 2390 13798 2424
rect 13832 2390 13866 2424
rect 13900 2390 13934 2424
rect 13968 2390 14002 2424
rect 14036 2390 14070 2424
rect 14104 2390 14138 2424
rect 14172 2390 14206 2424
rect 12268 2154 12302 2188
rect 12336 2154 12370 2188
rect 12404 2154 12438 2188
rect 12472 2154 12506 2188
rect 12540 2154 12574 2188
rect 12608 2154 12642 2188
rect 12676 2154 12710 2188
rect 12744 2154 12778 2188
rect 12812 2154 12846 2188
rect 12880 2154 12914 2188
rect 12948 2154 12982 2188
rect 13016 2154 13050 2188
rect 13084 2154 13118 2188
rect 13152 2154 13186 2188
rect 13220 2154 13254 2188
rect 13288 2154 13322 2188
rect 13356 2154 13390 2188
rect 13424 2154 13458 2188
rect 13492 2154 13526 2188
rect 13560 2154 13594 2188
rect 13628 2154 13662 2188
rect 13696 2154 13730 2188
rect 13764 2154 13798 2188
rect 13832 2154 13866 2188
rect 13900 2154 13934 2188
rect 13968 2154 14002 2188
rect 14036 2154 14070 2188
rect 14104 2154 14138 2188
rect 14172 2154 14206 2188
rect 12268 1918 12302 1952
rect 12336 1918 12370 1952
rect 12404 1918 12438 1952
rect 12472 1918 12506 1952
rect 12540 1918 12574 1952
rect 12608 1918 12642 1952
rect 12676 1918 12710 1952
rect 12744 1918 12778 1952
rect 12812 1918 12846 1952
rect 12880 1918 12914 1952
rect 12948 1918 12982 1952
rect 13016 1918 13050 1952
rect 13084 1918 13118 1952
rect 13152 1918 13186 1952
rect 13220 1918 13254 1952
rect 13288 1918 13322 1952
rect 13356 1918 13390 1952
rect 13424 1918 13458 1952
rect 13492 1918 13526 1952
rect 13560 1918 13594 1952
rect 13628 1918 13662 1952
rect 13696 1918 13730 1952
rect 13764 1918 13798 1952
rect 13832 1918 13866 1952
rect 13900 1918 13934 1952
rect 13968 1918 14002 1952
rect 14036 1918 14070 1952
rect 14104 1918 14138 1952
rect 14172 1918 14206 1952
rect 14912 2390 14946 2424
rect 14980 2390 15014 2424
rect 15048 2390 15082 2424
rect 15116 2390 15150 2424
rect 15184 2390 15218 2424
rect 15252 2390 15286 2424
rect 15320 2390 15354 2424
rect 15388 2390 15422 2424
rect 15456 2390 15490 2424
rect 15524 2390 15558 2424
rect 15592 2390 15626 2424
rect 15660 2390 15694 2424
rect 15728 2390 15762 2424
rect 15796 2390 15830 2424
rect 15864 2390 15898 2424
rect 15932 2390 15966 2424
rect 16000 2390 16034 2424
rect 16068 2390 16102 2424
rect 16136 2390 16170 2424
rect 16204 2390 16238 2424
rect 16272 2390 16306 2424
rect 16340 2390 16374 2424
rect 16408 2390 16442 2424
rect 16476 2390 16510 2424
rect 16544 2390 16578 2424
rect 16612 2390 16646 2424
rect 16680 2390 16714 2424
rect 16748 2390 16782 2424
rect 16816 2390 16850 2424
rect 14912 2154 14946 2188
rect 14980 2154 15014 2188
rect 15048 2154 15082 2188
rect 15116 2154 15150 2188
rect 15184 2154 15218 2188
rect 15252 2154 15286 2188
rect 15320 2154 15354 2188
rect 15388 2154 15422 2188
rect 15456 2154 15490 2188
rect 15524 2154 15558 2188
rect 15592 2154 15626 2188
rect 15660 2154 15694 2188
rect 15728 2154 15762 2188
rect 15796 2154 15830 2188
rect 15864 2154 15898 2188
rect 15932 2154 15966 2188
rect 16000 2154 16034 2188
rect 16068 2154 16102 2188
rect 16136 2154 16170 2188
rect 16204 2154 16238 2188
rect 16272 2154 16306 2188
rect 16340 2154 16374 2188
rect 16408 2154 16442 2188
rect 16476 2154 16510 2188
rect 16544 2154 16578 2188
rect 16612 2154 16646 2188
rect 16680 2154 16714 2188
rect 16748 2154 16782 2188
rect 16816 2154 16850 2188
rect 14912 1918 14946 1952
rect 14980 1918 15014 1952
rect 15048 1918 15082 1952
rect 15116 1918 15150 1952
rect 15184 1918 15218 1952
rect 15252 1918 15286 1952
rect 15320 1918 15354 1952
rect 15388 1918 15422 1952
rect 15456 1918 15490 1952
rect 15524 1918 15558 1952
rect 15592 1918 15626 1952
rect 15660 1918 15694 1952
rect 15728 1918 15762 1952
rect 15796 1918 15830 1952
rect 15864 1918 15898 1952
rect 15932 1918 15966 1952
rect 16000 1918 16034 1952
rect 16068 1918 16102 1952
rect 16136 1918 16170 1952
rect 16204 1918 16238 1952
rect 16272 1918 16306 1952
rect 16340 1918 16374 1952
rect 16408 1918 16442 1952
rect 16476 1918 16510 1952
rect 16544 1918 16578 1952
rect 16612 1918 16646 1952
rect 16680 1918 16714 1952
rect 16748 1918 16782 1952
rect 16816 1918 16850 1952
rect 5900 1096 5934 1130
rect 5900 1028 5934 1062
rect 5900 960 5934 994
rect 6116 1096 6150 1130
rect 6116 1028 6150 1062
rect 6116 960 6150 994
rect 6332 1096 6366 1130
rect 6332 1028 6366 1062
rect 6332 960 6366 994
rect 6548 1096 6582 1130
rect 6548 1028 6582 1062
rect 6548 960 6582 994
rect 6658 1036 6692 1070
rect 6658 968 6692 1002
rect 6658 900 6692 934
rect 6658 832 6692 866
rect 5900 766 5934 800
rect 5900 698 5934 732
rect 5900 630 5934 664
rect 6116 766 6150 800
rect 6116 698 6150 732
rect 6116 630 6150 664
rect 6332 766 6366 800
rect 6332 698 6366 732
rect 6332 630 6366 664
rect 6548 766 6582 800
rect 6548 698 6582 732
rect 6548 630 6582 664
rect 6658 764 6692 798
rect 6658 696 6692 730
rect 6658 628 6692 662
rect 6658 560 6692 594
rect 6814 1036 6848 1070
rect 6814 968 6848 1002
rect 6814 900 6848 934
rect 6814 832 6848 866
rect 6814 764 6848 798
rect 6814 696 6848 730
rect 6814 628 6848 662
rect 6814 560 6848 594
rect 6970 1036 7004 1070
rect 6970 968 7004 1002
rect 6970 900 7004 934
rect 6970 832 7004 866
rect 6970 764 7004 798
rect 6970 696 7004 730
rect 6970 628 7004 662
rect 6970 560 7004 594
rect 7126 1036 7160 1070
rect 7126 968 7160 1002
rect 7126 900 7160 934
rect 7126 832 7160 866
rect 7126 764 7160 798
rect 7126 696 7160 730
rect 7126 628 7160 662
rect 7126 560 7160 594
rect 7236 1044 7270 1078
rect 7236 976 7270 1010
rect 7236 908 7270 942
rect 7236 840 7270 874
rect 7236 772 7270 806
rect 7236 704 7270 738
rect 7236 636 7270 670
rect 7236 568 7270 602
rect 7236 500 7270 534
rect 5900 400 5934 434
rect 5900 332 5934 366
rect 5900 264 5934 298
rect 6116 400 6150 434
rect 6116 332 6150 366
rect 6116 264 6150 298
rect 6332 400 6366 434
rect 6332 332 6366 366
rect 6332 264 6366 298
rect 6548 400 6582 434
rect 6548 332 6582 366
rect 6548 264 6582 298
rect 7236 432 7270 466
rect 7236 364 7270 398
rect 7236 296 7270 330
rect 7236 228 7270 262
rect 7236 160 7270 194
rect 7392 1044 7426 1078
rect 7392 976 7426 1010
rect 7392 908 7426 942
rect 7392 840 7426 874
rect 7392 772 7426 806
rect 7392 704 7426 738
rect 7392 636 7426 670
rect 7392 568 7426 602
rect 7392 500 7426 534
rect 7392 432 7426 466
rect 7392 364 7426 398
rect 7392 296 7426 330
rect 7392 228 7426 262
rect 7392 160 7426 194
rect 7502 1044 7536 1078
rect 7502 976 7536 1010
rect 7502 908 7536 942
rect 7502 840 7536 874
rect 7502 772 7536 806
rect 7502 704 7536 738
rect 7502 636 7536 670
rect 7502 568 7536 602
rect 7502 500 7536 534
rect 7502 432 7536 466
rect 7502 364 7536 398
rect 7502 296 7536 330
rect 7502 228 7536 262
rect 7502 160 7536 194
rect 7718 1044 7752 1078
rect 7718 976 7752 1010
rect 7718 908 7752 942
rect 7718 840 7752 874
rect 7718 772 7752 806
rect 7718 704 7752 738
rect 7718 636 7752 670
rect 7718 568 7752 602
rect 7718 500 7752 534
rect 7718 432 7752 466
rect 7718 364 7752 398
rect 7718 296 7752 330
rect 7718 228 7752 262
rect 7718 160 7752 194
rect 7934 1044 7968 1078
rect 7934 976 7968 1010
rect 7934 908 7968 942
rect 7934 840 7968 874
rect 7934 772 7968 806
rect 7934 704 7968 738
rect 7934 636 7968 670
rect 7934 568 7968 602
rect 7934 500 7968 534
rect 7934 432 7968 466
rect 7934 364 7968 398
rect 7934 296 7968 330
rect 7934 228 7968 262
rect 7934 160 7968 194
rect 8150 1044 8184 1078
rect 8150 976 8184 1010
rect 8150 908 8184 942
rect 8150 840 8184 874
rect 8150 772 8184 806
rect 8150 704 8184 738
rect 8150 636 8184 670
rect 8150 568 8184 602
rect 8150 500 8184 534
rect 8150 432 8184 466
rect 8150 364 8184 398
rect 8150 296 8184 330
rect 8150 228 8184 262
rect 8150 160 8184 194
rect 8366 1044 8400 1078
rect 8366 976 8400 1010
rect 8366 908 8400 942
rect 8366 840 8400 874
rect 8366 772 8400 806
rect 8366 704 8400 738
rect 8366 636 8400 670
rect 8366 568 8400 602
rect 8366 500 8400 534
rect 8366 432 8400 466
rect 8366 364 8400 398
rect 8366 296 8400 330
rect 8366 228 8400 262
rect 8366 160 8400 194
rect 8582 1044 8616 1078
rect 8582 976 8616 1010
rect 8582 908 8616 942
rect 8582 840 8616 874
rect 8582 772 8616 806
rect 8582 704 8616 738
rect 8582 636 8616 670
rect 8582 568 8616 602
rect 8582 500 8616 534
rect 8582 432 8616 466
rect 8582 364 8616 398
rect 8582 296 8616 330
rect 8582 228 8616 262
rect 8582 160 8616 194
rect 8798 1044 8832 1078
rect 8798 976 8832 1010
rect 8798 908 8832 942
rect 8798 840 8832 874
rect 8798 772 8832 806
rect 8798 704 8832 738
rect 8798 636 8832 670
rect 8798 568 8832 602
rect 8798 500 8832 534
rect 8798 432 8832 466
rect 8798 364 8832 398
rect 8798 296 8832 330
rect 8798 228 8832 262
rect 8798 160 8832 194
rect 9014 1044 9048 1078
rect 9014 976 9048 1010
rect 9014 908 9048 942
rect 9014 840 9048 874
rect 9014 772 9048 806
rect 9014 704 9048 738
rect 9014 636 9048 670
rect 9014 568 9048 602
rect 9014 500 9048 534
rect 9014 432 9048 466
rect 9014 364 9048 398
rect 9014 296 9048 330
rect 9014 228 9048 262
rect 9014 160 9048 194
rect 9230 1044 9264 1078
rect 9230 976 9264 1010
rect 9230 908 9264 942
rect 9230 840 9264 874
rect 9230 772 9264 806
rect 9230 704 9264 738
rect 9230 636 9264 670
rect 9230 568 9264 602
rect 9230 500 9264 534
rect 9230 432 9264 466
rect 9230 364 9264 398
rect 9230 296 9264 330
rect 9230 228 9264 262
rect 9230 160 9264 194
rect 9446 1044 9480 1078
rect 9446 976 9480 1010
rect 9446 908 9480 942
rect 9446 840 9480 874
rect 9446 772 9480 806
rect 9446 704 9480 738
rect 9446 636 9480 670
rect 9446 568 9480 602
rect 9446 500 9480 534
rect 9446 432 9480 466
rect 9446 364 9480 398
rect 9446 296 9480 330
rect 9446 228 9480 262
rect 9446 160 9480 194
rect 9662 1044 9696 1078
rect 9662 976 9696 1010
rect 9662 908 9696 942
rect 9662 840 9696 874
rect 9662 772 9696 806
rect 9662 704 9696 738
rect 9662 636 9696 670
rect 9662 568 9696 602
rect 9662 500 9696 534
rect 9662 432 9696 466
rect 9662 364 9696 398
rect 9662 296 9696 330
rect 9662 228 9696 262
rect 9662 160 9696 194
rect 9878 1044 9912 1078
rect 9878 976 9912 1010
rect 9878 908 9912 942
rect 9878 840 9912 874
rect 9878 772 9912 806
rect 9878 704 9912 738
rect 9878 636 9912 670
rect 9878 568 9912 602
rect 9878 500 9912 534
rect 9878 432 9912 466
rect 9878 364 9912 398
rect 9878 296 9912 330
rect 9878 228 9912 262
rect 9878 160 9912 194
rect 10094 1044 10128 1078
rect 10094 976 10128 1010
rect 10094 908 10128 942
rect 10094 840 10128 874
rect 10094 772 10128 806
rect 10094 704 10128 738
rect 10094 636 10128 670
rect 10094 568 10128 602
rect 10094 500 10128 534
rect 10094 432 10128 466
rect 10094 364 10128 398
rect 10094 296 10128 330
rect 10094 228 10128 262
rect 10094 160 10128 194
rect 10310 1044 10344 1078
rect 10310 976 10344 1010
rect 10310 908 10344 942
rect 10310 840 10344 874
rect 10310 772 10344 806
rect 10310 704 10344 738
rect 10310 636 10344 670
rect 10310 568 10344 602
rect 10310 500 10344 534
rect 10310 432 10344 466
rect 10310 364 10344 398
rect 10310 296 10344 330
rect 10310 228 10344 262
rect 10310 160 10344 194
rect 10526 1044 10560 1078
rect 10526 976 10560 1010
rect 10526 908 10560 942
rect 10526 840 10560 874
rect 10526 772 10560 806
rect 10526 704 10560 738
rect 10526 636 10560 670
rect 10526 568 10560 602
rect 10526 500 10560 534
rect 10526 432 10560 466
rect 10526 364 10560 398
rect 10526 296 10560 330
rect 10526 228 10560 262
rect 10526 160 10560 194
rect 10742 1044 10776 1078
rect 10742 976 10776 1010
rect 10742 908 10776 942
rect 10742 840 10776 874
rect 10742 772 10776 806
rect 10742 704 10776 738
rect 10742 636 10776 670
rect 10742 568 10776 602
rect 10742 500 10776 534
rect 10742 432 10776 466
rect 10742 364 10776 398
rect 10742 296 10776 330
rect 10742 228 10776 262
rect 10742 160 10776 194
rect 10958 1044 10992 1078
rect 10958 976 10992 1010
rect 10958 908 10992 942
rect 10958 840 10992 874
rect 10958 772 10992 806
rect 10958 704 10992 738
rect 10958 636 10992 670
rect 10958 568 10992 602
rect 10958 500 10992 534
rect 10958 432 10992 466
rect 10958 364 10992 398
rect 10958 296 10992 330
rect 10958 228 10992 262
rect 10958 160 10992 194
rect 11174 1044 11208 1078
rect 11174 976 11208 1010
rect 11174 908 11208 942
rect 11174 840 11208 874
rect 11174 772 11208 806
rect 11174 704 11208 738
rect 11174 636 11208 670
rect 11174 568 11208 602
rect 11174 500 11208 534
rect 11174 432 11208 466
rect 11174 364 11208 398
rect 11174 296 11208 330
rect 11174 228 11208 262
rect 11174 160 11208 194
rect 11390 1044 11424 1078
rect 11390 976 11424 1010
rect 11390 908 11424 942
rect 11390 840 11424 874
rect 11390 772 11424 806
rect 11390 704 11424 738
rect 11390 636 11424 670
rect 11390 568 11424 602
rect 11390 500 11424 534
rect 11390 432 11424 466
rect 11390 364 11424 398
rect 11390 296 11424 330
rect 11390 228 11424 262
rect 11390 160 11424 194
rect 11606 1044 11640 1078
rect 11606 976 11640 1010
rect 11606 908 11640 942
rect 11606 840 11640 874
rect 11606 772 11640 806
rect 11606 704 11640 738
rect 11606 636 11640 670
rect 11606 568 11640 602
rect 11606 500 11640 534
rect 11606 432 11640 466
rect 11606 364 11640 398
rect 11606 296 11640 330
rect 11606 228 11640 262
rect 11606 160 11640 194
rect 11822 1044 11856 1078
rect 11822 976 11856 1010
rect 11822 908 11856 942
rect 11822 840 11856 874
rect 11822 772 11856 806
rect 11822 704 11856 738
rect 11822 636 11856 670
rect 11822 568 11856 602
rect 11822 500 11856 534
rect 11822 432 11856 466
rect 11822 364 11856 398
rect 11822 296 11856 330
rect 11822 228 11856 262
rect 11822 160 11856 194
rect 12038 1044 12072 1078
rect 12038 976 12072 1010
rect 12038 908 12072 942
rect 12038 840 12072 874
rect 12038 772 12072 806
rect 12038 704 12072 738
rect 12038 636 12072 670
rect 12038 568 12072 602
rect 12038 500 12072 534
rect 12038 432 12072 466
rect 12038 364 12072 398
rect 12038 296 12072 330
rect 12038 228 12072 262
rect 12038 160 12072 194
rect 12254 1044 12288 1078
rect 12254 976 12288 1010
rect 12254 908 12288 942
rect 12254 840 12288 874
rect 12254 772 12288 806
rect 12254 704 12288 738
rect 12254 636 12288 670
rect 12254 568 12288 602
rect 12254 500 12288 534
rect 12254 432 12288 466
rect 12254 364 12288 398
rect 12254 296 12288 330
rect 12254 228 12288 262
rect 12254 160 12288 194
rect 12470 1044 12504 1078
rect 12470 976 12504 1010
rect 12470 908 12504 942
rect 12470 840 12504 874
rect 12470 772 12504 806
rect 12470 704 12504 738
rect 12470 636 12504 670
rect 12470 568 12504 602
rect 12470 500 12504 534
rect 12470 432 12504 466
rect 12470 364 12504 398
rect 12470 296 12504 330
rect 12470 228 12504 262
rect 12470 160 12504 194
rect 12686 1044 12720 1078
rect 12686 976 12720 1010
rect 12686 908 12720 942
rect 12686 840 12720 874
rect 12686 772 12720 806
rect 12686 704 12720 738
rect 12686 636 12720 670
rect 12686 568 12720 602
rect 12686 500 12720 534
rect 12686 432 12720 466
rect 12686 364 12720 398
rect 12686 296 12720 330
rect 12686 228 12720 262
rect 12686 160 12720 194
rect 12902 1044 12936 1078
rect 12902 976 12936 1010
rect 12902 908 12936 942
rect 12902 840 12936 874
rect 12902 772 12936 806
rect 12902 704 12936 738
rect 12902 636 12936 670
rect 12902 568 12936 602
rect 12902 500 12936 534
rect 12902 432 12936 466
rect 12902 364 12936 398
rect 12902 296 12936 330
rect 12902 228 12936 262
rect 12902 160 12936 194
rect 13118 1044 13152 1078
rect 13118 976 13152 1010
rect 13118 908 13152 942
rect 13118 840 13152 874
rect 13118 772 13152 806
rect 13118 704 13152 738
rect 13118 636 13152 670
rect 13118 568 13152 602
rect 13118 500 13152 534
rect 13118 432 13152 466
rect 13118 364 13152 398
rect 13118 296 13152 330
rect 13118 228 13152 262
rect 13118 160 13152 194
rect 13334 1044 13368 1078
rect 13334 976 13368 1010
rect 13334 908 13368 942
rect 13334 840 13368 874
rect 13334 772 13368 806
rect 13334 704 13368 738
rect 13334 636 13368 670
rect 13334 568 13368 602
rect 13334 500 13368 534
rect 13334 432 13368 466
rect 13334 364 13368 398
rect 13334 296 13368 330
rect 13334 228 13368 262
rect 13334 160 13368 194
rect 13550 1044 13584 1078
rect 13550 976 13584 1010
rect 13550 908 13584 942
rect 13550 840 13584 874
rect 13550 772 13584 806
rect 13550 704 13584 738
rect 13550 636 13584 670
rect 13550 568 13584 602
rect 13550 500 13584 534
rect 13550 432 13584 466
rect 13550 364 13584 398
rect 13550 296 13584 330
rect 13550 228 13584 262
rect 13550 160 13584 194
rect 13766 1044 13800 1078
rect 13766 976 13800 1010
rect 13766 908 13800 942
rect 13766 840 13800 874
rect 13766 772 13800 806
rect 13766 704 13800 738
rect 13766 636 13800 670
rect 13766 568 13800 602
rect 13766 500 13800 534
rect 13766 432 13800 466
rect 13766 364 13800 398
rect 13766 296 13800 330
rect 13766 228 13800 262
rect 13766 160 13800 194
rect 13982 1044 14016 1078
rect 13982 976 14016 1010
rect 13982 908 14016 942
rect 13982 840 14016 874
rect 13982 772 14016 806
rect 13982 704 14016 738
rect 13982 636 14016 670
rect 13982 568 14016 602
rect 13982 500 14016 534
rect 13982 432 14016 466
rect 13982 364 14016 398
rect 13982 296 14016 330
rect 13982 228 14016 262
rect 13982 160 14016 194
rect 14198 1044 14232 1078
rect 14198 976 14232 1010
rect 14198 908 14232 942
rect 14198 840 14232 874
rect 14198 772 14232 806
rect 14198 704 14232 738
rect 14198 636 14232 670
rect 14198 568 14232 602
rect 14198 500 14232 534
rect 14198 432 14232 466
rect 14198 364 14232 398
rect 14198 296 14232 330
rect 14198 228 14232 262
rect 14198 160 14232 194
rect 14414 1044 14448 1078
rect 14414 976 14448 1010
rect 14414 908 14448 942
rect 14414 840 14448 874
rect 14414 772 14448 806
rect 14414 704 14448 738
rect 14414 636 14448 670
rect 14414 568 14448 602
rect 14414 500 14448 534
rect 14414 432 14448 466
rect 14414 364 14448 398
rect 14414 296 14448 330
rect 14414 228 14448 262
rect 14414 160 14448 194
rect 14630 1044 14664 1078
rect 14630 976 14664 1010
rect 14630 908 14664 942
rect 14630 840 14664 874
rect 14630 772 14664 806
rect 14630 704 14664 738
rect 14630 636 14664 670
rect 14630 568 14664 602
rect 14630 500 14664 534
rect 14630 432 14664 466
rect 14630 364 14664 398
rect 14630 296 14664 330
rect 14630 228 14664 262
rect 14630 160 14664 194
rect 14846 1044 14880 1078
rect 14846 976 14880 1010
rect 14846 908 14880 942
rect 14846 840 14880 874
rect 14846 772 14880 806
rect 14846 704 14880 738
rect 14846 636 14880 670
rect 14846 568 14880 602
rect 14846 500 14880 534
rect 14846 432 14880 466
rect 14846 364 14880 398
rect 14846 296 14880 330
rect 14846 228 14880 262
rect 14846 160 14880 194
rect 15062 1044 15096 1078
rect 15062 976 15096 1010
rect 15062 908 15096 942
rect 15062 840 15096 874
rect 15062 772 15096 806
rect 15062 704 15096 738
rect 15062 636 15096 670
rect 15062 568 15096 602
rect 15172 1036 15206 1070
rect 15172 968 15206 1002
rect 15172 900 15206 934
rect 15172 832 15206 866
rect 15172 764 15206 798
rect 15172 696 15206 730
rect 15172 628 15206 662
rect 15172 560 15206 594
rect 15428 1036 15462 1070
rect 15428 968 15462 1002
rect 15428 900 15462 934
rect 15428 832 15462 866
rect 15428 764 15462 798
rect 15428 696 15462 730
rect 15428 628 15462 662
rect 15428 560 15462 594
rect 15538 1044 15572 1078
rect 15538 976 15572 1010
rect 15538 908 15572 942
rect 15538 840 15572 874
rect 15538 772 15572 806
rect 15538 704 15572 738
rect 15538 636 15572 670
rect 15538 568 15572 602
rect 15062 500 15096 534
rect 15062 432 15096 466
rect 15062 364 15096 398
rect 15062 296 15096 330
rect 15062 228 15096 262
rect 15062 160 15096 194
rect 15538 500 15572 534
rect 15538 432 15572 466
rect 15538 364 15572 398
rect 15538 296 15572 330
rect 15538 228 15572 262
rect 15538 160 15572 194
rect 15754 1044 15788 1078
rect 15754 976 15788 1010
rect 15754 908 15788 942
rect 15754 840 15788 874
rect 15754 772 15788 806
rect 15754 704 15788 738
rect 15754 636 15788 670
rect 15754 568 15788 602
rect 15754 500 15788 534
rect 15754 432 15788 466
rect 15754 364 15788 398
rect 15754 296 15788 330
rect 15754 228 15788 262
rect 15754 160 15788 194
rect 15970 1044 16004 1078
rect 15970 976 16004 1010
rect 15970 908 16004 942
rect 15970 840 16004 874
rect 15970 772 16004 806
rect 15970 704 16004 738
rect 15970 636 16004 670
rect 15970 568 16004 602
rect 15970 500 16004 534
rect 15970 432 16004 466
rect 15970 364 16004 398
rect 15970 296 16004 330
rect 15970 228 16004 262
rect 15970 160 16004 194
<< mvpdiffc >>
rect 720 2817 754 2851
rect 720 2749 754 2783
rect 720 2681 754 2715
rect 720 2613 754 2647
rect 720 2545 754 2579
rect 720 2477 754 2511
rect 720 2409 754 2443
rect 720 2341 754 2375
rect 720 2273 754 2307
rect 720 2205 754 2239
rect 720 2137 754 2171
rect 720 2069 754 2103
rect 720 2001 754 2035
rect 720 1933 754 1967
rect 876 2817 910 2851
rect 876 2749 910 2783
rect 876 2681 910 2715
rect 876 2613 910 2647
rect 876 2545 910 2579
rect 876 2477 910 2511
rect 876 2409 910 2443
rect 876 2341 910 2375
rect 876 2273 910 2307
rect 876 2205 910 2239
rect 876 2137 910 2171
rect 876 2069 910 2103
rect 876 2001 910 2035
rect 876 1933 910 1967
rect 1032 2817 1066 2851
rect 1032 2749 1066 2783
rect 1032 2681 1066 2715
rect 1032 2613 1066 2647
rect 1032 2545 1066 2579
rect 1032 2477 1066 2511
rect 1032 2409 1066 2443
rect 1032 2341 1066 2375
rect 1032 2273 1066 2307
rect 1032 2205 1066 2239
rect 1032 2137 1066 2171
rect 1032 2069 1066 2103
rect 1032 2001 1066 2035
rect 1032 1933 1066 1967
rect 1142 2817 1176 2851
rect 1142 2749 1176 2783
rect 1142 2681 1176 2715
rect 1142 2613 1176 2647
rect 1142 2545 1176 2579
rect 1142 2477 1176 2511
rect 1142 2409 1176 2443
rect 1142 2341 1176 2375
rect 1142 2273 1176 2307
rect 1142 2205 1176 2239
rect 1142 2137 1176 2171
rect 1142 2069 1176 2103
rect 1142 2001 1176 2035
rect 1142 1933 1176 1967
rect 1298 2817 1332 2851
rect 1298 2749 1332 2783
rect 1298 2681 1332 2715
rect 1298 2613 1332 2647
rect 1298 2545 1332 2579
rect 1298 2477 1332 2511
rect 1298 2409 1332 2443
rect 1298 2341 1332 2375
rect 1298 2273 1332 2307
rect 1298 2205 1332 2239
rect 1298 2137 1332 2171
rect 1298 2069 1332 2103
rect 1298 2001 1332 2035
rect 1298 1933 1332 1967
rect 1454 2817 1488 2851
rect 1454 2749 1488 2783
rect 1454 2681 1488 2715
rect 1454 2613 1488 2647
rect 1454 2545 1488 2579
rect 1454 2477 1488 2511
rect 1454 2409 1488 2443
rect 1454 2341 1488 2375
rect 1454 2273 1488 2307
rect 1454 2205 1488 2239
rect 1454 2137 1488 2171
rect 1454 2069 1488 2103
rect 1454 2001 1488 2035
rect 1454 1933 1488 1967
rect 1610 2817 1644 2851
rect 1610 2749 1644 2783
rect 1610 2681 1644 2715
rect 1610 2613 1644 2647
rect 1610 2545 1644 2579
rect 1610 2477 1644 2511
rect 1610 2409 1644 2443
rect 1610 2341 1644 2375
rect 1610 2273 1644 2307
rect 1610 2205 1644 2239
rect 1610 2137 1644 2171
rect 1610 2069 1644 2103
rect 1610 2001 1644 2035
rect 1610 1933 1644 1967
rect 1766 2817 1800 2851
rect 1766 2749 1800 2783
rect 1766 2681 1800 2715
rect 1766 2613 1800 2647
rect 1766 2545 1800 2579
rect 1766 2477 1800 2511
rect 1766 2409 1800 2443
rect 1766 2341 1800 2375
rect 1766 2273 1800 2307
rect 1766 2205 1800 2239
rect 1766 2137 1800 2171
rect 1766 2069 1800 2103
rect 1766 2001 1800 2035
rect 1766 1933 1800 1967
rect 1922 2817 1956 2851
rect 1922 2749 1956 2783
rect 1922 2681 1956 2715
rect 1922 2613 1956 2647
rect 1922 2545 1956 2579
rect 1922 2477 1956 2511
rect 1922 2409 1956 2443
rect 1922 2341 1956 2375
rect 1922 2273 1956 2307
rect 1922 2205 1956 2239
rect 1922 2137 1956 2171
rect 1922 2069 1956 2103
rect 1922 2001 1956 2035
rect 1922 1933 1956 1967
rect 2078 2817 2112 2851
rect 2078 2749 2112 2783
rect 2078 2681 2112 2715
rect 2078 2613 2112 2647
rect 2078 2545 2112 2579
rect 2078 2477 2112 2511
rect 2078 2409 2112 2443
rect 2078 2341 2112 2375
rect 2078 2273 2112 2307
rect 2078 2205 2112 2239
rect 2078 2137 2112 2171
rect 2078 2069 2112 2103
rect 2078 2001 2112 2035
rect 2078 1933 2112 1967
rect 2234 2817 2268 2851
rect 2234 2749 2268 2783
rect 2234 2681 2268 2715
rect 2234 2613 2268 2647
rect 2234 2545 2268 2579
rect 2234 2477 2268 2511
rect 2234 2409 2268 2443
rect 2234 2341 2268 2375
rect 2234 2273 2268 2307
rect 2234 2205 2268 2239
rect 2234 2137 2268 2171
rect 2234 2069 2268 2103
rect 2234 2001 2268 2035
rect 2234 1933 2268 1967
rect 2390 2817 2424 2851
rect 2390 2749 2424 2783
rect 2390 2681 2424 2715
rect 2390 2613 2424 2647
rect 2390 2545 2424 2579
rect 2390 2477 2424 2511
rect 2390 2409 2424 2443
rect 2390 2341 2424 2375
rect 2390 2273 2424 2307
rect 2390 2205 2424 2239
rect 2390 2137 2424 2171
rect 2390 2069 2424 2103
rect 2390 2001 2424 2035
rect 2390 1933 2424 1967
rect 2546 2817 2580 2851
rect 2546 2749 2580 2783
rect 2546 2681 2580 2715
rect 2546 2613 2580 2647
rect 2546 2545 2580 2579
rect 2546 2477 2580 2511
rect 2546 2409 2580 2443
rect 2546 2341 2580 2375
rect 2546 2273 2580 2307
rect 2546 2205 2580 2239
rect 2546 2137 2580 2171
rect 2546 2069 2580 2103
rect 2546 2001 2580 2035
rect 2546 1933 2580 1967
rect 2702 2817 2736 2851
rect 2702 2749 2736 2783
rect 2702 2681 2736 2715
rect 2702 2613 2736 2647
rect 2702 2545 2736 2579
rect 2702 2477 2736 2511
rect 2702 2409 2736 2443
rect 2702 2341 2736 2375
rect 2702 2273 2736 2307
rect 2702 2205 2736 2239
rect 2702 2137 2736 2171
rect 2702 2069 2736 2103
rect 2702 2001 2736 2035
rect 2702 1933 2736 1967
rect 2858 2817 2892 2851
rect 2858 2749 2892 2783
rect 2858 2681 2892 2715
rect 2858 2613 2892 2647
rect 2858 2545 2892 2579
rect 2858 2477 2892 2511
rect 2858 2409 2892 2443
rect 2858 2341 2892 2375
rect 2858 2273 2892 2307
rect 2858 2205 2892 2239
rect 2858 2137 2892 2171
rect 2858 2069 2892 2103
rect 2858 2001 2892 2035
rect 2858 1933 2892 1967
rect 3014 2817 3048 2851
rect 3014 2749 3048 2783
rect 3014 2681 3048 2715
rect 3014 2613 3048 2647
rect 3014 2545 3048 2579
rect 3014 2477 3048 2511
rect 3014 2409 3048 2443
rect 3014 2341 3048 2375
rect 3014 2273 3048 2307
rect 3014 2205 3048 2239
rect 3014 2137 3048 2171
rect 3014 2069 3048 2103
rect 3014 2001 3048 2035
rect 3014 1933 3048 1967
rect 3170 2817 3204 2851
rect 3170 2749 3204 2783
rect 3170 2681 3204 2715
rect 3170 2613 3204 2647
rect 3170 2545 3204 2579
rect 3170 2477 3204 2511
rect 3170 2409 3204 2443
rect 3170 2341 3204 2375
rect 3170 2273 3204 2307
rect 3170 2205 3204 2239
rect 3170 2137 3204 2171
rect 3170 2069 3204 2103
rect 3170 2001 3204 2035
rect 3170 1933 3204 1967
rect 3326 2817 3360 2851
rect 3326 2749 3360 2783
rect 3326 2681 3360 2715
rect 3326 2613 3360 2647
rect 3326 2545 3360 2579
rect 3326 2477 3360 2511
rect 3326 2409 3360 2443
rect 3326 2341 3360 2375
rect 3326 2273 3360 2307
rect 3326 2205 3360 2239
rect 3326 2137 3360 2171
rect 3326 2069 3360 2103
rect 3326 2001 3360 2035
rect 3326 1933 3360 1967
rect 3482 2817 3516 2851
rect 3482 2749 3516 2783
rect 3482 2681 3516 2715
rect 3482 2613 3516 2647
rect 3482 2545 3516 2579
rect 3482 2477 3516 2511
rect 3482 2409 3516 2443
rect 3482 2341 3516 2375
rect 3482 2273 3516 2307
rect 3482 2205 3516 2239
rect 3482 2137 3516 2171
rect 3482 2069 3516 2103
rect 3482 2001 3516 2035
rect 3482 1933 3516 1967
rect 3638 2817 3672 2851
rect 3638 2749 3672 2783
rect 3638 2681 3672 2715
rect 3638 2613 3672 2647
rect 3638 2545 3672 2579
rect 3638 2477 3672 2511
rect 3638 2409 3672 2443
rect 3638 2341 3672 2375
rect 3638 2273 3672 2307
rect 3638 2205 3672 2239
rect 3638 2137 3672 2171
rect 3638 2069 3672 2103
rect 3638 2001 3672 2035
rect 3638 1933 3672 1967
rect 3794 2817 3828 2851
rect 3794 2749 3828 2783
rect 3794 2681 3828 2715
rect 3794 2613 3828 2647
rect 3794 2545 3828 2579
rect 3794 2477 3828 2511
rect 3794 2409 3828 2443
rect 3794 2341 3828 2375
rect 3794 2273 3828 2307
rect 3794 2205 3828 2239
rect 3794 2137 3828 2171
rect 3794 2069 3828 2103
rect 3794 2001 3828 2035
rect 3794 1933 3828 1967
rect 3950 2817 3984 2851
rect 3950 2749 3984 2783
rect 3950 2681 3984 2715
rect 3950 2613 3984 2647
rect 3950 2545 3984 2579
rect 3950 2477 3984 2511
rect 3950 2409 3984 2443
rect 3950 2341 3984 2375
rect 3950 2273 3984 2307
rect 3950 2205 3984 2239
rect 3950 2137 3984 2171
rect 3950 2069 3984 2103
rect 3950 2001 3984 2035
rect 3950 1933 3984 1967
rect 4106 2817 4140 2851
rect 4106 2749 4140 2783
rect 4106 2681 4140 2715
rect 4106 2613 4140 2647
rect 4106 2545 4140 2579
rect 4106 2477 4140 2511
rect 4106 2409 4140 2443
rect 4106 2341 4140 2375
rect 4106 2273 4140 2307
rect 4106 2205 4140 2239
rect 4106 2137 4140 2171
rect 4106 2069 4140 2103
rect 4106 2001 4140 2035
rect 4106 1933 4140 1967
rect 4216 2409 4250 2443
rect 4216 2341 4250 2375
rect 4216 2273 4250 2307
rect 4216 2205 4250 2239
rect 4216 2137 4250 2171
rect 4216 2069 4250 2103
rect 4216 2001 4250 2035
rect 4216 1933 4250 1967
rect 4372 2409 4406 2443
rect 4372 2341 4406 2375
rect 4372 2273 4406 2307
rect 4372 2205 4406 2239
rect 4372 2137 4406 2171
rect 4372 2069 4406 2103
rect 4372 2001 4406 2035
rect 4372 1933 4406 1967
rect 4528 2409 4562 2443
rect 4528 2341 4562 2375
rect 4528 2273 4562 2307
rect 4528 2205 4562 2239
rect 4528 2137 4562 2171
rect 4528 2069 4562 2103
rect 4528 2001 4562 2035
rect 4528 1933 4562 1967
rect 5502 2817 5536 2851
rect 5502 2749 5536 2783
rect 5502 2681 5536 2715
rect 5502 2613 5536 2647
rect 5502 2545 5536 2579
rect 5502 2477 5536 2511
rect 5502 2409 5536 2443
rect 5502 2341 5536 2375
rect 5502 2273 5536 2307
rect 5502 2205 5536 2239
rect 5502 2137 5536 2171
rect 5502 2069 5536 2103
rect 5502 2001 5536 2035
rect 5502 1933 5536 1967
rect 5658 2817 5692 2851
rect 5658 2749 5692 2783
rect 5658 2681 5692 2715
rect 5658 2613 5692 2647
rect 5658 2545 5692 2579
rect 5658 2477 5692 2511
rect 5658 2409 5692 2443
rect 5658 2341 5692 2375
rect 5658 2273 5692 2307
rect 5658 2205 5692 2239
rect 5658 2137 5692 2171
rect 5658 2069 5692 2103
rect 5658 2001 5692 2035
rect 5658 1933 5692 1967
rect 5814 2817 5848 2851
rect 5814 2749 5848 2783
rect 5814 2681 5848 2715
rect 5814 2613 5848 2647
rect 5814 2545 5848 2579
rect 5814 2477 5848 2511
rect 5814 2409 5848 2443
rect 5814 2341 5848 2375
rect 5814 2273 5848 2307
rect 5814 2205 5848 2239
rect 5814 2137 5848 2171
rect 5814 2069 5848 2103
rect 5814 2001 5848 2035
rect 5814 1933 5848 1967
rect 6030 2817 6064 2851
rect 6030 2749 6064 2783
rect 6030 2681 6064 2715
rect 6030 2613 6064 2647
rect 6030 2545 6064 2579
rect 6030 2477 6064 2511
rect 6030 2409 6064 2443
rect 6030 2341 6064 2375
rect 6030 2273 6064 2307
rect 6030 2205 6064 2239
rect 6030 2137 6064 2171
rect 6030 2069 6064 2103
rect 6030 2001 6064 2035
rect 6030 1933 6064 1967
rect 6246 2817 6280 2851
rect 6246 2749 6280 2783
rect 6246 2681 6280 2715
rect 6246 2613 6280 2647
rect 6246 2545 6280 2579
rect 6246 2477 6280 2511
rect 6246 2409 6280 2443
rect 6246 2341 6280 2375
rect 6356 2469 6390 2503
rect 6356 2401 6390 2435
rect 6356 2333 6390 2367
rect 6512 2469 6546 2503
rect 6512 2401 6546 2435
rect 6512 2333 6546 2367
rect 6246 2273 6280 2307
rect 6246 2205 6280 2239
rect 6246 2137 6280 2171
rect 6246 2069 6280 2103
rect 6246 2001 6280 2035
rect 6246 1933 6280 1967
rect 7370 2817 7404 2851
rect 7370 2749 7404 2783
rect 7370 2681 7404 2715
rect 7370 2613 7404 2647
rect 7370 2545 7404 2579
rect 7370 2477 7404 2511
rect 7370 2409 7404 2443
rect 7370 2341 7404 2375
rect 7370 2273 7404 2307
rect 7370 2205 7404 2239
rect 7370 2137 7404 2171
rect 7370 2069 7404 2103
rect 7370 2001 7404 2035
rect 7370 1933 7404 1967
rect 7586 2817 7620 2851
rect 7586 2749 7620 2783
rect 7586 2681 7620 2715
rect 7586 2613 7620 2647
rect 7586 2545 7620 2579
rect 7586 2477 7620 2511
rect 7586 2409 7620 2443
rect 7586 2341 7620 2375
rect 7586 2273 7620 2307
rect 7586 2205 7620 2239
rect 7586 2137 7620 2171
rect 7586 2069 7620 2103
rect 7586 2001 7620 2035
rect 7586 1933 7620 1967
rect 7802 2817 7836 2851
rect 7802 2749 7836 2783
rect 7802 2681 7836 2715
rect 7802 2613 7836 2647
rect 7802 2545 7836 2579
rect 7802 2477 7836 2511
rect 7802 2409 7836 2443
rect 7802 2341 7836 2375
rect 7802 2273 7836 2307
rect 7802 2205 7836 2239
rect 7802 2137 7836 2171
rect 7802 2069 7836 2103
rect 7802 2001 7836 2035
rect 7802 1933 7836 1967
rect 8018 2817 8052 2851
rect 8018 2749 8052 2783
rect 8018 2681 8052 2715
rect 8018 2613 8052 2647
rect 8018 2545 8052 2579
rect 8018 2477 8052 2511
rect 8018 2409 8052 2443
rect 8018 2341 8052 2375
rect 8018 2273 8052 2307
rect 8018 2205 8052 2239
rect 8018 2137 8052 2171
rect 8018 2069 8052 2103
rect 8018 2001 8052 2035
rect 8018 1933 8052 1967
rect 8174 2817 8208 2851
rect 8174 2749 8208 2783
rect 8174 2681 8208 2715
rect 8174 2613 8208 2647
rect 8174 2545 8208 2579
rect 8174 2477 8208 2511
rect 8174 2409 8208 2443
rect 8174 2341 8208 2375
rect 8174 2273 8208 2307
rect 8174 2205 8208 2239
rect 8174 2137 8208 2171
rect 8174 2069 8208 2103
rect 8174 2001 8208 2035
rect 8174 1933 8208 1967
rect 8330 2817 8364 2851
rect 8330 2749 8364 2783
rect 8330 2681 8364 2715
rect 8330 2613 8364 2647
rect 8330 2545 8364 2579
rect 8330 2477 8364 2511
rect 8330 2409 8364 2443
rect 8330 2341 8364 2375
rect 8330 2273 8364 2307
rect 8330 2205 8364 2239
rect 8330 2137 8364 2171
rect 8330 2069 8364 2103
rect 8330 2001 8364 2035
rect 8330 1933 8364 1967
rect 8486 2817 8520 2851
rect 8486 2749 8520 2783
rect 8486 2681 8520 2715
rect 8486 2613 8520 2647
rect 8486 2545 8520 2579
rect 8486 2477 8520 2511
rect 8486 2409 8520 2443
rect 8486 2341 8520 2375
rect 8486 2273 8520 2307
rect 8486 2205 8520 2239
rect 8486 2137 8520 2171
rect 8486 2069 8520 2103
rect 8486 2001 8520 2035
rect 8486 1933 8520 1967
rect 8642 2817 8676 2851
rect 8642 2749 8676 2783
rect 8642 2681 8676 2715
rect 8642 2613 8676 2647
rect 8642 2545 8676 2579
rect 8642 2477 8676 2511
rect 8642 2409 8676 2443
rect 8642 2341 8676 2375
rect 8642 2273 8676 2307
rect 8642 2205 8676 2239
rect 8642 2137 8676 2171
rect 8642 2069 8676 2103
rect 8642 2001 8676 2035
rect 8642 1933 8676 1967
rect 9648 2817 9682 2851
rect 9648 2749 9682 2783
rect 9648 2681 9682 2715
rect 9648 2613 9682 2647
rect 9648 2545 9682 2579
rect 9648 2477 9682 2511
rect 9648 2409 9682 2443
rect 9648 2341 9682 2375
rect 9648 2273 9682 2307
rect 9648 2205 9682 2239
rect 9648 2137 9682 2171
rect 9648 2069 9682 2103
rect 9648 2001 9682 2035
rect 9648 1933 9682 1967
rect 9804 2817 9838 2851
rect 9804 2749 9838 2783
rect 9804 2681 9838 2715
rect 9804 2613 9838 2647
rect 9804 2545 9838 2579
rect 9804 2477 9838 2511
rect 9804 2409 9838 2443
rect 9804 2341 9838 2375
rect 9804 2273 9838 2307
rect 9804 2205 9838 2239
rect 9804 2137 9838 2171
rect 9804 2069 9838 2103
rect 9804 2001 9838 2035
rect 9804 1933 9838 1967
rect 9960 2817 9994 2851
rect 9960 2749 9994 2783
rect 9960 2681 9994 2715
rect 9960 2613 9994 2647
rect 9960 2545 9994 2579
rect 9960 2477 9994 2511
rect 9960 2409 9994 2443
rect 9960 2341 9994 2375
rect 9960 2273 9994 2307
rect 9960 2205 9994 2239
rect 9960 2137 9994 2171
rect 9960 2069 9994 2103
rect 9960 2001 9994 2035
rect 9960 1933 9994 1967
rect 10116 2817 10150 2851
rect 10116 2749 10150 2783
rect 10116 2681 10150 2715
rect 10116 2613 10150 2647
rect 10116 2545 10150 2579
rect 10116 2477 10150 2511
rect 10116 2409 10150 2443
rect 10116 2341 10150 2375
rect 10116 2273 10150 2307
rect 10116 2205 10150 2239
rect 10116 2137 10150 2171
rect 10116 2069 10150 2103
rect 10116 2001 10150 2035
rect 10116 1933 10150 1967
rect 10272 2817 10306 2851
rect 10272 2749 10306 2783
rect 10272 2681 10306 2715
rect 10272 2613 10306 2647
rect 10272 2545 10306 2579
rect 10272 2477 10306 2511
rect 10272 2409 10306 2443
rect 10272 2341 10306 2375
rect 10272 2273 10306 2307
rect 10272 2205 10306 2239
rect 10272 2137 10306 2171
rect 10272 2069 10306 2103
rect 10272 2001 10306 2035
rect 10272 1933 10306 1967
rect 10428 2817 10462 2851
rect 10428 2749 10462 2783
rect 10428 2681 10462 2715
rect 10428 2613 10462 2647
rect 10428 2545 10462 2579
rect 10428 2477 10462 2511
rect 10428 2409 10462 2443
rect 10428 2341 10462 2375
rect 10428 2273 10462 2307
rect 10428 2205 10462 2239
rect 10428 2137 10462 2171
rect 10428 2069 10462 2103
rect 10428 2001 10462 2035
rect 10428 1933 10462 1967
rect 10584 2817 10618 2851
rect 10584 2749 10618 2783
rect 10584 2681 10618 2715
rect 10584 2613 10618 2647
rect 10584 2545 10618 2579
rect 10584 2477 10618 2511
rect 10584 2409 10618 2443
rect 10584 2341 10618 2375
rect 10584 2273 10618 2307
rect 10584 2205 10618 2239
rect 10584 2137 10618 2171
rect 10584 2069 10618 2103
rect 10584 2001 10618 2035
rect 10584 1933 10618 1967
rect 10740 2817 10774 2851
rect 10740 2749 10774 2783
rect 10740 2681 10774 2715
rect 10740 2613 10774 2647
rect 10740 2545 10774 2579
rect 10740 2477 10774 2511
rect 10740 2409 10774 2443
rect 10740 2341 10774 2375
rect 10740 2273 10774 2307
rect 10740 2205 10774 2239
rect 10740 2137 10774 2171
rect 10740 2069 10774 2103
rect 10740 2001 10774 2035
rect 10740 1933 10774 1967
rect 10896 2817 10930 2851
rect 10896 2749 10930 2783
rect 10896 2681 10930 2715
rect 10896 2613 10930 2647
rect 10896 2545 10930 2579
rect 10896 2477 10930 2511
rect 10896 2409 10930 2443
rect 10896 2341 10930 2375
rect 10896 2273 10930 2307
rect 10896 2205 10930 2239
rect 10896 2137 10930 2171
rect 10896 2069 10930 2103
rect 10896 2001 10930 2035
rect 10896 1933 10930 1967
rect 11052 2817 11086 2851
rect 11052 2749 11086 2783
rect 11052 2681 11086 2715
rect 11052 2613 11086 2647
rect 11052 2545 11086 2579
rect 11052 2477 11086 2511
rect 11052 2409 11086 2443
rect 11052 2341 11086 2375
rect 11052 2273 11086 2307
rect 11052 2205 11086 2239
rect 11052 2137 11086 2171
rect 11052 2069 11086 2103
rect 11052 2001 11086 2035
rect 11052 1933 11086 1967
rect 11208 2817 11242 2851
rect 11208 2749 11242 2783
rect 11208 2681 11242 2715
rect 11208 2613 11242 2647
rect 11208 2545 11242 2579
rect 11208 2477 11242 2511
rect 11208 2409 11242 2443
rect 11208 2341 11242 2375
rect 11208 2273 11242 2307
rect 11208 2205 11242 2239
rect 11208 2137 11242 2171
rect 11208 2069 11242 2103
rect 11208 2001 11242 2035
rect 11208 1933 11242 1967
rect 11364 2817 11398 2851
rect 11364 2749 11398 2783
rect 11364 2681 11398 2715
rect 11364 2613 11398 2647
rect 11364 2545 11398 2579
rect 11364 2477 11398 2511
rect 11364 2409 11398 2443
rect 11364 2341 11398 2375
rect 11364 2273 11398 2307
rect 11364 2205 11398 2239
rect 11364 2137 11398 2171
rect 11364 2069 11398 2103
rect 11364 2001 11398 2035
rect 11364 1933 11398 1967
rect 11520 2817 11554 2851
rect 11520 2749 11554 2783
rect 11520 2681 11554 2715
rect 11520 2613 11554 2647
rect 11520 2545 11554 2579
rect 11520 2477 11554 2511
rect 11520 2409 11554 2443
rect 11520 2341 11554 2375
rect 11520 2273 11554 2307
rect 11520 2205 11554 2239
rect 11520 2137 11554 2171
rect 11520 2069 11554 2103
rect 11520 2001 11554 2035
rect 11520 1933 11554 1967
<< nsubdiff >>
rect 3934 40 3958 74
rect 3992 40 4028 74
rect 4062 40 4098 74
rect 4132 40 4168 74
rect 4202 40 4238 74
rect 4272 40 4308 74
rect 4342 40 4378 74
rect 4412 40 4448 74
rect 4482 40 4518 74
rect 4552 40 4587 74
rect 4621 40 4656 74
rect 4690 40 4725 74
rect 4759 40 4794 74
rect 4828 40 4863 74
rect 4897 40 4932 74
rect 4966 40 5001 74
rect 5035 40 5070 74
rect 5104 40 5139 74
rect 5173 40 5208 74
rect 5242 40 5277 74
rect 5311 40 5346 74
rect 5380 40 5415 74
rect 5449 40 5484 74
rect 5518 40 5553 74
rect 5587 40 5622 74
rect 5656 40 5680 74
<< mvpsubdiff >>
rect 210 3238 278 3272
rect 312 3238 346 3272
rect 380 3238 414 3272
rect 448 3238 482 3272
rect 516 3238 550 3272
rect 584 3238 618 3272
rect 652 3238 686 3272
rect 720 3238 754 3272
rect 788 3238 822 3272
rect 856 3238 890 3272
rect 924 3238 958 3272
rect 992 3238 1026 3272
rect 1060 3238 1094 3272
rect 1128 3238 1162 3272
rect 1196 3238 1230 3272
rect 1264 3238 1298 3272
rect 1332 3238 1366 3272
rect 1400 3238 1434 3272
rect 1468 3238 1502 3272
rect 1536 3238 1570 3272
rect 1604 3238 1638 3272
rect 1672 3238 1706 3272
rect 1740 3238 1774 3272
rect 1808 3238 1842 3272
rect 1876 3238 1910 3272
rect 1944 3238 1978 3272
rect 2012 3238 2046 3272
rect 2080 3238 2114 3272
rect 2148 3238 2182 3272
rect 2216 3238 2250 3272
rect 2284 3238 2318 3272
rect 2352 3238 2386 3272
rect 2420 3238 2454 3272
rect 2488 3238 2522 3272
rect 2556 3238 2590 3272
rect 2624 3238 2658 3272
rect 2692 3238 2726 3272
rect 2760 3238 2794 3272
rect 2828 3238 2862 3272
rect 2896 3238 2930 3272
rect 2964 3238 2998 3272
rect 3032 3238 3066 3272
rect 3100 3238 3134 3272
rect 3168 3238 3202 3272
rect 3236 3238 3270 3272
rect 3304 3238 3338 3272
rect 3372 3238 3406 3272
rect 3440 3238 3474 3272
rect 3508 3238 3542 3272
rect 3576 3238 3610 3272
rect 3644 3238 3678 3272
rect 3712 3238 3746 3272
rect 3780 3238 3814 3272
rect 3848 3238 3882 3272
rect 3916 3238 3950 3272
rect 3984 3238 4018 3272
rect 4052 3238 4086 3272
rect 4120 3238 4154 3272
rect 4188 3238 4222 3272
rect 4256 3238 4290 3272
rect 4324 3238 4358 3272
rect 4392 3238 4426 3272
rect 4460 3238 4494 3272
rect 4528 3238 4562 3272
rect 4596 3238 4630 3272
rect 4664 3238 4698 3272
rect 4732 3238 4766 3272
rect 4800 3238 4930 3272
rect 210 3191 244 3238
rect 210 3123 244 3157
rect 210 3055 244 3089
rect 4896 3204 4930 3238
rect 4896 3136 4930 3170
rect 4896 3068 4930 3102
rect 210 2987 244 3021
rect 210 2919 244 2953
rect 210 2851 244 2885
rect 210 2783 244 2817
rect 210 2715 244 2749
rect 210 2647 244 2681
rect 210 2579 244 2613
rect 210 2511 244 2545
rect 210 2443 244 2477
rect 210 2375 244 2409
rect 210 2307 244 2341
rect 210 2239 244 2273
rect 210 2171 244 2205
rect 210 2103 244 2137
rect 210 2035 244 2069
rect 210 1967 244 2001
rect 210 1899 244 1933
rect 210 1831 244 1865
rect 210 1763 244 1797
rect 210 1695 244 1729
rect 4896 3000 4930 3034
rect 4896 2932 4930 2966
rect 4896 2864 4930 2898
rect 4896 2796 4930 2830
rect 4896 2728 4930 2762
rect 4896 2660 4930 2694
rect 4896 2592 4930 2626
rect 4896 2524 4930 2558
rect 4896 2456 4930 2490
rect 4896 2388 4930 2422
rect 4896 2320 4930 2354
rect 4896 2252 4930 2286
rect 4896 2184 4930 2218
rect 4896 2116 4930 2150
rect 4896 2048 4930 2082
rect 4896 1980 4930 2014
rect 4896 1912 4930 1946
rect 4896 1844 4930 1878
rect 4896 1776 4930 1810
rect 4896 1708 4930 1742
rect 210 1627 244 1661
rect 210 1559 244 1593
rect 210 1491 244 1525
rect 4896 1640 4930 1674
rect 4896 1491 4930 1606
rect 210 1457 340 1491
rect 374 1457 408 1491
rect 442 1457 476 1491
rect 510 1457 544 1491
rect 578 1457 612 1491
rect 646 1457 680 1491
rect 714 1457 748 1491
rect 782 1457 816 1491
rect 850 1457 884 1491
rect 918 1457 952 1491
rect 986 1457 1020 1491
rect 1054 1457 1088 1491
rect 1122 1457 1156 1491
rect 1190 1457 1224 1491
rect 1258 1457 1292 1491
rect 1326 1457 1360 1491
rect 1394 1457 1428 1491
rect 1462 1457 1496 1491
rect 1530 1457 1564 1491
rect 1598 1457 1632 1491
rect 1666 1457 1700 1491
rect 1734 1457 1768 1491
rect 1802 1457 1836 1491
rect 1870 1457 1904 1491
rect 1938 1457 1972 1491
rect 2006 1457 2040 1491
rect 2074 1457 2108 1491
rect 2142 1457 2176 1491
rect 2210 1457 2244 1491
rect 2278 1457 2312 1491
rect 2346 1457 2380 1491
rect 2414 1457 2448 1491
rect 2482 1457 2516 1491
rect 2550 1457 2584 1491
rect 2618 1457 2652 1491
rect 2686 1457 2720 1491
rect 2754 1457 2788 1491
rect 2822 1457 2856 1491
rect 2890 1457 2924 1491
rect 2958 1457 2992 1491
rect 3026 1457 3060 1491
rect 3094 1457 3128 1491
rect 3162 1457 3196 1491
rect 3230 1457 3264 1491
rect 3298 1457 3332 1491
rect 3366 1457 3400 1491
rect 3434 1457 3468 1491
rect 3502 1457 3536 1491
rect 3570 1457 3604 1491
rect 3638 1457 3672 1491
rect 3706 1457 3740 1491
rect 3774 1457 3808 1491
rect 3842 1457 3876 1491
rect 3910 1457 3944 1491
rect 3978 1457 4012 1491
rect 4046 1457 4080 1491
rect 4114 1457 4148 1491
rect 4182 1457 4216 1491
rect 4250 1457 4284 1491
rect 4318 1457 4352 1491
rect 4386 1457 4420 1491
rect 4454 1457 4488 1491
rect 4522 1457 4556 1491
rect 4590 1457 4624 1491
rect 4658 1457 4692 1491
rect 4726 1457 4760 1491
rect 4794 1457 4828 1491
rect 4862 1457 4930 1491
rect 5099 3238 5177 3272
rect 5211 3238 5245 3272
rect 5279 3238 5313 3272
rect 5347 3238 5381 3272
rect 5415 3238 5449 3272
rect 5483 3238 5517 3272
rect 5551 3238 5585 3272
rect 5619 3238 5653 3272
rect 5687 3238 5721 3272
rect 5755 3238 5789 3272
rect 5823 3238 5857 3272
rect 5891 3238 5925 3272
rect 5959 3238 5993 3272
rect 6027 3238 6061 3272
rect 6095 3238 6129 3272
rect 6163 3238 6197 3272
rect 6231 3238 6265 3272
rect 6299 3238 6333 3272
rect 6367 3238 6401 3272
rect 6435 3238 6469 3272
rect 6503 3238 6537 3272
rect 6571 3238 6605 3272
rect 6639 3238 6673 3272
rect 6707 3238 6741 3272
rect 6775 3238 6809 3272
rect 6843 3238 6911 3272
rect 5099 3204 5133 3238
rect 5099 3136 5133 3170
rect 5099 3068 5133 3102
rect 6877 3191 6911 3238
rect 6877 3123 6911 3157
rect 6877 3055 6911 3089
rect 5099 3000 5133 3034
rect 5099 2932 5133 2966
rect 5099 2864 5133 2898
rect 5099 2796 5133 2830
rect 5099 2728 5133 2762
rect 5099 2660 5133 2694
rect 5099 2592 5133 2626
rect 5099 2524 5133 2558
rect 5099 2456 5133 2490
rect 5099 2388 5133 2422
rect 5099 2320 5133 2354
rect 5099 2252 5133 2286
rect 5099 2184 5133 2218
rect 5099 2116 5133 2150
rect 5099 2048 5133 2082
rect 5099 1980 5133 2014
rect 5099 1912 5133 1946
rect 5099 1844 5133 1878
rect 5099 1776 5133 1810
rect 5099 1708 5133 1742
rect 6877 2987 6911 3021
rect 6877 2919 6911 2953
rect 6877 2851 6911 2885
rect 6877 2783 6911 2817
rect 6877 2715 6911 2749
rect 6877 2647 6911 2681
rect 6877 2579 6911 2613
rect 6877 2511 6911 2545
rect 6877 2443 6911 2477
rect 6877 2375 6911 2409
rect 6877 2307 6911 2341
rect 6877 2239 6911 2273
rect 6877 2171 6911 2205
rect 6877 2103 6911 2137
rect 6877 2035 6911 2069
rect 6877 1967 6911 2001
rect 6877 1899 6911 1933
rect 6877 1831 6911 1865
rect 6877 1763 6911 1797
rect 6877 1695 6911 1729
rect 5099 1640 5133 1674
rect 5099 1491 5133 1606
rect 6877 1627 6911 1661
rect 6877 1559 6911 1593
rect 6877 1491 6911 1525
rect 5099 1457 5167 1491
rect 5201 1457 5235 1491
rect 5269 1457 5303 1491
rect 5337 1457 5371 1491
rect 5405 1457 5439 1491
rect 5473 1457 5507 1491
rect 5541 1457 5575 1491
rect 5609 1457 5643 1491
rect 5677 1457 5711 1491
rect 5745 1457 5779 1491
rect 5813 1457 5847 1491
rect 5881 1457 5915 1491
rect 5949 1457 5983 1491
rect 6017 1457 6051 1491
rect 6085 1457 6119 1491
rect 6153 1457 6187 1491
rect 6221 1457 6255 1491
rect 6289 1457 6323 1491
rect 6357 1457 6391 1491
rect 6425 1457 6459 1491
rect 6493 1457 6527 1491
rect 6561 1457 6595 1491
rect 6629 1457 6663 1491
rect 6697 1457 6731 1491
rect 6765 1457 6799 1491
rect 6833 1457 6911 1491
rect 6999 3238 7114 3272
rect 7148 3238 7182 3272
rect 7216 3238 7250 3272
rect 7284 3238 7318 3272
rect 7352 3238 7386 3272
rect 7420 3238 7454 3272
rect 7488 3238 7522 3272
rect 7556 3238 7590 3272
rect 7624 3238 7658 3272
rect 7692 3238 7726 3272
rect 7760 3238 7794 3272
rect 7828 3238 7862 3272
rect 7896 3238 7930 3272
rect 7964 3238 7998 3272
rect 8032 3238 8066 3272
rect 8100 3238 8134 3272
rect 8168 3238 8202 3272
rect 8236 3238 8270 3272
rect 8304 3238 8338 3272
rect 8372 3238 8406 3272
rect 8440 3238 8474 3272
rect 8508 3238 8542 3272
rect 8576 3238 8610 3272
rect 8644 3238 8678 3272
rect 8712 3238 8746 3272
rect 8780 3238 8814 3272
rect 8848 3238 8882 3272
rect 8916 3238 8950 3272
rect 8984 3238 9052 3272
rect 6999 3204 7033 3238
rect 6999 3136 7033 3170
rect 6999 3068 7033 3102
rect 9018 3191 9052 3238
rect 9018 3123 9052 3157
rect 9018 3055 9052 3089
rect 6999 3000 7033 3034
rect 6999 2932 7033 2966
rect 6999 2864 7033 2898
rect 6999 2796 7033 2830
rect 6999 2728 7033 2762
rect 6999 2660 7033 2694
rect 6999 2592 7033 2626
rect 6999 2524 7033 2558
rect 6999 2456 7033 2490
rect 6999 2388 7033 2422
rect 6999 2320 7033 2354
rect 6999 2252 7033 2286
rect 6999 2184 7033 2218
rect 6999 2116 7033 2150
rect 6999 2048 7033 2082
rect 6999 1980 7033 2014
rect 6999 1912 7033 1946
rect 6999 1844 7033 1878
rect 6999 1776 7033 1810
rect 6999 1708 7033 1742
rect 9018 2987 9052 3021
rect 9018 2919 9052 2953
rect 9018 2851 9052 2885
rect 9018 2783 9052 2817
rect 9018 2715 9052 2749
rect 9018 2647 9052 2681
rect 9018 2579 9052 2613
rect 9018 2511 9052 2545
rect 9018 2443 9052 2477
rect 9018 2375 9052 2409
rect 9018 2307 9052 2341
rect 9018 2239 9052 2273
rect 9018 2171 9052 2205
rect 9018 2103 9052 2137
rect 9018 2035 9052 2069
rect 9018 1967 9052 2001
rect 9018 1899 9052 1933
rect 9018 1831 9052 1865
rect 9018 1763 9052 1797
rect 9018 1695 9052 1729
rect 6999 1640 7033 1674
rect 6999 1491 7033 1606
rect 12208 2744 12232 2778
rect 12266 2744 12302 2778
rect 12336 2744 12372 2778
rect 12406 2744 12442 2778
rect 12476 2744 12512 2778
rect 12546 2744 12582 2778
rect 12616 2744 12651 2778
rect 12685 2744 12720 2778
rect 12754 2744 12789 2778
rect 12823 2744 12858 2778
rect 12892 2744 12927 2778
rect 12961 2744 12996 2778
rect 13030 2744 13065 2778
rect 13099 2744 13134 2778
rect 13168 2744 13203 2778
rect 13237 2744 13272 2778
rect 13306 2744 13341 2778
rect 13375 2744 13410 2778
rect 13444 2744 13479 2778
rect 13513 2744 13548 2778
rect 13582 2744 13617 2778
rect 13651 2744 13686 2778
rect 13720 2744 13755 2778
rect 13789 2744 13824 2778
rect 13858 2744 13893 2778
rect 13927 2744 13962 2778
rect 13996 2744 14031 2778
rect 14065 2744 14100 2778
rect 14134 2744 14169 2778
rect 14203 2744 14227 2778
rect 14853 2744 14877 2778
rect 14911 2744 14947 2778
rect 14981 2744 15017 2778
rect 15051 2744 15087 2778
rect 15121 2744 15157 2778
rect 15191 2744 15227 2778
rect 15261 2744 15296 2778
rect 15330 2744 15365 2778
rect 15399 2744 15434 2778
rect 15468 2744 15503 2778
rect 15537 2744 15572 2778
rect 15606 2744 15641 2778
rect 15675 2744 15710 2778
rect 15744 2744 15779 2778
rect 15813 2744 15848 2778
rect 15882 2744 15917 2778
rect 15951 2744 15986 2778
rect 16020 2744 16055 2778
rect 16089 2744 16124 2778
rect 16158 2744 16193 2778
rect 16227 2744 16262 2778
rect 16296 2744 16331 2778
rect 16365 2744 16400 2778
rect 16434 2744 16469 2778
rect 16503 2744 16538 2778
rect 16572 2744 16607 2778
rect 16641 2744 16676 2778
rect 16710 2744 16745 2778
rect 16779 2744 16814 2778
rect 16848 2744 16872 2778
rect 9018 1627 9052 1661
rect 9018 1559 9052 1593
rect 9018 1491 9052 1525
rect 6999 1457 7067 1491
rect 7101 1457 7135 1491
rect 7169 1457 7203 1491
rect 7237 1457 7271 1491
rect 7305 1457 7339 1491
rect 7373 1457 7407 1491
rect 7441 1457 7475 1491
rect 7509 1457 7543 1491
rect 7577 1457 7611 1491
rect 7645 1457 7679 1491
rect 7713 1457 7747 1491
rect 7781 1457 7815 1491
rect 7849 1457 7883 1491
rect 7917 1457 7951 1491
rect 7985 1457 8019 1491
rect 8053 1457 8087 1491
rect 8121 1457 8155 1491
rect 8189 1457 8223 1491
rect 8257 1457 8291 1491
rect 8325 1457 8359 1491
rect 8393 1457 8427 1491
rect 8461 1457 8495 1491
rect 8529 1457 8563 1491
rect 8597 1457 8631 1491
rect 8665 1457 8699 1491
rect 8733 1457 8767 1491
rect 8801 1457 8835 1491
rect 8869 1457 8903 1491
rect 8937 1457 9052 1491
rect 1499 48 1523 82
rect 1557 48 1597 82
rect 1631 48 1671 82
rect 1705 48 1745 82
rect 1779 48 1819 82
rect 1853 48 1893 82
rect 1927 48 1967 82
rect 2001 48 2040 82
rect 2074 48 2113 82
rect 2147 48 2186 82
rect 2220 48 2259 82
rect 2293 48 2317 82
rect 2979 48 3003 82
rect 3037 48 3072 82
rect 3106 48 3141 82
rect 3175 48 3210 82
rect 3244 48 3279 82
rect 3313 48 3348 82
rect 3382 48 3406 82
rect 5916 40 5940 74
rect 5974 40 6009 74
rect 6043 40 6078 74
rect 6112 40 6147 74
rect 6181 40 6216 74
rect 6250 40 6284 74
rect 6318 40 6352 74
rect 6386 40 6420 74
rect 6454 40 6488 74
rect 6522 40 6556 74
rect 6590 40 6624 74
rect 6658 40 6692 74
rect 6726 40 6760 74
rect 6794 40 6828 74
rect 6862 40 6896 74
rect 6930 40 6964 74
rect 6998 40 7032 74
rect 7066 40 7100 74
rect 7134 40 7168 74
rect 7202 40 7236 74
rect 7270 40 7304 74
rect 7338 40 7372 74
rect 7406 40 7440 74
rect 7474 40 7508 74
rect 7542 40 7576 74
rect 7610 40 7644 74
rect 7678 40 7712 74
rect 7746 40 7780 74
rect 7814 40 7848 74
rect 7882 40 7916 74
rect 7950 40 7984 74
rect 8018 40 8052 74
rect 8086 40 8120 74
rect 8154 40 8188 74
rect 8222 40 8256 74
rect 8290 40 8324 74
rect 8358 40 8392 74
rect 8426 40 8460 74
rect 8494 40 8528 74
rect 8562 40 8596 74
rect 8630 40 8664 74
rect 8698 40 8732 74
rect 8766 40 8800 74
rect 8834 40 8868 74
rect 8902 40 8936 74
rect 8970 40 9004 74
rect 9038 40 9072 74
rect 9106 40 9140 74
rect 9174 40 9208 74
rect 9242 40 9276 74
rect 9310 40 9344 74
rect 9378 40 9412 74
rect 9446 40 9480 74
rect 9514 40 9548 74
rect 9582 40 9616 74
rect 9650 40 9684 74
rect 9718 40 9752 74
rect 9786 40 9820 74
rect 9854 40 9888 74
rect 9922 40 9956 74
rect 9990 40 10024 74
rect 10058 40 10092 74
rect 10126 40 10160 74
rect 10194 40 10228 74
rect 10262 40 10296 74
rect 10330 40 10364 74
rect 10398 40 10432 74
rect 10466 40 10500 74
rect 10534 40 10568 74
rect 10602 40 10636 74
rect 10670 40 10704 74
rect 10738 40 10772 74
rect 10806 40 10840 74
rect 10874 40 10908 74
rect 10942 40 10976 74
rect 11010 40 11044 74
rect 11078 40 11112 74
rect 11146 40 11180 74
rect 11214 40 11248 74
rect 11282 40 11316 74
rect 11350 40 11384 74
rect 11418 40 11452 74
rect 11486 40 11520 74
rect 11554 40 11588 74
rect 11622 40 11656 74
rect 11690 40 11724 74
rect 11758 40 11792 74
rect 11826 40 11860 74
rect 11894 40 11928 74
rect 11962 40 11996 74
rect 12030 40 12064 74
rect 12098 40 12132 74
rect 12166 40 12200 74
rect 12234 40 12268 74
rect 12302 40 12336 74
rect 12370 40 12404 74
rect 12438 40 12472 74
rect 12506 40 12540 74
rect 12574 40 12608 74
rect 12642 40 12676 74
rect 12710 40 12744 74
rect 12778 40 12812 74
rect 12846 40 12880 74
rect 12914 40 12948 74
rect 12982 40 13016 74
rect 13050 40 13084 74
rect 13118 40 13152 74
rect 13186 40 13220 74
rect 13254 40 13288 74
rect 13322 40 13356 74
rect 13390 40 13424 74
rect 13458 40 13492 74
rect 13526 40 13560 74
rect 13594 40 13628 74
rect 13662 40 13696 74
rect 13730 40 13764 74
rect 13798 40 13832 74
rect 13866 40 13900 74
rect 13934 40 13968 74
rect 14002 40 14036 74
rect 14070 40 14104 74
rect 14138 40 14172 74
rect 14206 40 14240 74
rect 14274 40 14308 74
rect 14342 40 14376 74
rect 14410 40 14444 74
rect 14478 40 14512 74
rect 14546 40 14580 74
rect 14614 40 14648 74
rect 14682 40 14716 74
rect 14750 40 14784 74
rect 14818 40 14852 74
rect 14886 40 14920 74
rect 14954 40 14988 74
rect 15022 40 15056 74
rect 15090 40 15124 74
rect 15158 40 15192 74
rect 15226 40 15260 74
rect 15294 40 15328 74
rect 15362 40 15396 74
rect 15430 40 15464 74
rect 15498 40 15532 74
rect 15566 40 15600 74
rect 15634 40 15668 74
rect 15702 40 15736 74
rect 15770 40 15804 74
rect 15838 40 15872 74
rect 15906 40 15940 74
rect 15974 40 15998 74
<< mvnsubdiff >>
rect 433 3015 501 3049
rect 535 3015 569 3049
rect 603 3015 637 3049
rect 671 3015 705 3049
rect 739 3015 773 3049
rect 807 3015 841 3049
rect 875 3015 909 3049
rect 943 3015 977 3049
rect 1011 3015 1045 3049
rect 1079 3015 1113 3049
rect 1147 3015 1181 3049
rect 1215 3015 1249 3049
rect 1283 3015 1317 3049
rect 1351 3015 1385 3049
rect 1419 3015 1453 3049
rect 1487 3015 1521 3049
rect 1555 3015 1589 3049
rect 1623 3015 1657 3049
rect 1691 3015 1725 3049
rect 1759 3015 1793 3049
rect 1827 3015 1861 3049
rect 1895 3015 1929 3049
rect 1963 3015 1997 3049
rect 2031 3015 2065 3049
rect 2099 3015 2133 3049
rect 2167 3015 2201 3049
rect 2235 3015 2269 3049
rect 2303 3015 2337 3049
rect 2371 3015 2405 3049
rect 2439 3015 2473 3049
rect 2507 3015 2541 3049
rect 2575 3015 2609 3049
rect 2643 3015 2677 3049
rect 2711 3015 2745 3049
rect 2779 3015 2813 3049
rect 2847 3015 2881 3049
rect 2915 3015 2949 3049
rect 2983 3015 3017 3049
rect 3051 3015 3085 3049
rect 3119 3015 3153 3049
rect 3187 3015 3221 3049
rect 3255 3015 3289 3049
rect 3323 3015 3357 3049
rect 3391 3015 3425 3049
rect 3459 3015 3493 3049
rect 3527 3015 3561 3049
rect 3595 3015 3629 3049
rect 3663 3015 3697 3049
rect 3731 3015 3765 3049
rect 3799 3015 3833 3049
rect 3867 3015 3901 3049
rect 3935 3015 3969 3049
rect 4003 3015 4037 3049
rect 4071 3015 4105 3049
rect 4139 3015 4173 3049
rect 4207 3015 4241 3049
rect 4275 3015 4309 3049
rect 4343 3015 4377 3049
rect 4411 3015 4445 3049
rect 4479 3015 4513 3049
rect 4547 3015 4581 3049
rect 4615 3015 4707 3049
rect 433 2938 467 3015
rect 4673 2981 4707 3015
rect 433 2870 467 2904
rect 433 2802 467 2836
rect 433 2734 467 2768
rect 433 2666 467 2700
rect 433 2598 467 2632
rect 433 2530 467 2564
rect 433 2462 467 2496
rect 433 2394 467 2428
rect 433 2326 467 2360
rect 433 2258 467 2292
rect 433 2190 467 2224
rect 433 2122 467 2156
rect 433 2054 467 2088
rect 433 1986 467 2020
rect 433 1918 467 1952
rect 4673 2913 4707 2947
rect 4673 2845 4707 2879
rect 4673 2777 4707 2811
rect 4673 2709 4707 2743
rect 4673 2641 4707 2675
rect 4673 2573 4707 2607
rect 4673 2505 4707 2539
rect 4673 2437 4707 2471
rect 4673 2369 4707 2403
rect 4673 2301 4707 2335
rect 4673 2233 4707 2267
rect 4673 2165 4707 2199
rect 4673 2097 4707 2131
rect 4673 2029 4707 2063
rect 4673 1961 4707 1995
rect 433 1850 467 1884
rect 4673 1893 4707 1927
rect 433 1782 467 1816
rect 433 1714 467 1748
rect 4673 1788 4707 1859
rect 4673 1714 4707 1754
rect 433 1680 525 1714
rect 559 1680 593 1714
rect 627 1680 661 1714
rect 695 1680 729 1714
rect 763 1680 797 1714
rect 831 1680 865 1714
rect 899 1680 933 1714
rect 967 1680 1001 1714
rect 1035 1680 1069 1714
rect 1103 1680 1137 1714
rect 1171 1680 1205 1714
rect 1239 1680 1273 1714
rect 1307 1680 1341 1714
rect 1375 1680 1409 1714
rect 1443 1680 1477 1714
rect 1511 1680 1545 1714
rect 1579 1680 1613 1714
rect 1647 1680 1681 1714
rect 1715 1680 1749 1714
rect 1783 1680 1817 1714
rect 1851 1680 1885 1714
rect 1919 1680 1953 1714
rect 1987 1680 2021 1714
rect 2055 1680 2089 1714
rect 2123 1680 2157 1714
rect 2191 1680 2225 1714
rect 2259 1680 2293 1714
rect 2327 1680 2361 1714
rect 2395 1680 2429 1714
rect 2463 1680 2497 1714
rect 2531 1680 2565 1714
rect 2599 1680 2633 1714
rect 2667 1680 2701 1714
rect 2735 1680 2769 1714
rect 2803 1680 2837 1714
rect 2871 1680 2905 1714
rect 2939 1680 2973 1714
rect 3007 1680 3041 1714
rect 3075 1680 3109 1714
rect 3143 1680 3177 1714
rect 3211 1680 3245 1714
rect 3279 1680 3313 1714
rect 3347 1680 3381 1714
rect 3415 1680 3449 1714
rect 3483 1680 3517 1714
rect 3551 1680 3585 1714
rect 3619 1680 3653 1714
rect 3687 1680 3721 1714
rect 3755 1680 3789 1714
rect 3823 1680 3857 1714
rect 3891 1680 3925 1714
rect 3959 1680 3993 1714
rect 4027 1680 4061 1714
rect 4095 1680 4129 1714
rect 4163 1680 4197 1714
rect 4231 1680 4265 1714
rect 4299 1680 4333 1714
rect 4367 1680 4401 1714
rect 4435 1680 4469 1714
rect 4503 1680 4537 1714
rect 4571 1680 4605 1714
rect 4639 1680 4707 1714
rect 5357 3015 5433 3049
rect 5467 3015 5501 3049
rect 5535 3015 5569 3049
rect 5603 3015 5637 3049
rect 5671 3015 5705 3049
rect 5739 3015 5773 3049
rect 5807 3015 5841 3049
rect 5875 3015 5909 3049
rect 5943 3015 5977 3049
rect 6011 3015 6045 3049
rect 6079 3015 6113 3049
rect 6147 3015 6181 3049
rect 6215 3015 6249 3049
rect 6283 3015 6317 3049
rect 6351 3015 6385 3049
rect 6419 3015 6453 3049
rect 6487 3015 6521 3049
rect 6555 3015 6589 3049
rect 6623 3015 6691 3049
rect 5357 2981 5391 3015
rect 5357 2913 5391 2947
rect 6657 2938 6691 3015
rect 5357 2845 5391 2879
rect 5357 2777 5391 2811
rect 5357 2709 5391 2743
rect 5357 2641 5391 2675
rect 5357 2573 5391 2607
rect 5357 2505 5391 2539
rect 5357 2437 5391 2471
rect 5357 2369 5391 2403
rect 5357 2301 5391 2335
rect 5357 2233 5391 2267
rect 5357 2165 5391 2199
rect 5357 2097 5391 2131
rect 5357 2029 5391 2063
rect 5357 1961 5391 1995
rect 5357 1893 5391 1927
rect 6657 2870 6691 2904
rect 6657 2802 6691 2836
rect 6657 2734 6691 2768
rect 6657 2666 6691 2700
rect 6657 2598 6691 2632
rect 6657 2530 6691 2564
rect 6657 2462 6691 2496
rect 6657 2394 6691 2428
rect 6657 2326 6691 2360
rect 6657 2258 6691 2292
rect 6657 2190 6691 2224
rect 6657 2122 6691 2156
rect 6657 2054 6691 2088
rect 6657 1986 6691 2020
rect 5357 1788 5391 1859
rect 6657 1918 6691 1952
rect 6657 1850 6691 1884
rect 5357 1714 5391 1754
rect 6657 1782 6691 1816
rect 6657 1714 6691 1748
rect 5357 1680 5425 1714
rect 5459 1680 5493 1714
rect 5527 1680 5561 1714
rect 5595 1680 5629 1714
rect 5663 1680 5697 1714
rect 5731 1680 5765 1714
rect 5799 1680 5833 1714
rect 5867 1680 5901 1714
rect 5935 1680 5969 1714
rect 6003 1680 6037 1714
rect 6071 1680 6105 1714
rect 6139 1680 6173 1714
rect 6207 1680 6241 1714
rect 6275 1680 6309 1714
rect 6343 1680 6377 1714
rect 6411 1680 6445 1714
rect 6479 1680 6513 1714
rect 6547 1680 6581 1714
rect 6615 1680 6691 1714
rect 7225 3015 7299 3049
rect 7333 3015 7367 3049
rect 7401 3015 7435 3049
rect 7469 3015 7503 3049
rect 7537 3015 7571 3049
rect 7605 3015 7639 3049
rect 7673 3015 7707 3049
rect 7741 3015 7775 3049
rect 7809 3015 7843 3049
rect 7877 3015 7911 3049
rect 7945 3015 7979 3049
rect 8013 3015 8047 3049
rect 8081 3015 8115 3049
rect 8149 3015 8183 3049
rect 8217 3015 8251 3049
rect 8285 3015 8319 3049
rect 8353 3015 8387 3049
rect 8421 3015 8455 3049
rect 8489 3015 8523 3049
rect 8557 3015 8591 3049
rect 8625 3015 8659 3049
rect 8693 3015 8727 3049
rect 8761 3015 8829 3049
rect 7225 2981 7259 3015
rect 7225 2913 7259 2947
rect 8795 2938 8829 3015
rect 7225 2845 7259 2879
rect 7225 2777 7259 2811
rect 7225 2709 7259 2743
rect 7225 2641 7259 2675
rect 7225 2573 7259 2607
rect 7225 2505 7259 2539
rect 7225 2437 7259 2471
rect 7225 2369 7259 2403
rect 7225 2301 7259 2335
rect 7225 2233 7259 2267
rect 7225 2165 7259 2199
rect 7225 2097 7259 2131
rect 7225 2029 7259 2063
rect 7225 1961 7259 1995
rect 7225 1893 7259 1927
rect 8795 2870 8829 2904
rect 8795 2802 8829 2836
rect 8795 2734 8829 2768
rect 8795 2666 8829 2700
rect 8795 2598 8829 2632
rect 8795 2530 8829 2564
rect 8795 2462 8829 2496
rect 8795 2394 8829 2428
rect 8795 2326 8829 2360
rect 8795 2258 8829 2292
rect 8795 2190 8829 2224
rect 8795 2122 8829 2156
rect 8795 2054 8829 2088
rect 8795 1986 8829 2020
rect 7225 1788 7259 1859
rect 8795 1918 8829 1952
rect 8795 1850 8829 1884
rect 7225 1714 7259 1754
rect 8795 1782 8829 1816
rect 8795 1714 8829 1748
rect 7225 1680 7293 1714
rect 7327 1680 7361 1714
rect 7395 1680 7429 1714
rect 7463 1680 7497 1714
rect 7531 1680 7565 1714
rect 7599 1680 7633 1714
rect 7667 1680 7701 1714
rect 7735 1680 7769 1714
rect 7803 1680 7837 1714
rect 7871 1680 7905 1714
rect 7939 1680 7973 1714
rect 8007 1680 8041 1714
rect 8075 1680 8109 1714
rect 8143 1680 8177 1714
rect 8211 1680 8245 1714
rect 8279 1680 8313 1714
rect 8347 1680 8381 1714
rect 8415 1680 8449 1714
rect 8483 1680 8517 1714
rect 8551 1680 8585 1714
rect 8619 1680 8653 1714
rect 8687 1680 8721 1714
rect 8755 1680 8829 1714
rect 9503 3015 9571 3049
rect 9605 3015 9639 3049
rect 9673 3015 9707 3049
rect 9741 3015 9775 3049
rect 9809 3015 9843 3049
rect 9877 3015 9911 3049
rect 9945 3015 9979 3049
rect 10013 3015 10047 3049
rect 10081 3015 10115 3049
rect 10149 3015 10183 3049
rect 10217 3015 10251 3049
rect 10285 3015 10319 3049
rect 10353 3015 10387 3049
rect 10421 3015 10455 3049
rect 10489 3015 10523 3049
rect 10557 3015 10591 3049
rect 10625 3015 10659 3049
rect 10693 3015 10727 3049
rect 10761 3015 10795 3049
rect 10829 3015 10863 3049
rect 10897 3015 10931 3049
rect 10965 3015 10999 3049
rect 11033 3015 11067 3049
rect 11101 3015 11135 3049
rect 11169 3015 11203 3049
rect 11237 3015 11271 3049
rect 11305 3015 11339 3049
rect 11373 3015 11407 3049
rect 11441 3015 11475 3049
rect 11509 3015 11543 3049
rect 11577 3015 11611 3049
rect 11645 3015 11729 3049
rect 9503 2938 9537 3015
rect 11695 2981 11729 3015
rect 9503 2870 9537 2904
rect 9503 2802 9537 2836
rect 9503 2734 9537 2768
rect 9503 2666 9537 2700
rect 9503 2598 9537 2632
rect 9503 2530 9537 2564
rect 9503 2462 9537 2496
rect 9503 2394 9537 2428
rect 9503 2326 9537 2360
rect 9503 2258 9537 2292
rect 9503 2190 9537 2224
rect 9503 2122 9537 2156
rect 9503 2054 9537 2088
rect 9503 1986 9537 2020
rect 9503 1918 9537 1952
rect 11695 2913 11729 2947
rect 11695 2845 11729 2879
rect 11695 2777 11729 2811
rect 11695 2709 11729 2743
rect 11695 2641 11729 2675
rect 11695 2573 11729 2607
rect 11695 2505 11729 2539
rect 11695 2437 11729 2471
rect 11695 2369 11729 2403
rect 11695 2301 11729 2335
rect 11695 2233 11729 2267
rect 11695 2165 11729 2199
rect 11695 2097 11729 2131
rect 11695 2029 11729 2063
rect 9503 1850 9537 1884
rect 11695 1862 11729 1995
rect 9503 1782 9537 1816
rect 9503 1714 9537 1748
rect 11695 1794 11729 1828
rect 11695 1714 11729 1760
rect 9503 1680 9587 1714
rect 9621 1680 9655 1714
rect 9689 1680 9723 1714
rect 9757 1680 9791 1714
rect 9825 1680 9859 1714
rect 9893 1680 9927 1714
rect 9961 1680 9995 1714
rect 10029 1680 10063 1714
rect 10097 1680 10131 1714
rect 10165 1680 10199 1714
rect 10233 1680 10267 1714
rect 10301 1680 10335 1714
rect 10369 1680 10403 1714
rect 10437 1680 10471 1714
rect 10505 1680 10539 1714
rect 10573 1680 10607 1714
rect 10641 1680 10675 1714
rect 10709 1680 10743 1714
rect 10777 1680 10811 1714
rect 10845 1680 10879 1714
rect 10913 1680 10947 1714
rect 10981 1680 11015 1714
rect 11049 1680 11083 1714
rect 11117 1680 11151 1714
rect 11185 1680 11219 1714
rect 11253 1680 11287 1714
rect 11321 1680 11355 1714
rect 11389 1680 11423 1714
rect 11457 1680 11491 1714
rect 11525 1680 11559 1714
rect 11593 1680 11627 1714
rect 11661 1680 11729 1714
rect 11922 3030 12056 3064
rect 12090 3030 12124 3064
rect 12158 3030 12192 3064
rect 12226 3030 12260 3064
rect 12294 3030 12328 3064
rect 12362 3030 12396 3064
rect 12430 3030 12464 3064
rect 12498 3030 12532 3064
rect 12566 3030 12600 3064
rect 12634 3030 12668 3064
rect 12702 3030 12736 3064
rect 12770 3030 12804 3064
rect 12838 3030 12872 3064
rect 12906 3030 12940 3064
rect 12974 3030 13008 3064
rect 13042 3030 13076 3064
rect 13110 3030 13144 3064
rect 13178 3030 13212 3064
rect 13246 3030 13280 3064
rect 13314 3030 13348 3064
rect 13382 3030 13416 3064
rect 13450 3030 13484 3064
rect 13518 3030 13552 3064
rect 13586 3030 13620 3064
rect 13654 3030 13688 3064
rect 13722 3030 13756 3064
rect 13790 3030 13824 3064
rect 13858 3030 13892 3064
rect 13926 3030 13960 3064
rect 13994 3030 14028 3064
rect 14062 3030 14096 3064
rect 14130 3030 14164 3064
rect 14198 3030 14232 3064
rect 14266 3030 14300 3064
rect 14334 3030 14368 3064
rect 14402 3030 14436 3064
rect 14470 3030 14504 3064
rect 14538 3030 14572 3064
rect 14606 3030 14640 3064
rect 14674 3030 14708 3064
rect 14742 3030 14776 3064
rect 14810 3030 14844 3064
rect 14878 3030 14912 3064
rect 14946 3030 14980 3064
rect 15014 3030 15048 3064
rect 15082 3030 15116 3064
rect 15150 3030 15184 3064
rect 15218 3030 15252 3064
rect 15286 3030 15320 3064
rect 15354 3030 15388 3064
rect 15422 3030 15456 3064
rect 15490 3030 15524 3064
rect 15558 3030 15592 3064
rect 15626 3030 15660 3064
rect 15694 3030 15728 3064
rect 15762 3030 15796 3064
rect 15830 3030 15864 3064
rect 15898 3030 15932 3064
rect 15966 3030 16000 3064
rect 16034 3030 16068 3064
rect 16102 3030 16136 3064
rect 16170 3030 16204 3064
rect 16238 3030 16272 3064
rect 16306 3030 16340 3064
rect 16374 3030 16408 3064
rect 16442 3030 16476 3064
rect 16510 3030 16544 3064
rect 16578 3030 16612 3064
rect 16646 3030 16680 3064
rect 16714 3030 16748 3064
rect 16782 3030 16816 3064
rect 16850 3030 16884 3064
rect 16918 3030 16952 3064
rect 16986 3030 17020 3064
rect 17054 3030 17122 3064
rect 11922 2996 11956 3030
rect 11922 2928 11956 2962
rect 11922 2860 11956 2894
rect 11922 2792 11956 2826
rect 14535 2996 14569 3030
rect 14535 2926 14569 2962
rect 14535 2856 14569 2892
rect 14535 2787 14569 2822
rect 11922 2724 11956 2758
rect 17088 2976 17122 3030
rect 17088 2908 17122 2942
rect 17088 2840 17122 2874
rect 11922 2656 11956 2690
rect 14535 2718 14569 2753
rect 17088 2772 17122 2806
rect 11922 2588 11956 2622
rect 14535 2649 14569 2684
rect 17088 2704 17122 2738
rect 17088 2636 17122 2670
rect 11922 2520 11956 2554
rect 11922 2452 11956 2486
rect 11922 2384 11956 2418
rect 11922 2316 11956 2350
rect 11922 2248 11956 2282
rect 11922 2180 11956 2214
rect 11922 2112 11956 2146
rect 11922 2044 11956 2078
rect 11922 1976 11956 2010
rect 14535 2580 14569 2615
rect 14535 2511 14569 2546
rect 14535 2442 14569 2477
rect 14535 2373 14569 2408
rect 14535 2304 14569 2339
rect 14535 2235 14569 2270
rect 14535 2166 14569 2201
rect 14535 2097 14569 2132
rect 14535 2028 14569 2063
rect 11922 1908 11956 1942
rect 14535 1959 14569 1994
rect 17088 2568 17122 2602
rect 17088 2500 17122 2534
rect 17088 2432 17122 2466
rect 17088 2364 17122 2398
rect 17088 2296 17122 2330
rect 17088 2228 17122 2262
rect 17088 2160 17122 2194
rect 17088 2092 17122 2126
rect 17088 2024 17122 2058
rect 11922 1776 11956 1874
rect 11922 1684 11956 1742
rect 14535 1890 14569 1925
rect 17088 1956 17122 1990
rect 14535 1821 14569 1856
rect 14535 1752 14569 1787
rect 14535 1684 14569 1718
rect 17088 1888 17122 1922
rect 17088 1820 17122 1854
rect 17088 1752 17122 1786
rect 17088 1684 17122 1718
rect 11922 1650 11990 1684
rect 12024 1650 12058 1684
rect 12092 1650 12126 1684
rect 12160 1650 12194 1684
rect 12228 1650 12262 1684
rect 12296 1650 12330 1684
rect 12364 1650 12398 1684
rect 12432 1650 12466 1684
rect 12500 1650 12534 1684
rect 12568 1650 12602 1684
rect 12636 1650 12670 1684
rect 12704 1650 12738 1684
rect 12772 1650 12806 1684
rect 12840 1650 12874 1684
rect 12908 1650 12942 1684
rect 12976 1650 13010 1684
rect 13044 1650 13078 1684
rect 13112 1650 13146 1684
rect 13180 1650 13214 1684
rect 13248 1650 13282 1684
rect 13316 1650 13350 1684
rect 13384 1650 13418 1684
rect 13452 1650 13486 1684
rect 13520 1650 13554 1684
rect 13588 1650 13622 1684
rect 13656 1650 13690 1684
rect 13724 1650 13758 1684
rect 13792 1650 13826 1684
rect 13860 1650 13894 1684
rect 13928 1650 13962 1684
rect 13996 1650 14030 1684
rect 14064 1650 14098 1684
rect 14132 1650 14166 1684
rect 14200 1650 14234 1684
rect 14268 1650 14302 1684
rect 14336 1650 14370 1684
rect 14404 1650 14438 1684
rect 14472 1650 14506 1684
rect 14540 1650 14574 1684
rect 14608 1650 14642 1684
rect 14676 1650 14710 1684
rect 14744 1650 14778 1684
rect 14812 1650 14846 1684
rect 14880 1650 14914 1684
rect 14948 1650 14982 1684
rect 15016 1650 15050 1684
rect 15084 1650 15118 1684
rect 15152 1650 15186 1684
rect 15220 1650 15254 1684
rect 15288 1650 15322 1684
rect 15356 1650 15390 1684
rect 15424 1650 15458 1684
rect 15492 1650 15526 1684
rect 15560 1650 15594 1684
rect 15628 1650 15662 1684
rect 15696 1650 15730 1684
rect 15764 1650 15798 1684
rect 15832 1650 15866 1684
rect 15900 1650 15934 1684
rect 15968 1650 16002 1684
rect 16036 1650 16070 1684
rect 16104 1650 16138 1684
rect 16172 1650 16206 1684
rect 16240 1650 16274 1684
rect 16308 1650 16342 1684
rect 16376 1650 16410 1684
rect 16444 1650 16478 1684
rect 16512 1650 16546 1684
rect 16580 1650 16614 1684
rect 16648 1650 16682 1684
rect 16716 1650 16750 1684
rect 16784 1650 16818 1684
rect 16852 1650 16886 1684
rect 16920 1650 16954 1684
rect 16988 1650 17122 1684
rect 1524 1032 1588 1066
rect 1622 1032 1656 1066
rect 1690 1032 1724 1066
rect 1758 1032 1792 1066
rect 1826 1032 1860 1066
rect 1894 1032 1928 1066
rect 1962 1032 1996 1066
rect 2030 1032 2064 1066
rect 2098 1032 2132 1066
rect 2166 1032 2200 1066
rect 2234 1032 2268 1066
rect 2302 1032 2336 1066
rect 2954 1032 3023 1066
rect 3057 1032 3091 1066
rect 3125 1032 3159 1066
rect 3193 1032 3227 1066
rect 3261 1032 3295 1066
rect 3329 1032 3363 1066
rect 3397 1032 3431 1066
<< nsubdiffcont >>
rect 3958 40 3992 74
rect 4028 40 4062 74
rect 4098 40 4132 74
rect 4168 40 4202 74
rect 4238 40 4272 74
rect 4308 40 4342 74
rect 4378 40 4412 74
rect 4448 40 4482 74
rect 4518 40 4552 74
rect 4587 40 4621 74
rect 4656 40 4690 74
rect 4725 40 4759 74
rect 4794 40 4828 74
rect 4863 40 4897 74
rect 4932 40 4966 74
rect 5001 40 5035 74
rect 5070 40 5104 74
rect 5139 40 5173 74
rect 5208 40 5242 74
rect 5277 40 5311 74
rect 5346 40 5380 74
rect 5415 40 5449 74
rect 5484 40 5518 74
rect 5553 40 5587 74
rect 5622 40 5656 74
<< mvpsubdiffcont >>
rect 278 3238 312 3272
rect 346 3238 380 3272
rect 414 3238 448 3272
rect 482 3238 516 3272
rect 550 3238 584 3272
rect 618 3238 652 3272
rect 686 3238 720 3272
rect 754 3238 788 3272
rect 822 3238 856 3272
rect 890 3238 924 3272
rect 958 3238 992 3272
rect 1026 3238 1060 3272
rect 1094 3238 1128 3272
rect 1162 3238 1196 3272
rect 1230 3238 1264 3272
rect 1298 3238 1332 3272
rect 1366 3238 1400 3272
rect 1434 3238 1468 3272
rect 1502 3238 1536 3272
rect 1570 3238 1604 3272
rect 1638 3238 1672 3272
rect 1706 3238 1740 3272
rect 1774 3238 1808 3272
rect 1842 3238 1876 3272
rect 1910 3238 1944 3272
rect 1978 3238 2012 3272
rect 2046 3238 2080 3272
rect 2114 3238 2148 3272
rect 2182 3238 2216 3272
rect 2250 3238 2284 3272
rect 2318 3238 2352 3272
rect 2386 3238 2420 3272
rect 2454 3238 2488 3272
rect 2522 3238 2556 3272
rect 2590 3238 2624 3272
rect 2658 3238 2692 3272
rect 2726 3238 2760 3272
rect 2794 3238 2828 3272
rect 2862 3238 2896 3272
rect 2930 3238 2964 3272
rect 2998 3238 3032 3272
rect 3066 3238 3100 3272
rect 3134 3238 3168 3272
rect 3202 3238 3236 3272
rect 3270 3238 3304 3272
rect 3338 3238 3372 3272
rect 3406 3238 3440 3272
rect 3474 3238 3508 3272
rect 3542 3238 3576 3272
rect 3610 3238 3644 3272
rect 3678 3238 3712 3272
rect 3746 3238 3780 3272
rect 3814 3238 3848 3272
rect 3882 3238 3916 3272
rect 3950 3238 3984 3272
rect 4018 3238 4052 3272
rect 4086 3238 4120 3272
rect 4154 3238 4188 3272
rect 4222 3238 4256 3272
rect 4290 3238 4324 3272
rect 4358 3238 4392 3272
rect 4426 3238 4460 3272
rect 4494 3238 4528 3272
rect 4562 3238 4596 3272
rect 4630 3238 4664 3272
rect 4698 3238 4732 3272
rect 4766 3238 4800 3272
rect 210 3157 244 3191
rect 210 3089 244 3123
rect 210 3021 244 3055
rect 4896 3170 4930 3204
rect 4896 3102 4930 3136
rect 210 2953 244 2987
rect 210 2885 244 2919
rect 210 2817 244 2851
rect 210 2749 244 2783
rect 210 2681 244 2715
rect 210 2613 244 2647
rect 210 2545 244 2579
rect 210 2477 244 2511
rect 210 2409 244 2443
rect 210 2341 244 2375
rect 210 2273 244 2307
rect 210 2205 244 2239
rect 210 2137 244 2171
rect 210 2069 244 2103
rect 210 2001 244 2035
rect 210 1933 244 1967
rect 210 1865 244 1899
rect 210 1797 244 1831
rect 210 1729 244 1763
rect 210 1661 244 1695
rect 4896 3034 4930 3068
rect 4896 2966 4930 3000
rect 4896 2898 4930 2932
rect 4896 2830 4930 2864
rect 4896 2762 4930 2796
rect 4896 2694 4930 2728
rect 4896 2626 4930 2660
rect 4896 2558 4930 2592
rect 4896 2490 4930 2524
rect 4896 2422 4930 2456
rect 4896 2354 4930 2388
rect 4896 2286 4930 2320
rect 4896 2218 4930 2252
rect 4896 2150 4930 2184
rect 4896 2082 4930 2116
rect 4896 2014 4930 2048
rect 4896 1946 4930 1980
rect 4896 1878 4930 1912
rect 4896 1810 4930 1844
rect 4896 1742 4930 1776
rect 210 1593 244 1627
rect 210 1525 244 1559
rect 4896 1674 4930 1708
rect 4896 1606 4930 1640
rect 340 1457 374 1491
rect 408 1457 442 1491
rect 476 1457 510 1491
rect 544 1457 578 1491
rect 612 1457 646 1491
rect 680 1457 714 1491
rect 748 1457 782 1491
rect 816 1457 850 1491
rect 884 1457 918 1491
rect 952 1457 986 1491
rect 1020 1457 1054 1491
rect 1088 1457 1122 1491
rect 1156 1457 1190 1491
rect 1224 1457 1258 1491
rect 1292 1457 1326 1491
rect 1360 1457 1394 1491
rect 1428 1457 1462 1491
rect 1496 1457 1530 1491
rect 1564 1457 1598 1491
rect 1632 1457 1666 1491
rect 1700 1457 1734 1491
rect 1768 1457 1802 1491
rect 1836 1457 1870 1491
rect 1904 1457 1938 1491
rect 1972 1457 2006 1491
rect 2040 1457 2074 1491
rect 2108 1457 2142 1491
rect 2176 1457 2210 1491
rect 2244 1457 2278 1491
rect 2312 1457 2346 1491
rect 2380 1457 2414 1491
rect 2448 1457 2482 1491
rect 2516 1457 2550 1491
rect 2584 1457 2618 1491
rect 2652 1457 2686 1491
rect 2720 1457 2754 1491
rect 2788 1457 2822 1491
rect 2856 1457 2890 1491
rect 2924 1457 2958 1491
rect 2992 1457 3026 1491
rect 3060 1457 3094 1491
rect 3128 1457 3162 1491
rect 3196 1457 3230 1491
rect 3264 1457 3298 1491
rect 3332 1457 3366 1491
rect 3400 1457 3434 1491
rect 3468 1457 3502 1491
rect 3536 1457 3570 1491
rect 3604 1457 3638 1491
rect 3672 1457 3706 1491
rect 3740 1457 3774 1491
rect 3808 1457 3842 1491
rect 3876 1457 3910 1491
rect 3944 1457 3978 1491
rect 4012 1457 4046 1491
rect 4080 1457 4114 1491
rect 4148 1457 4182 1491
rect 4216 1457 4250 1491
rect 4284 1457 4318 1491
rect 4352 1457 4386 1491
rect 4420 1457 4454 1491
rect 4488 1457 4522 1491
rect 4556 1457 4590 1491
rect 4624 1457 4658 1491
rect 4692 1457 4726 1491
rect 4760 1457 4794 1491
rect 4828 1457 4862 1491
rect 5177 3238 5211 3272
rect 5245 3238 5279 3272
rect 5313 3238 5347 3272
rect 5381 3238 5415 3272
rect 5449 3238 5483 3272
rect 5517 3238 5551 3272
rect 5585 3238 5619 3272
rect 5653 3238 5687 3272
rect 5721 3238 5755 3272
rect 5789 3238 5823 3272
rect 5857 3238 5891 3272
rect 5925 3238 5959 3272
rect 5993 3238 6027 3272
rect 6061 3238 6095 3272
rect 6129 3238 6163 3272
rect 6197 3238 6231 3272
rect 6265 3238 6299 3272
rect 6333 3238 6367 3272
rect 6401 3238 6435 3272
rect 6469 3238 6503 3272
rect 6537 3238 6571 3272
rect 6605 3238 6639 3272
rect 6673 3238 6707 3272
rect 6741 3238 6775 3272
rect 6809 3238 6843 3272
rect 5099 3170 5133 3204
rect 5099 3102 5133 3136
rect 5099 3034 5133 3068
rect 6877 3157 6911 3191
rect 6877 3089 6911 3123
rect 5099 2966 5133 3000
rect 5099 2898 5133 2932
rect 5099 2830 5133 2864
rect 5099 2762 5133 2796
rect 5099 2694 5133 2728
rect 5099 2626 5133 2660
rect 5099 2558 5133 2592
rect 5099 2490 5133 2524
rect 5099 2422 5133 2456
rect 5099 2354 5133 2388
rect 5099 2286 5133 2320
rect 5099 2218 5133 2252
rect 5099 2150 5133 2184
rect 5099 2082 5133 2116
rect 5099 2014 5133 2048
rect 5099 1946 5133 1980
rect 5099 1878 5133 1912
rect 5099 1810 5133 1844
rect 5099 1742 5133 1776
rect 5099 1674 5133 1708
rect 6877 3021 6911 3055
rect 6877 2953 6911 2987
rect 6877 2885 6911 2919
rect 6877 2817 6911 2851
rect 6877 2749 6911 2783
rect 6877 2681 6911 2715
rect 6877 2613 6911 2647
rect 6877 2545 6911 2579
rect 6877 2477 6911 2511
rect 6877 2409 6911 2443
rect 6877 2341 6911 2375
rect 6877 2273 6911 2307
rect 6877 2205 6911 2239
rect 6877 2137 6911 2171
rect 6877 2069 6911 2103
rect 6877 2001 6911 2035
rect 6877 1933 6911 1967
rect 6877 1865 6911 1899
rect 6877 1797 6911 1831
rect 6877 1729 6911 1763
rect 5099 1606 5133 1640
rect 6877 1661 6911 1695
rect 6877 1593 6911 1627
rect 6877 1525 6911 1559
rect 5167 1457 5201 1491
rect 5235 1457 5269 1491
rect 5303 1457 5337 1491
rect 5371 1457 5405 1491
rect 5439 1457 5473 1491
rect 5507 1457 5541 1491
rect 5575 1457 5609 1491
rect 5643 1457 5677 1491
rect 5711 1457 5745 1491
rect 5779 1457 5813 1491
rect 5847 1457 5881 1491
rect 5915 1457 5949 1491
rect 5983 1457 6017 1491
rect 6051 1457 6085 1491
rect 6119 1457 6153 1491
rect 6187 1457 6221 1491
rect 6255 1457 6289 1491
rect 6323 1457 6357 1491
rect 6391 1457 6425 1491
rect 6459 1457 6493 1491
rect 6527 1457 6561 1491
rect 6595 1457 6629 1491
rect 6663 1457 6697 1491
rect 6731 1457 6765 1491
rect 6799 1457 6833 1491
rect 7114 3238 7148 3272
rect 7182 3238 7216 3272
rect 7250 3238 7284 3272
rect 7318 3238 7352 3272
rect 7386 3238 7420 3272
rect 7454 3238 7488 3272
rect 7522 3238 7556 3272
rect 7590 3238 7624 3272
rect 7658 3238 7692 3272
rect 7726 3238 7760 3272
rect 7794 3238 7828 3272
rect 7862 3238 7896 3272
rect 7930 3238 7964 3272
rect 7998 3238 8032 3272
rect 8066 3238 8100 3272
rect 8134 3238 8168 3272
rect 8202 3238 8236 3272
rect 8270 3238 8304 3272
rect 8338 3238 8372 3272
rect 8406 3238 8440 3272
rect 8474 3238 8508 3272
rect 8542 3238 8576 3272
rect 8610 3238 8644 3272
rect 8678 3238 8712 3272
rect 8746 3238 8780 3272
rect 8814 3238 8848 3272
rect 8882 3238 8916 3272
rect 8950 3238 8984 3272
rect 6999 3170 7033 3204
rect 6999 3102 7033 3136
rect 6999 3034 7033 3068
rect 9018 3157 9052 3191
rect 9018 3089 9052 3123
rect 6999 2966 7033 3000
rect 6999 2898 7033 2932
rect 6999 2830 7033 2864
rect 6999 2762 7033 2796
rect 6999 2694 7033 2728
rect 6999 2626 7033 2660
rect 6999 2558 7033 2592
rect 6999 2490 7033 2524
rect 6999 2422 7033 2456
rect 6999 2354 7033 2388
rect 6999 2286 7033 2320
rect 6999 2218 7033 2252
rect 6999 2150 7033 2184
rect 6999 2082 7033 2116
rect 6999 2014 7033 2048
rect 6999 1946 7033 1980
rect 6999 1878 7033 1912
rect 6999 1810 7033 1844
rect 6999 1742 7033 1776
rect 6999 1674 7033 1708
rect 9018 3021 9052 3055
rect 9018 2953 9052 2987
rect 9018 2885 9052 2919
rect 9018 2817 9052 2851
rect 9018 2749 9052 2783
rect 9018 2681 9052 2715
rect 9018 2613 9052 2647
rect 9018 2545 9052 2579
rect 9018 2477 9052 2511
rect 9018 2409 9052 2443
rect 9018 2341 9052 2375
rect 9018 2273 9052 2307
rect 9018 2205 9052 2239
rect 9018 2137 9052 2171
rect 9018 2069 9052 2103
rect 9018 2001 9052 2035
rect 9018 1933 9052 1967
rect 9018 1865 9052 1899
rect 9018 1797 9052 1831
rect 9018 1729 9052 1763
rect 6999 1606 7033 1640
rect 9018 1661 9052 1695
rect 12232 2744 12266 2778
rect 12302 2744 12336 2778
rect 12372 2744 12406 2778
rect 12442 2744 12476 2778
rect 12512 2744 12546 2778
rect 12582 2744 12616 2778
rect 12651 2744 12685 2778
rect 12720 2744 12754 2778
rect 12789 2744 12823 2778
rect 12858 2744 12892 2778
rect 12927 2744 12961 2778
rect 12996 2744 13030 2778
rect 13065 2744 13099 2778
rect 13134 2744 13168 2778
rect 13203 2744 13237 2778
rect 13272 2744 13306 2778
rect 13341 2744 13375 2778
rect 13410 2744 13444 2778
rect 13479 2744 13513 2778
rect 13548 2744 13582 2778
rect 13617 2744 13651 2778
rect 13686 2744 13720 2778
rect 13755 2744 13789 2778
rect 13824 2744 13858 2778
rect 13893 2744 13927 2778
rect 13962 2744 13996 2778
rect 14031 2744 14065 2778
rect 14100 2744 14134 2778
rect 14169 2744 14203 2778
rect 14877 2744 14911 2778
rect 14947 2744 14981 2778
rect 15017 2744 15051 2778
rect 15087 2744 15121 2778
rect 15157 2744 15191 2778
rect 15227 2744 15261 2778
rect 15296 2744 15330 2778
rect 15365 2744 15399 2778
rect 15434 2744 15468 2778
rect 15503 2744 15537 2778
rect 15572 2744 15606 2778
rect 15641 2744 15675 2778
rect 15710 2744 15744 2778
rect 15779 2744 15813 2778
rect 15848 2744 15882 2778
rect 15917 2744 15951 2778
rect 15986 2744 16020 2778
rect 16055 2744 16089 2778
rect 16124 2744 16158 2778
rect 16193 2744 16227 2778
rect 16262 2744 16296 2778
rect 16331 2744 16365 2778
rect 16400 2744 16434 2778
rect 16469 2744 16503 2778
rect 16538 2744 16572 2778
rect 16607 2744 16641 2778
rect 16676 2744 16710 2778
rect 16745 2744 16779 2778
rect 16814 2744 16848 2778
rect 9018 1593 9052 1627
rect 9018 1525 9052 1559
rect 7067 1457 7101 1491
rect 7135 1457 7169 1491
rect 7203 1457 7237 1491
rect 7271 1457 7305 1491
rect 7339 1457 7373 1491
rect 7407 1457 7441 1491
rect 7475 1457 7509 1491
rect 7543 1457 7577 1491
rect 7611 1457 7645 1491
rect 7679 1457 7713 1491
rect 7747 1457 7781 1491
rect 7815 1457 7849 1491
rect 7883 1457 7917 1491
rect 7951 1457 7985 1491
rect 8019 1457 8053 1491
rect 8087 1457 8121 1491
rect 8155 1457 8189 1491
rect 8223 1457 8257 1491
rect 8291 1457 8325 1491
rect 8359 1457 8393 1491
rect 8427 1457 8461 1491
rect 8495 1457 8529 1491
rect 8563 1457 8597 1491
rect 8631 1457 8665 1491
rect 8699 1457 8733 1491
rect 8767 1457 8801 1491
rect 8835 1457 8869 1491
rect 8903 1457 8937 1491
rect 1523 48 1557 82
rect 1597 48 1631 82
rect 1671 48 1705 82
rect 1745 48 1779 82
rect 1819 48 1853 82
rect 1893 48 1927 82
rect 1967 48 2001 82
rect 2040 48 2074 82
rect 2113 48 2147 82
rect 2186 48 2220 82
rect 2259 48 2293 82
rect 3003 48 3037 82
rect 3072 48 3106 82
rect 3141 48 3175 82
rect 3210 48 3244 82
rect 3279 48 3313 82
rect 3348 48 3382 82
rect 5940 40 5974 74
rect 6009 40 6043 74
rect 6078 40 6112 74
rect 6147 40 6181 74
rect 6216 40 6250 74
rect 6284 40 6318 74
rect 6352 40 6386 74
rect 6420 40 6454 74
rect 6488 40 6522 74
rect 6556 40 6590 74
rect 6624 40 6658 74
rect 6692 40 6726 74
rect 6760 40 6794 74
rect 6828 40 6862 74
rect 6896 40 6930 74
rect 6964 40 6998 74
rect 7032 40 7066 74
rect 7100 40 7134 74
rect 7168 40 7202 74
rect 7236 40 7270 74
rect 7304 40 7338 74
rect 7372 40 7406 74
rect 7440 40 7474 74
rect 7508 40 7542 74
rect 7576 40 7610 74
rect 7644 40 7678 74
rect 7712 40 7746 74
rect 7780 40 7814 74
rect 7848 40 7882 74
rect 7916 40 7950 74
rect 7984 40 8018 74
rect 8052 40 8086 74
rect 8120 40 8154 74
rect 8188 40 8222 74
rect 8256 40 8290 74
rect 8324 40 8358 74
rect 8392 40 8426 74
rect 8460 40 8494 74
rect 8528 40 8562 74
rect 8596 40 8630 74
rect 8664 40 8698 74
rect 8732 40 8766 74
rect 8800 40 8834 74
rect 8868 40 8902 74
rect 8936 40 8970 74
rect 9004 40 9038 74
rect 9072 40 9106 74
rect 9140 40 9174 74
rect 9208 40 9242 74
rect 9276 40 9310 74
rect 9344 40 9378 74
rect 9412 40 9446 74
rect 9480 40 9514 74
rect 9548 40 9582 74
rect 9616 40 9650 74
rect 9684 40 9718 74
rect 9752 40 9786 74
rect 9820 40 9854 74
rect 9888 40 9922 74
rect 9956 40 9990 74
rect 10024 40 10058 74
rect 10092 40 10126 74
rect 10160 40 10194 74
rect 10228 40 10262 74
rect 10296 40 10330 74
rect 10364 40 10398 74
rect 10432 40 10466 74
rect 10500 40 10534 74
rect 10568 40 10602 74
rect 10636 40 10670 74
rect 10704 40 10738 74
rect 10772 40 10806 74
rect 10840 40 10874 74
rect 10908 40 10942 74
rect 10976 40 11010 74
rect 11044 40 11078 74
rect 11112 40 11146 74
rect 11180 40 11214 74
rect 11248 40 11282 74
rect 11316 40 11350 74
rect 11384 40 11418 74
rect 11452 40 11486 74
rect 11520 40 11554 74
rect 11588 40 11622 74
rect 11656 40 11690 74
rect 11724 40 11758 74
rect 11792 40 11826 74
rect 11860 40 11894 74
rect 11928 40 11962 74
rect 11996 40 12030 74
rect 12064 40 12098 74
rect 12132 40 12166 74
rect 12200 40 12234 74
rect 12268 40 12302 74
rect 12336 40 12370 74
rect 12404 40 12438 74
rect 12472 40 12506 74
rect 12540 40 12574 74
rect 12608 40 12642 74
rect 12676 40 12710 74
rect 12744 40 12778 74
rect 12812 40 12846 74
rect 12880 40 12914 74
rect 12948 40 12982 74
rect 13016 40 13050 74
rect 13084 40 13118 74
rect 13152 40 13186 74
rect 13220 40 13254 74
rect 13288 40 13322 74
rect 13356 40 13390 74
rect 13424 40 13458 74
rect 13492 40 13526 74
rect 13560 40 13594 74
rect 13628 40 13662 74
rect 13696 40 13730 74
rect 13764 40 13798 74
rect 13832 40 13866 74
rect 13900 40 13934 74
rect 13968 40 14002 74
rect 14036 40 14070 74
rect 14104 40 14138 74
rect 14172 40 14206 74
rect 14240 40 14274 74
rect 14308 40 14342 74
rect 14376 40 14410 74
rect 14444 40 14478 74
rect 14512 40 14546 74
rect 14580 40 14614 74
rect 14648 40 14682 74
rect 14716 40 14750 74
rect 14784 40 14818 74
rect 14852 40 14886 74
rect 14920 40 14954 74
rect 14988 40 15022 74
rect 15056 40 15090 74
rect 15124 40 15158 74
rect 15192 40 15226 74
rect 15260 40 15294 74
rect 15328 40 15362 74
rect 15396 40 15430 74
rect 15464 40 15498 74
rect 15532 40 15566 74
rect 15600 40 15634 74
rect 15668 40 15702 74
rect 15736 40 15770 74
rect 15804 40 15838 74
rect 15872 40 15906 74
rect 15940 40 15974 74
<< mvnsubdiffcont >>
rect 501 3015 535 3049
rect 569 3015 603 3049
rect 637 3015 671 3049
rect 705 3015 739 3049
rect 773 3015 807 3049
rect 841 3015 875 3049
rect 909 3015 943 3049
rect 977 3015 1011 3049
rect 1045 3015 1079 3049
rect 1113 3015 1147 3049
rect 1181 3015 1215 3049
rect 1249 3015 1283 3049
rect 1317 3015 1351 3049
rect 1385 3015 1419 3049
rect 1453 3015 1487 3049
rect 1521 3015 1555 3049
rect 1589 3015 1623 3049
rect 1657 3015 1691 3049
rect 1725 3015 1759 3049
rect 1793 3015 1827 3049
rect 1861 3015 1895 3049
rect 1929 3015 1963 3049
rect 1997 3015 2031 3049
rect 2065 3015 2099 3049
rect 2133 3015 2167 3049
rect 2201 3015 2235 3049
rect 2269 3015 2303 3049
rect 2337 3015 2371 3049
rect 2405 3015 2439 3049
rect 2473 3015 2507 3049
rect 2541 3015 2575 3049
rect 2609 3015 2643 3049
rect 2677 3015 2711 3049
rect 2745 3015 2779 3049
rect 2813 3015 2847 3049
rect 2881 3015 2915 3049
rect 2949 3015 2983 3049
rect 3017 3015 3051 3049
rect 3085 3015 3119 3049
rect 3153 3015 3187 3049
rect 3221 3015 3255 3049
rect 3289 3015 3323 3049
rect 3357 3015 3391 3049
rect 3425 3015 3459 3049
rect 3493 3015 3527 3049
rect 3561 3015 3595 3049
rect 3629 3015 3663 3049
rect 3697 3015 3731 3049
rect 3765 3015 3799 3049
rect 3833 3015 3867 3049
rect 3901 3015 3935 3049
rect 3969 3015 4003 3049
rect 4037 3015 4071 3049
rect 4105 3015 4139 3049
rect 4173 3015 4207 3049
rect 4241 3015 4275 3049
rect 4309 3015 4343 3049
rect 4377 3015 4411 3049
rect 4445 3015 4479 3049
rect 4513 3015 4547 3049
rect 4581 3015 4615 3049
rect 433 2904 467 2938
rect 4673 2947 4707 2981
rect 433 2836 467 2870
rect 433 2768 467 2802
rect 433 2700 467 2734
rect 433 2632 467 2666
rect 433 2564 467 2598
rect 433 2496 467 2530
rect 433 2428 467 2462
rect 433 2360 467 2394
rect 433 2292 467 2326
rect 433 2224 467 2258
rect 433 2156 467 2190
rect 433 2088 467 2122
rect 433 2020 467 2054
rect 433 1952 467 1986
rect 4673 2879 4707 2913
rect 4673 2811 4707 2845
rect 4673 2743 4707 2777
rect 4673 2675 4707 2709
rect 4673 2607 4707 2641
rect 4673 2539 4707 2573
rect 4673 2471 4707 2505
rect 4673 2403 4707 2437
rect 4673 2335 4707 2369
rect 4673 2267 4707 2301
rect 4673 2199 4707 2233
rect 4673 2131 4707 2165
rect 4673 2063 4707 2097
rect 4673 1995 4707 2029
rect 4673 1927 4707 1961
rect 433 1884 467 1918
rect 433 1816 467 1850
rect 4673 1859 4707 1893
rect 433 1748 467 1782
rect 4673 1754 4707 1788
rect 525 1680 559 1714
rect 593 1680 627 1714
rect 661 1680 695 1714
rect 729 1680 763 1714
rect 797 1680 831 1714
rect 865 1680 899 1714
rect 933 1680 967 1714
rect 1001 1680 1035 1714
rect 1069 1680 1103 1714
rect 1137 1680 1171 1714
rect 1205 1680 1239 1714
rect 1273 1680 1307 1714
rect 1341 1680 1375 1714
rect 1409 1680 1443 1714
rect 1477 1680 1511 1714
rect 1545 1680 1579 1714
rect 1613 1680 1647 1714
rect 1681 1680 1715 1714
rect 1749 1680 1783 1714
rect 1817 1680 1851 1714
rect 1885 1680 1919 1714
rect 1953 1680 1987 1714
rect 2021 1680 2055 1714
rect 2089 1680 2123 1714
rect 2157 1680 2191 1714
rect 2225 1680 2259 1714
rect 2293 1680 2327 1714
rect 2361 1680 2395 1714
rect 2429 1680 2463 1714
rect 2497 1680 2531 1714
rect 2565 1680 2599 1714
rect 2633 1680 2667 1714
rect 2701 1680 2735 1714
rect 2769 1680 2803 1714
rect 2837 1680 2871 1714
rect 2905 1680 2939 1714
rect 2973 1680 3007 1714
rect 3041 1680 3075 1714
rect 3109 1680 3143 1714
rect 3177 1680 3211 1714
rect 3245 1680 3279 1714
rect 3313 1680 3347 1714
rect 3381 1680 3415 1714
rect 3449 1680 3483 1714
rect 3517 1680 3551 1714
rect 3585 1680 3619 1714
rect 3653 1680 3687 1714
rect 3721 1680 3755 1714
rect 3789 1680 3823 1714
rect 3857 1680 3891 1714
rect 3925 1680 3959 1714
rect 3993 1680 4027 1714
rect 4061 1680 4095 1714
rect 4129 1680 4163 1714
rect 4197 1680 4231 1714
rect 4265 1680 4299 1714
rect 4333 1680 4367 1714
rect 4401 1680 4435 1714
rect 4469 1680 4503 1714
rect 4537 1680 4571 1714
rect 4605 1680 4639 1714
rect 5433 3015 5467 3049
rect 5501 3015 5535 3049
rect 5569 3015 5603 3049
rect 5637 3015 5671 3049
rect 5705 3015 5739 3049
rect 5773 3015 5807 3049
rect 5841 3015 5875 3049
rect 5909 3015 5943 3049
rect 5977 3015 6011 3049
rect 6045 3015 6079 3049
rect 6113 3015 6147 3049
rect 6181 3015 6215 3049
rect 6249 3015 6283 3049
rect 6317 3015 6351 3049
rect 6385 3015 6419 3049
rect 6453 3015 6487 3049
rect 6521 3015 6555 3049
rect 6589 3015 6623 3049
rect 5357 2947 5391 2981
rect 5357 2879 5391 2913
rect 5357 2811 5391 2845
rect 5357 2743 5391 2777
rect 5357 2675 5391 2709
rect 5357 2607 5391 2641
rect 5357 2539 5391 2573
rect 5357 2471 5391 2505
rect 5357 2403 5391 2437
rect 5357 2335 5391 2369
rect 5357 2267 5391 2301
rect 5357 2199 5391 2233
rect 5357 2131 5391 2165
rect 5357 2063 5391 2097
rect 5357 1995 5391 2029
rect 5357 1927 5391 1961
rect 6657 2904 6691 2938
rect 6657 2836 6691 2870
rect 6657 2768 6691 2802
rect 6657 2700 6691 2734
rect 6657 2632 6691 2666
rect 6657 2564 6691 2598
rect 6657 2496 6691 2530
rect 6657 2428 6691 2462
rect 6657 2360 6691 2394
rect 6657 2292 6691 2326
rect 6657 2224 6691 2258
rect 6657 2156 6691 2190
rect 6657 2088 6691 2122
rect 6657 2020 6691 2054
rect 6657 1952 6691 1986
rect 5357 1859 5391 1893
rect 6657 1884 6691 1918
rect 5357 1754 5391 1788
rect 6657 1816 6691 1850
rect 6657 1748 6691 1782
rect 5425 1680 5459 1714
rect 5493 1680 5527 1714
rect 5561 1680 5595 1714
rect 5629 1680 5663 1714
rect 5697 1680 5731 1714
rect 5765 1680 5799 1714
rect 5833 1680 5867 1714
rect 5901 1680 5935 1714
rect 5969 1680 6003 1714
rect 6037 1680 6071 1714
rect 6105 1680 6139 1714
rect 6173 1680 6207 1714
rect 6241 1680 6275 1714
rect 6309 1680 6343 1714
rect 6377 1680 6411 1714
rect 6445 1680 6479 1714
rect 6513 1680 6547 1714
rect 6581 1680 6615 1714
rect 7299 3015 7333 3049
rect 7367 3015 7401 3049
rect 7435 3015 7469 3049
rect 7503 3015 7537 3049
rect 7571 3015 7605 3049
rect 7639 3015 7673 3049
rect 7707 3015 7741 3049
rect 7775 3015 7809 3049
rect 7843 3015 7877 3049
rect 7911 3015 7945 3049
rect 7979 3015 8013 3049
rect 8047 3015 8081 3049
rect 8115 3015 8149 3049
rect 8183 3015 8217 3049
rect 8251 3015 8285 3049
rect 8319 3015 8353 3049
rect 8387 3015 8421 3049
rect 8455 3015 8489 3049
rect 8523 3015 8557 3049
rect 8591 3015 8625 3049
rect 8659 3015 8693 3049
rect 8727 3015 8761 3049
rect 7225 2947 7259 2981
rect 7225 2879 7259 2913
rect 7225 2811 7259 2845
rect 7225 2743 7259 2777
rect 7225 2675 7259 2709
rect 7225 2607 7259 2641
rect 7225 2539 7259 2573
rect 7225 2471 7259 2505
rect 7225 2403 7259 2437
rect 7225 2335 7259 2369
rect 7225 2267 7259 2301
rect 7225 2199 7259 2233
rect 7225 2131 7259 2165
rect 7225 2063 7259 2097
rect 7225 1995 7259 2029
rect 7225 1927 7259 1961
rect 8795 2904 8829 2938
rect 8795 2836 8829 2870
rect 8795 2768 8829 2802
rect 8795 2700 8829 2734
rect 8795 2632 8829 2666
rect 8795 2564 8829 2598
rect 8795 2496 8829 2530
rect 8795 2428 8829 2462
rect 8795 2360 8829 2394
rect 8795 2292 8829 2326
rect 8795 2224 8829 2258
rect 8795 2156 8829 2190
rect 8795 2088 8829 2122
rect 8795 2020 8829 2054
rect 8795 1952 8829 1986
rect 7225 1859 7259 1893
rect 8795 1884 8829 1918
rect 7225 1754 7259 1788
rect 8795 1816 8829 1850
rect 8795 1748 8829 1782
rect 7293 1680 7327 1714
rect 7361 1680 7395 1714
rect 7429 1680 7463 1714
rect 7497 1680 7531 1714
rect 7565 1680 7599 1714
rect 7633 1680 7667 1714
rect 7701 1680 7735 1714
rect 7769 1680 7803 1714
rect 7837 1680 7871 1714
rect 7905 1680 7939 1714
rect 7973 1680 8007 1714
rect 8041 1680 8075 1714
rect 8109 1680 8143 1714
rect 8177 1680 8211 1714
rect 8245 1680 8279 1714
rect 8313 1680 8347 1714
rect 8381 1680 8415 1714
rect 8449 1680 8483 1714
rect 8517 1680 8551 1714
rect 8585 1680 8619 1714
rect 8653 1680 8687 1714
rect 8721 1680 8755 1714
rect 9571 3015 9605 3049
rect 9639 3015 9673 3049
rect 9707 3015 9741 3049
rect 9775 3015 9809 3049
rect 9843 3015 9877 3049
rect 9911 3015 9945 3049
rect 9979 3015 10013 3049
rect 10047 3015 10081 3049
rect 10115 3015 10149 3049
rect 10183 3015 10217 3049
rect 10251 3015 10285 3049
rect 10319 3015 10353 3049
rect 10387 3015 10421 3049
rect 10455 3015 10489 3049
rect 10523 3015 10557 3049
rect 10591 3015 10625 3049
rect 10659 3015 10693 3049
rect 10727 3015 10761 3049
rect 10795 3015 10829 3049
rect 10863 3015 10897 3049
rect 10931 3015 10965 3049
rect 10999 3015 11033 3049
rect 11067 3015 11101 3049
rect 11135 3015 11169 3049
rect 11203 3015 11237 3049
rect 11271 3015 11305 3049
rect 11339 3015 11373 3049
rect 11407 3015 11441 3049
rect 11475 3015 11509 3049
rect 11543 3015 11577 3049
rect 11611 3015 11645 3049
rect 9503 2904 9537 2938
rect 11695 2947 11729 2981
rect 9503 2836 9537 2870
rect 9503 2768 9537 2802
rect 9503 2700 9537 2734
rect 9503 2632 9537 2666
rect 9503 2564 9537 2598
rect 9503 2496 9537 2530
rect 9503 2428 9537 2462
rect 9503 2360 9537 2394
rect 9503 2292 9537 2326
rect 9503 2224 9537 2258
rect 9503 2156 9537 2190
rect 9503 2088 9537 2122
rect 9503 2020 9537 2054
rect 9503 1952 9537 1986
rect 11695 2879 11729 2913
rect 11695 2811 11729 2845
rect 11695 2743 11729 2777
rect 11695 2675 11729 2709
rect 11695 2607 11729 2641
rect 11695 2539 11729 2573
rect 11695 2471 11729 2505
rect 11695 2403 11729 2437
rect 11695 2335 11729 2369
rect 11695 2267 11729 2301
rect 11695 2199 11729 2233
rect 11695 2131 11729 2165
rect 11695 2063 11729 2097
rect 11695 1995 11729 2029
rect 9503 1884 9537 1918
rect 9503 1816 9537 1850
rect 11695 1828 11729 1862
rect 9503 1748 9537 1782
rect 11695 1760 11729 1794
rect 9587 1680 9621 1714
rect 9655 1680 9689 1714
rect 9723 1680 9757 1714
rect 9791 1680 9825 1714
rect 9859 1680 9893 1714
rect 9927 1680 9961 1714
rect 9995 1680 10029 1714
rect 10063 1680 10097 1714
rect 10131 1680 10165 1714
rect 10199 1680 10233 1714
rect 10267 1680 10301 1714
rect 10335 1680 10369 1714
rect 10403 1680 10437 1714
rect 10471 1680 10505 1714
rect 10539 1680 10573 1714
rect 10607 1680 10641 1714
rect 10675 1680 10709 1714
rect 10743 1680 10777 1714
rect 10811 1680 10845 1714
rect 10879 1680 10913 1714
rect 10947 1680 10981 1714
rect 11015 1680 11049 1714
rect 11083 1680 11117 1714
rect 11151 1680 11185 1714
rect 11219 1680 11253 1714
rect 11287 1680 11321 1714
rect 11355 1680 11389 1714
rect 11423 1680 11457 1714
rect 11491 1680 11525 1714
rect 11559 1680 11593 1714
rect 11627 1680 11661 1714
rect 12056 3030 12090 3064
rect 12124 3030 12158 3064
rect 12192 3030 12226 3064
rect 12260 3030 12294 3064
rect 12328 3030 12362 3064
rect 12396 3030 12430 3064
rect 12464 3030 12498 3064
rect 12532 3030 12566 3064
rect 12600 3030 12634 3064
rect 12668 3030 12702 3064
rect 12736 3030 12770 3064
rect 12804 3030 12838 3064
rect 12872 3030 12906 3064
rect 12940 3030 12974 3064
rect 13008 3030 13042 3064
rect 13076 3030 13110 3064
rect 13144 3030 13178 3064
rect 13212 3030 13246 3064
rect 13280 3030 13314 3064
rect 13348 3030 13382 3064
rect 13416 3030 13450 3064
rect 13484 3030 13518 3064
rect 13552 3030 13586 3064
rect 13620 3030 13654 3064
rect 13688 3030 13722 3064
rect 13756 3030 13790 3064
rect 13824 3030 13858 3064
rect 13892 3030 13926 3064
rect 13960 3030 13994 3064
rect 14028 3030 14062 3064
rect 14096 3030 14130 3064
rect 14164 3030 14198 3064
rect 14232 3030 14266 3064
rect 14300 3030 14334 3064
rect 14368 3030 14402 3064
rect 14436 3030 14470 3064
rect 14504 3030 14538 3064
rect 14572 3030 14606 3064
rect 14640 3030 14674 3064
rect 14708 3030 14742 3064
rect 14776 3030 14810 3064
rect 14844 3030 14878 3064
rect 14912 3030 14946 3064
rect 14980 3030 15014 3064
rect 15048 3030 15082 3064
rect 15116 3030 15150 3064
rect 15184 3030 15218 3064
rect 15252 3030 15286 3064
rect 15320 3030 15354 3064
rect 15388 3030 15422 3064
rect 15456 3030 15490 3064
rect 15524 3030 15558 3064
rect 15592 3030 15626 3064
rect 15660 3030 15694 3064
rect 15728 3030 15762 3064
rect 15796 3030 15830 3064
rect 15864 3030 15898 3064
rect 15932 3030 15966 3064
rect 16000 3030 16034 3064
rect 16068 3030 16102 3064
rect 16136 3030 16170 3064
rect 16204 3030 16238 3064
rect 16272 3030 16306 3064
rect 16340 3030 16374 3064
rect 16408 3030 16442 3064
rect 16476 3030 16510 3064
rect 16544 3030 16578 3064
rect 16612 3030 16646 3064
rect 16680 3030 16714 3064
rect 16748 3030 16782 3064
rect 16816 3030 16850 3064
rect 16884 3030 16918 3064
rect 16952 3030 16986 3064
rect 17020 3030 17054 3064
rect 11922 2962 11956 2996
rect 11922 2894 11956 2928
rect 11922 2826 11956 2860
rect 11922 2758 11956 2792
rect 14535 2962 14569 2996
rect 14535 2892 14569 2926
rect 14535 2822 14569 2856
rect 14535 2753 14569 2787
rect 17088 2942 17122 2976
rect 17088 2874 17122 2908
rect 17088 2806 17122 2840
rect 11922 2690 11956 2724
rect 14535 2684 14569 2718
rect 11922 2622 11956 2656
rect 17088 2738 17122 2772
rect 17088 2670 17122 2704
rect 14535 2615 14569 2649
rect 11922 2554 11956 2588
rect 11922 2486 11956 2520
rect 11922 2418 11956 2452
rect 11922 2350 11956 2384
rect 11922 2282 11956 2316
rect 11922 2214 11956 2248
rect 11922 2146 11956 2180
rect 11922 2078 11956 2112
rect 11922 2010 11956 2044
rect 11922 1942 11956 1976
rect 14535 2546 14569 2580
rect 14535 2477 14569 2511
rect 14535 2408 14569 2442
rect 14535 2339 14569 2373
rect 14535 2270 14569 2304
rect 14535 2201 14569 2235
rect 14535 2132 14569 2166
rect 14535 2063 14569 2097
rect 14535 1994 14569 2028
rect 17088 2602 17122 2636
rect 17088 2534 17122 2568
rect 17088 2466 17122 2500
rect 17088 2398 17122 2432
rect 17088 2330 17122 2364
rect 17088 2262 17122 2296
rect 17088 2194 17122 2228
rect 17088 2126 17122 2160
rect 17088 2058 17122 2092
rect 17088 1990 17122 2024
rect 14535 1925 14569 1959
rect 11922 1874 11956 1908
rect 11922 1742 11956 1776
rect 17088 1922 17122 1956
rect 14535 1856 14569 1890
rect 14535 1787 14569 1821
rect 14535 1718 14569 1752
rect 17088 1854 17122 1888
rect 17088 1786 17122 1820
rect 17088 1718 17122 1752
rect 11990 1650 12024 1684
rect 12058 1650 12092 1684
rect 12126 1650 12160 1684
rect 12194 1650 12228 1684
rect 12262 1650 12296 1684
rect 12330 1650 12364 1684
rect 12398 1650 12432 1684
rect 12466 1650 12500 1684
rect 12534 1650 12568 1684
rect 12602 1650 12636 1684
rect 12670 1650 12704 1684
rect 12738 1650 12772 1684
rect 12806 1650 12840 1684
rect 12874 1650 12908 1684
rect 12942 1650 12976 1684
rect 13010 1650 13044 1684
rect 13078 1650 13112 1684
rect 13146 1650 13180 1684
rect 13214 1650 13248 1684
rect 13282 1650 13316 1684
rect 13350 1650 13384 1684
rect 13418 1650 13452 1684
rect 13486 1650 13520 1684
rect 13554 1650 13588 1684
rect 13622 1650 13656 1684
rect 13690 1650 13724 1684
rect 13758 1650 13792 1684
rect 13826 1650 13860 1684
rect 13894 1650 13928 1684
rect 13962 1650 13996 1684
rect 14030 1650 14064 1684
rect 14098 1650 14132 1684
rect 14166 1650 14200 1684
rect 14234 1650 14268 1684
rect 14302 1650 14336 1684
rect 14370 1650 14404 1684
rect 14438 1650 14472 1684
rect 14506 1650 14540 1684
rect 14574 1650 14608 1684
rect 14642 1650 14676 1684
rect 14710 1650 14744 1684
rect 14778 1650 14812 1684
rect 14846 1650 14880 1684
rect 14914 1650 14948 1684
rect 14982 1650 15016 1684
rect 15050 1650 15084 1684
rect 15118 1650 15152 1684
rect 15186 1650 15220 1684
rect 15254 1650 15288 1684
rect 15322 1650 15356 1684
rect 15390 1650 15424 1684
rect 15458 1650 15492 1684
rect 15526 1650 15560 1684
rect 15594 1650 15628 1684
rect 15662 1650 15696 1684
rect 15730 1650 15764 1684
rect 15798 1650 15832 1684
rect 15866 1650 15900 1684
rect 15934 1650 15968 1684
rect 16002 1650 16036 1684
rect 16070 1650 16104 1684
rect 16138 1650 16172 1684
rect 16206 1650 16240 1684
rect 16274 1650 16308 1684
rect 16342 1650 16376 1684
rect 16410 1650 16444 1684
rect 16478 1650 16512 1684
rect 16546 1650 16580 1684
rect 16614 1650 16648 1684
rect 16682 1650 16716 1684
rect 16750 1650 16784 1684
rect 16818 1650 16852 1684
rect 16886 1650 16920 1684
rect 16954 1650 16988 1684
rect 1588 1032 1622 1066
rect 1656 1032 1690 1066
rect 1724 1032 1758 1066
rect 1792 1032 1826 1066
rect 1860 1032 1894 1066
rect 1928 1032 1962 1066
rect 1996 1032 2030 1066
rect 2064 1032 2098 1066
rect 2132 1032 2166 1066
rect 2200 1032 2234 1066
rect 2268 1032 2302 1066
rect 3023 1032 3057 1066
rect 3091 1032 3125 1066
rect 3159 1032 3193 1066
rect 3227 1032 3261 1066
rect 3295 1032 3329 1066
rect 3363 1032 3397 1066
<< poly >>
rect -56 2838 44 2870
rect -56 2206 44 2238
rect -71 2190 63 2206
rect -71 2156 -55 2190
rect -21 2156 13 2190
rect 47 2156 63 2190
rect -71 2140 63 2156
rect 765 2921 865 2953
rect 921 2921 1021 2953
rect 1187 2921 1287 2953
rect 1343 2921 1443 2953
rect 1499 2921 1599 2953
rect 1655 2921 1755 2953
rect 1811 2921 1911 2953
rect 1967 2921 2067 2953
rect 2123 2921 2223 2953
rect 2279 2921 2379 2953
rect 2435 2921 2535 2953
rect 2591 2921 2691 2953
rect 2747 2921 2847 2953
rect 2903 2921 3003 2953
rect 3059 2921 3159 2953
rect 3215 2921 3315 2953
rect 3371 2921 3471 2953
rect 3527 2921 3627 2953
rect 3683 2921 3783 2953
rect 3839 2921 3939 2953
rect 3995 2921 4095 2953
rect 4261 2603 4517 2619
rect 4261 2569 4277 2603
rect 4311 2569 4372 2603
rect 4406 2569 4467 2603
rect 4501 2569 4517 2603
rect 4261 2553 4517 2569
rect 4261 2521 4361 2553
rect 4417 2521 4517 2553
rect 765 1889 865 1921
rect 921 1889 1021 1921
rect 765 1873 1021 1889
rect 765 1839 781 1873
rect 815 1839 876 1873
rect 910 1839 971 1873
rect 1005 1839 1021 1873
rect 765 1823 1021 1839
rect 1187 1889 1287 1921
rect 1343 1889 1443 1921
rect 1499 1889 1599 1921
rect 1655 1889 1755 1921
rect 1811 1889 1911 1921
rect 1967 1889 2067 1921
rect 1187 1873 2067 1889
rect 1187 1839 1203 1873
rect 1237 1839 1277 1873
rect 1311 1839 1351 1873
rect 1385 1839 1425 1873
rect 1459 1839 1499 1873
rect 1533 1839 1573 1873
rect 1607 1839 1647 1873
rect 1681 1839 1721 1873
rect 1755 1839 1795 1873
rect 1829 1839 1869 1873
rect 1903 1839 1943 1873
rect 1977 1839 2017 1873
rect 2051 1839 2067 1873
rect 1187 1823 2067 1839
rect 2123 1889 2223 1921
rect 2279 1889 2379 1921
rect 2435 1889 2535 1921
rect 2591 1889 2691 1921
rect 2123 1873 2691 1889
rect 2123 1839 2139 1873
rect 2173 1839 2210 1873
rect 2244 1839 2281 1873
rect 2315 1839 2353 1873
rect 2387 1839 2425 1873
rect 2459 1839 2497 1873
rect 2531 1839 2569 1873
rect 2603 1839 2641 1873
rect 2675 1839 2691 1873
rect 2123 1823 2691 1839
rect 2747 1889 2847 1921
rect 2903 1889 3003 1921
rect 3059 1889 3159 1921
rect 3215 1889 3315 1921
rect 2747 1873 3315 1889
rect 2747 1839 2763 1873
rect 2797 1839 2835 1873
rect 2869 1839 2907 1873
rect 2941 1839 2979 1873
rect 3013 1839 3051 1873
rect 3085 1839 3123 1873
rect 3157 1839 3194 1873
rect 3228 1839 3265 1873
rect 3299 1839 3315 1873
rect 2747 1823 3315 1839
rect 3371 1889 3471 1921
rect 3527 1889 3627 1921
rect 3683 1889 3783 1921
rect 3839 1889 3939 1921
rect 3995 1889 4095 1921
rect 4261 1889 4361 1921
rect 4417 1889 4517 1921
rect 3371 1873 4095 1889
rect 3371 1839 3387 1873
rect 3421 1839 3461 1873
rect 3495 1839 3534 1873
rect 3568 1839 3607 1873
rect 3641 1839 3680 1873
rect 3714 1839 3753 1873
rect 3787 1839 3826 1873
rect 3860 1839 3899 1873
rect 3933 1839 3972 1873
rect 4006 1839 4045 1873
rect 4079 1839 4095 1873
rect 3371 1823 4095 1839
rect 5547 2921 5647 2953
rect 5703 2921 5803 2953
rect 5859 2921 6019 2953
rect 6075 2921 6235 2953
rect 6401 2521 6501 2553
rect 6401 2289 6501 2321
rect 6401 2273 6535 2289
rect 6401 2239 6417 2273
rect 6451 2239 6485 2273
rect 6519 2239 6535 2273
rect 6401 2223 6535 2239
rect 5547 1889 5647 1921
rect 5703 1889 5803 1921
rect 5547 1873 5803 1889
rect 5547 1839 5563 1873
rect 5597 1839 5658 1873
rect 5692 1839 5753 1873
rect 5787 1839 5803 1873
rect 5547 1823 5803 1839
rect 5859 1889 6019 1921
rect 6075 1889 6235 1921
rect 5859 1873 6235 1889
rect 5859 1839 5875 1873
rect 5909 1839 5953 1873
rect 5987 1839 6031 1873
rect 6065 1839 6108 1873
rect 6142 1839 6185 1873
rect 6219 1839 6235 1873
rect 5859 1823 6235 1839
rect 7415 2921 7575 2953
rect 7631 2921 7791 2953
rect 7847 2921 8007 2953
rect 8063 2921 8163 2953
rect 8219 2921 8319 2953
rect 8375 2921 8475 2953
rect 8531 2921 8631 2953
rect 7415 1889 7575 1921
rect 7631 1889 7791 1921
rect 7847 1889 8007 1921
rect 7415 1873 8007 1889
rect 7415 1839 7431 1873
rect 7465 1839 7507 1873
rect 7541 1839 7582 1873
rect 7616 1839 7657 1873
rect 7691 1839 7732 1873
rect 7766 1839 7807 1873
rect 7841 1839 7882 1873
rect 7916 1839 7957 1873
rect 7991 1839 8007 1873
rect 7415 1823 8007 1839
rect 8063 1889 8163 1921
rect 8219 1889 8319 1921
rect 8375 1889 8475 1921
rect 8531 1889 8631 1921
rect 8063 1873 8631 1889
rect 8063 1839 8079 1873
rect 8113 1839 8151 1873
rect 8185 1839 8223 1873
rect 8257 1839 8295 1873
rect 8329 1839 8367 1873
rect 8401 1839 8439 1873
rect 8473 1839 8510 1873
rect 8544 1839 8581 1873
rect 8615 1839 8631 1873
rect 8063 1823 8631 1839
rect 9693 2921 9793 2953
rect 9849 2921 9949 2953
rect 10005 2921 10105 2953
rect 10161 2921 10261 2953
rect 10317 2921 10417 2953
rect 10473 2921 10573 2953
rect 10629 2921 10729 2953
rect 10785 2921 10885 2953
rect 10941 2921 11041 2953
rect 11097 2921 11197 2953
rect 11253 2921 11353 2953
rect 11409 2921 11509 2953
rect 9693 1889 9793 1921
rect 9849 1889 9949 1921
rect 9693 1873 9949 1889
rect 9693 1839 9709 1873
rect 9743 1839 9804 1873
rect 9838 1839 9899 1873
rect 9933 1839 9949 1873
rect 9693 1823 9949 1839
rect 10005 1889 10105 1921
rect 10161 1889 10261 1921
rect 10317 1889 10417 1921
rect 10473 1889 10573 1921
rect 10629 1889 10729 1921
rect 10785 1889 10885 1921
rect 10941 1889 11041 1921
rect 11097 1889 11197 1921
rect 10005 1873 10886 1889
rect 10005 1839 10021 1873
rect 10055 1839 10096 1873
rect 10130 1839 10170 1873
rect 10204 1839 10244 1873
rect 10278 1839 10318 1873
rect 10352 1839 10392 1873
rect 10426 1839 10466 1873
rect 10500 1839 10540 1873
rect 10574 1839 10614 1873
rect 10648 1839 10688 1873
rect 10722 1839 10762 1873
rect 10796 1839 10836 1873
rect 10870 1839 10886 1873
rect 10005 1823 10886 1839
rect 10941 1873 11197 1889
rect 10941 1839 10957 1873
rect 10991 1839 11052 1873
rect 11086 1839 11147 1873
rect 11181 1839 11197 1873
rect 10941 1823 11197 1839
rect 11253 1889 11353 1921
rect 11409 1889 11509 1921
rect 11253 1873 11509 1889
rect 11253 1839 11269 1873
rect 11303 1839 11364 1873
rect 11398 1839 11459 1873
rect 11493 1839 11509 1873
rect 11253 1823 11509 1839
rect 12186 2435 12218 2615
rect 14218 2599 14316 2615
rect 14218 2565 14266 2599
rect 14300 2565 14316 2599
rect 14218 2526 14316 2565
rect 14218 2492 14266 2526
rect 14300 2492 14316 2526
rect 14218 2453 14316 2492
rect 14218 2435 14266 2453
rect 14250 2419 14266 2435
rect 14300 2419 14316 2453
rect 14250 2380 14316 2419
rect 14250 2379 14266 2380
rect 12186 2199 12218 2379
rect 14218 2346 14266 2379
rect 14300 2346 14316 2380
rect 14218 2307 14316 2346
rect 14218 2273 14266 2307
rect 14300 2273 14316 2307
rect 14218 2234 14316 2273
rect 14218 2200 14266 2234
rect 14300 2200 14316 2234
rect 14218 2199 14316 2200
rect 14250 2161 14316 2199
rect 14250 2143 14266 2161
rect 12186 1963 12218 2143
rect 14218 2127 14266 2143
rect 14300 2127 14316 2161
rect 14218 2087 14316 2127
rect 14218 2053 14266 2087
rect 14300 2053 14316 2087
rect 14218 2013 14316 2053
rect 14218 1979 14266 2013
rect 14300 1979 14316 2013
rect 14218 1963 14316 1979
rect 14764 2599 14862 2615
rect 14764 2565 14780 2599
rect 14814 2565 14862 2599
rect 14764 2526 14862 2565
rect 14764 2492 14780 2526
rect 14814 2492 14862 2526
rect 14764 2453 14862 2492
rect 14764 2419 14780 2453
rect 14814 2435 14862 2453
rect 16862 2435 16894 2615
rect 14814 2419 14830 2435
rect 14764 2380 14830 2419
rect 14764 2346 14780 2380
rect 14814 2379 14830 2380
rect 14814 2346 14862 2379
rect 14764 2307 14862 2346
rect 14764 2273 14780 2307
rect 14814 2273 14862 2307
rect 14764 2234 14862 2273
rect 14764 2200 14780 2234
rect 14814 2200 14862 2234
rect 14764 2199 14862 2200
rect 16862 2199 16894 2379
rect 14764 2161 14830 2199
rect 14764 2127 14780 2161
rect 14814 2143 14830 2161
rect 14814 2127 14862 2143
rect 14764 2087 14862 2127
rect 14764 2053 14780 2087
rect 14814 2053 14862 2087
rect 14764 2013 14862 2053
rect 14764 1979 14780 2013
rect 14814 1979 14862 2013
rect 14764 1963 14862 1979
rect 16862 1963 16894 2143
rect 3987 1230 5627 1246
rect 3987 1196 4003 1230
rect 4037 1196 4072 1230
rect 4106 1196 4141 1230
rect 4175 1196 4210 1230
rect 4244 1196 4279 1230
rect 4313 1196 4348 1230
rect 4382 1196 4417 1230
rect 4451 1196 4486 1230
rect 4520 1196 4555 1230
rect 4589 1196 4624 1230
rect 4658 1196 4693 1230
rect 4727 1196 4761 1230
rect 4795 1196 4829 1230
rect 4863 1196 4897 1230
rect 4931 1196 4965 1230
rect 4999 1196 5033 1230
rect 5067 1196 5101 1230
rect 5135 1196 5169 1230
rect 5203 1196 5237 1230
rect 5271 1196 5305 1230
rect 5339 1196 5373 1230
rect 5407 1196 5441 1230
rect 5475 1196 5509 1230
rect 5543 1196 5577 1230
rect 5611 1196 5627 1230
rect 3987 1180 5627 1196
rect 6703 1230 6959 1246
rect 6703 1196 6719 1230
rect 6753 1196 6814 1230
rect 6848 1196 6909 1230
rect 6943 1196 6959 1230
rect 6703 1180 6959 1196
rect 3987 1148 4037 1180
rect 4093 1148 4143 1180
rect 4199 1148 4249 1180
rect 4305 1148 4355 1180
rect 4411 1148 4461 1180
rect 4517 1148 4567 1180
rect 4623 1148 4673 1180
rect 4729 1148 4779 1180
rect 4835 1148 4885 1180
rect 4941 1148 4991 1180
rect 5047 1148 5097 1180
rect 5153 1148 5203 1180
rect 5259 1148 5309 1180
rect 5365 1148 5415 1180
rect 5471 1148 5521 1180
rect 5577 1148 5627 1180
rect 5945 1148 6105 1180
rect 6161 1148 6321 1180
rect 6377 1148 6537 1180
rect 6703 1148 6803 1180
rect 6859 1148 6959 1180
rect 7015 1230 7149 1246
rect 7015 1196 7031 1230
rect 7065 1196 7099 1230
rect 7133 1196 7149 1230
rect 7015 1180 7149 1196
rect 7281 1230 7415 1246
rect 7281 1196 7297 1230
rect 7331 1196 7365 1230
rect 7399 1196 7415 1230
rect 7281 1180 7415 1196
rect 7547 1230 8571 1246
rect 7547 1196 7563 1230
rect 7597 1196 7631 1230
rect 7665 1196 7699 1230
rect 7733 1196 7767 1230
rect 7801 1196 7835 1230
rect 7869 1196 7903 1230
rect 7937 1196 7971 1230
rect 8005 1196 8039 1230
rect 8073 1196 8107 1230
rect 8141 1196 8176 1230
rect 8210 1196 8245 1230
rect 8279 1196 8314 1230
rect 8348 1196 8383 1230
rect 8417 1196 8452 1230
rect 8486 1196 8521 1230
rect 8555 1196 8571 1230
rect 7547 1180 8571 1196
rect 7015 1148 7115 1180
rect 7281 1148 7381 1180
rect 7547 1148 7707 1180
rect 7763 1148 7923 1180
rect 7979 1148 8139 1180
rect 8195 1148 8355 1180
rect 8411 1148 8571 1180
rect 8627 1230 11163 1246
rect 8627 1196 8643 1230
rect 8677 1196 8711 1230
rect 8745 1196 8779 1230
rect 8813 1196 8847 1230
rect 8881 1196 8915 1230
rect 8949 1196 8983 1230
rect 9017 1196 9051 1230
rect 9085 1196 9119 1230
rect 9153 1196 9187 1230
rect 9221 1196 9255 1230
rect 9289 1196 9323 1230
rect 9357 1196 9391 1230
rect 9425 1196 9459 1230
rect 9493 1196 9527 1230
rect 9561 1196 9595 1230
rect 9629 1196 9664 1230
rect 9698 1196 9733 1230
rect 9767 1196 9802 1230
rect 9836 1196 9871 1230
rect 9905 1196 9940 1230
rect 9974 1196 10009 1230
rect 10043 1196 10078 1230
rect 10112 1196 10147 1230
rect 10181 1196 10216 1230
rect 10250 1196 10285 1230
rect 10319 1196 10354 1230
rect 10388 1196 10423 1230
rect 10457 1196 10492 1230
rect 10526 1196 10561 1230
rect 10595 1196 10630 1230
rect 10664 1196 10699 1230
rect 10733 1196 10768 1230
rect 10802 1196 10837 1230
rect 10871 1196 10906 1230
rect 10940 1196 10975 1230
rect 11009 1196 11044 1230
rect 11078 1196 11113 1230
rect 11147 1196 11163 1230
rect 8627 1180 11163 1196
rect 8627 1148 8787 1180
rect 8843 1148 9003 1180
rect 9059 1148 9219 1180
rect 9275 1148 9435 1180
rect 9491 1148 9651 1180
rect 9707 1148 9867 1180
rect 9923 1148 10083 1180
rect 10139 1148 10299 1180
rect 10355 1148 10515 1180
rect 10571 1148 10731 1180
rect 10787 1148 10947 1180
rect 11003 1148 11163 1180
rect 11219 1230 15051 1246
rect 11219 1196 11235 1230
rect 11269 1196 11303 1230
rect 11337 1196 11371 1230
rect 11405 1196 11439 1230
rect 11473 1196 11507 1230
rect 11541 1196 11575 1230
rect 11609 1196 11643 1230
rect 11677 1196 11711 1230
rect 11745 1196 11779 1230
rect 11813 1196 11847 1230
rect 11881 1196 11915 1230
rect 11949 1196 11983 1230
rect 12017 1196 12051 1230
rect 12085 1196 12119 1230
rect 12153 1196 12187 1230
rect 12221 1196 12255 1230
rect 12289 1196 12323 1230
rect 12357 1196 12391 1230
rect 12425 1196 12459 1230
rect 12493 1196 12527 1230
rect 12561 1196 12595 1230
rect 12629 1196 12663 1230
rect 12697 1196 12731 1230
rect 12765 1196 12799 1230
rect 12833 1196 12867 1230
rect 12901 1196 12935 1230
rect 12969 1196 13003 1230
rect 13037 1196 13071 1230
rect 13105 1196 13139 1230
rect 13173 1196 13207 1230
rect 13241 1196 13276 1230
rect 13310 1196 13345 1230
rect 13379 1196 13414 1230
rect 13448 1196 13483 1230
rect 13517 1196 13552 1230
rect 13586 1196 13621 1230
rect 13655 1196 13690 1230
rect 13724 1196 13759 1230
rect 13793 1196 13828 1230
rect 13862 1196 13897 1230
rect 13931 1196 13966 1230
rect 14000 1196 14035 1230
rect 14069 1196 14104 1230
rect 14138 1196 14173 1230
rect 14207 1196 14242 1230
rect 14276 1196 14311 1230
rect 14345 1196 14380 1230
rect 14414 1196 14449 1230
rect 14483 1196 14518 1230
rect 14552 1196 14587 1230
rect 14621 1196 14656 1230
rect 14690 1196 14725 1230
rect 14759 1196 14794 1230
rect 14828 1196 14863 1230
rect 14897 1196 14932 1230
rect 14966 1196 15001 1230
rect 15035 1196 15051 1230
rect 11219 1180 15051 1196
rect 11219 1148 11379 1180
rect 11435 1148 11595 1180
rect 11651 1148 11811 1180
rect 11867 1148 12027 1180
rect 12083 1148 12243 1180
rect 12299 1148 12459 1180
rect 12515 1148 12675 1180
rect 12731 1148 12891 1180
rect 12947 1148 13107 1180
rect 13163 1148 13323 1180
rect 13379 1148 13539 1180
rect 13595 1148 13755 1180
rect 13811 1148 13971 1180
rect 14027 1148 14187 1180
rect 14243 1148 14403 1180
rect 14459 1148 14619 1180
rect 14675 1148 14835 1180
rect 14891 1148 15051 1180
rect 15217 1230 15417 1246
rect 15217 1196 15233 1230
rect 15267 1196 15367 1230
rect 15401 1196 15417 1230
rect 15217 1148 15417 1196
rect 15583 1230 15959 1246
rect 15583 1196 15599 1230
rect 15633 1196 15677 1230
rect 15711 1196 15755 1230
rect 15789 1196 15832 1230
rect 15866 1196 15909 1230
rect 15943 1196 15959 1230
rect 15583 1180 15959 1196
rect 15583 1148 15743 1180
rect 15799 1148 15959 1180
rect 5945 916 6105 948
rect 6161 916 6321 948
rect 6377 916 6537 948
rect 5945 900 6537 916
rect 5945 866 5961 900
rect 5995 866 6037 900
rect 6071 866 6112 900
rect 6146 866 6187 900
rect 6221 866 6262 900
rect 6296 866 6337 900
rect 6371 866 6412 900
rect 6446 866 6487 900
rect 6521 866 6537 900
rect 5945 850 6537 866
rect 5945 818 6105 850
rect 6161 818 6321 850
rect 6377 818 6537 850
rect 5945 586 6105 618
rect 6161 586 6321 618
rect 6377 586 6537 618
rect 5945 528 6537 544
rect 5945 494 5961 528
rect 5995 494 6037 528
rect 6071 494 6112 528
rect 6146 494 6187 528
rect 6221 494 6262 528
rect 6296 494 6337 528
rect 6371 494 6412 528
rect 6446 494 6487 528
rect 6521 494 6537 528
rect 6703 516 6803 548
rect 6859 516 6959 548
rect 7015 516 7115 548
rect 5945 478 6537 494
rect 5945 446 6105 478
rect 6161 446 6321 478
rect 6377 446 6537 478
rect 5945 214 6105 246
rect 6161 214 6321 246
rect 6377 214 6537 246
rect 15217 516 15417 548
rect 3987 116 4037 148
rect 4093 116 4143 148
rect 4199 116 4249 148
rect 4305 116 4355 148
rect 4411 116 4461 148
rect 4517 116 4567 148
rect 4623 116 4673 148
rect 4729 116 4779 148
rect 4835 116 4885 148
rect 4941 116 4991 148
rect 5047 116 5097 148
rect 5153 116 5203 148
rect 5259 116 5309 148
rect 5365 116 5415 148
rect 5471 116 5521 148
rect 5577 116 5627 148
rect 7281 116 7381 148
rect 7547 116 7707 148
rect 7763 116 7923 148
rect 7979 116 8139 148
rect 8195 116 8355 148
rect 8411 116 8571 148
rect 8627 116 8787 148
rect 8843 116 9003 148
rect 9059 116 9219 148
rect 9275 116 9435 148
rect 9491 116 9651 148
rect 9707 116 9867 148
rect 9923 116 10083 148
rect 10139 116 10299 148
rect 10355 116 10515 148
rect 10571 116 10731 148
rect 10787 116 10947 148
rect 11003 116 11163 148
rect 11219 116 11379 148
rect 11435 116 11595 148
rect 11651 116 11811 148
rect 11867 116 12027 148
rect 12083 116 12243 148
rect 12299 116 12459 148
rect 12515 116 12675 148
rect 12731 116 12891 148
rect 12947 116 13107 148
rect 13163 116 13323 148
rect 13379 116 13539 148
rect 13595 116 13755 148
rect 13811 116 13971 148
rect 14027 116 14187 148
rect 14243 116 14403 148
rect 14459 116 14619 148
rect 14675 116 14835 148
rect 14891 116 15051 148
rect 15583 116 15743 148
rect 15799 116 15959 148
<< polycont >>
rect -55 2156 -21 2190
rect 13 2156 47 2190
rect 4277 2569 4311 2603
rect 4372 2569 4406 2603
rect 4467 2569 4501 2603
rect 781 1839 815 1873
rect 876 1839 910 1873
rect 971 1839 1005 1873
rect 1203 1839 1237 1873
rect 1277 1839 1311 1873
rect 1351 1839 1385 1873
rect 1425 1839 1459 1873
rect 1499 1839 1533 1873
rect 1573 1839 1607 1873
rect 1647 1839 1681 1873
rect 1721 1839 1755 1873
rect 1795 1839 1829 1873
rect 1869 1839 1903 1873
rect 1943 1839 1977 1873
rect 2017 1839 2051 1873
rect 2139 1839 2173 1873
rect 2210 1839 2244 1873
rect 2281 1839 2315 1873
rect 2353 1839 2387 1873
rect 2425 1839 2459 1873
rect 2497 1839 2531 1873
rect 2569 1839 2603 1873
rect 2641 1839 2675 1873
rect 2763 1839 2797 1873
rect 2835 1839 2869 1873
rect 2907 1839 2941 1873
rect 2979 1839 3013 1873
rect 3051 1839 3085 1873
rect 3123 1839 3157 1873
rect 3194 1839 3228 1873
rect 3265 1839 3299 1873
rect 3387 1839 3421 1873
rect 3461 1839 3495 1873
rect 3534 1839 3568 1873
rect 3607 1839 3641 1873
rect 3680 1839 3714 1873
rect 3753 1839 3787 1873
rect 3826 1839 3860 1873
rect 3899 1839 3933 1873
rect 3972 1839 4006 1873
rect 4045 1839 4079 1873
rect 6417 2239 6451 2273
rect 6485 2239 6519 2273
rect 5563 1839 5597 1873
rect 5658 1839 5692 1873
rect 5753 1839 5787 1873
rect 5875 1839 5909 1873
rect 5953 1839 5987 1873
rect 6031 1839 6065 1873
rect 6108 1839 6142 1873
rect 6185 1839 6219 1873
rect 7431 1839 7465 1873
rect 7507 1839 7541 1873
rect 7582 1839 7616 1873
rect 7657 1839 7691 1873
rect 7732 1839 7766 1873
rect 7807 1839 7841 1873
rect 7882 1839 7916 1873
rect 7957 1839 7991 1873
rect 8079 1839 8113 1873
rect 8151 1839 8185 1873
rect 8223 1839 8257 1873
rect 8295 1839 8329 1873
rect 8367 1839 8401 1873
rect 8439 1839 8473 1873
rect 8510 1839 8544 1873
rect 8581 1839 8615 1873
rect 9709 1839 9743 1873
rect 9804 1839 9838 1873
rect 9899 1839 9933 1873
rect 10021 1839 10055 1873
rect 10096 1839 10130 1873
rect 10170 1839 10204 1873
rect 10244 1839 10278 1873
rect 10318 1839 10352 1873
rect 10392 1839 10426 1873
rect 10466 1839 10500 1873
rect 10540 1839 10574 1873
rect 10614 1839 10648 1873
rect 10688 1839 10722 1873
rect 10762 1839 10796 1873
rect 10836 1839 10870 1873
rect 10957 1839 10991 1873
rect 11052 1839 11086 1873
rect 11147 1839 11181 1873
rect 11269 1839 11303 1873
rect 11364 1839 11398 1873
rect 11459 1839 11493 1873
rect 14266 2565 14300 2599
rect 14266 2492 14300 2526
rect 14266 2419 14300 2453
rect 14266 2346 14300 2380
rect 14266 2273 14300 2307
rect 14266 2200 14300 2234
rect 14266 2127 14300 2161
rect 14266 2053 14300 2087
rect 14266 1979 14300 2013
rect 14780 2565 14814 2599
rect 14780 2492 14814 2526
rect 14780 2419 14814 2453
rect 14780 2346 14814 2380
rect 14780 2273 14814 2307
rect 14780 2200 14814 2234
rect 14780 2127 14814 2161
rect 14780 2053 14814 2087
rect 14780 1979 14814 2013
rect 4003 1196 4037 1230
rect 4072 1196 4106 1230
rect 4141 1196 4175 1230
rect 4210 1196 4244 1230
rect 4279 1196 4313 1230
rect 4348 1196 4382 1230
rect 4417 1196 4451 1230
rect 4486 1196 4520 1230
rect 4555 1196 4589 1230
rect 4624 1196 4658 1230
rect 4693 1196 4727 1230
rect 4761 1196 4795 1230
rect 4829 1196 4863 1230
rect 4897 1196 4931 1230
rect 4965 1196 4999 1230
rect 5033 1196 5067 1230
rect 5101 1196 5135 1230
rect 5169 1196 5203 1230
rect 5237 1196 5271 1230
rect 5305 1196 5339 1230
rect 5373 1196 5407 1230
rect 5441 1196 5475 1230
rect 5509 1196 5543 1230
rect 5577 1196 5611 1230
rect 6719 1196 6753 1230
rect 6814 1196 6848 1230
rect 6909 1196 6943 1230
rect 7031 1196 7065 1230
rect 7099 1196 7133 1230
rect 7297 1196 7331 1230
rect 7365 1196 7399 1230
rect 7563 1196 7597 1230
rect 7631 1196 7665 1230
rect 7699 1196 7733 1230
rect 7767 1196 7801 1230
rect 7835 1196 7869 1230
rect 7903 1196 7937 1230
rect 7971 1196 8005 1230
rect 8039 1196 8073 1230
rect 8107 1196 8141 1230
rect 8176 1196 8210 1230
rect 8245 1196 8279 1230
rect 8314 1196 8348 1230
rect 8383 1196 8417 1230
rect 8452 1196 8486 1230
rect 8521 1196 8555 1230
rect 8643 1196 8677 1230
rect 8711 1196 8745 1230
rect 8779 1196 8813 1230
rect 8847 1196 8881 1230
rect 8915 1196 8949 1230
rect 8983 1196 9017 1230
rect 9051 1196 9085 1230
rect 9119 1196 9153 1230
rect 9187 1196 9221 1230
rect 9255 1196 9289 1230
rect 9323 1196 9357 1230
rect 9391 1196 9425 1230
rect 9459 1196 9493 1230
rect 9527 1196 9561 1230
rect 9595 1196 9629 1230
rect 9664 1196 9698 1230
rect 9733 1196 9767 1230
rect 9802 1196 9836 1230
rect 9871 1196 9905 1230
rect 9940 1196 9974 1230
rect 10009 1196 10043 1230
rect 10078 1196 10112 1230
rect 10147 1196 10181 1230
rect 10216 1196 10250 1230
rect 10285 1196 10319 1230
rect 10354 1196 10388 1230
rect 10423 1196 10457 1230
rect 10492 1196 10526 1230
rect 10561 1196 10595 1230
rect 10630 1196 10664 1230
rect 10699 1196 10733 1230
rect 10768 1196 10802 1230
rect 10837 1196 10871 1230
rect 10906 1196 10940 1230
rect 10975 1196 11009 1230
rect 11044 1196 11078 1230
rect 11113 1196 11147 1230
rect 11235 1196 11269 1230
rect 11303 1196 11337 1230
rect 11371 1196 11405 1230
rect 11439 1196 11473 1230
rect 11507 1196 11541 1230
rect 11575 1196 11609 1230
rect 11643 1196 11677 1230
rect 11711 1196 11745 1230
rect 11779 1196 11813 1230
rect 11847 1196 11881 1230
rect 11915 1196 11949 1230
rect 11983 1196 12017 1230
rect 12051 1196 12085 1230
rect 12119 1196 12153 1230
rect 12187 1196 12221 1230
rect 12255 1196 12289 1230
rect 12323 1196 12357 1230
rect 12391 1196 12425 1230
rect 12459 1196 12493 1230
rect 12527 1196 12561 1230
rect 12595 1196 12629 1230
rect 12663 1196 12697 1230
rect 12731 1196 12765 1230
rect 12799 1196 12833 1230
rect 12867 1196 12901 1230
rect 12935 1196 12969 1230
rect 13003 1196 13037 1230
rect 13071 1196 13105 1230
rect 13139 1196 13173 1230
rect 13207 1196 13241 1230
rect 13276 1196 13310 1230
rect 13345 1196 13379 1230
rect 13414 1196 13448 1230
rect 13483 1196 13517 1230
rect 13552 1196 13586 1230
rect 13621 1196 13655 1230
rect 13690 1196 13724 1230
rect 13759 1196 13793 1230
rect 13828 1196 13862 1230
rect 13897 1196 13931 1230
rect 13966 1196 14000 1230
rect 14035 1196 14069 1230
rect 14104 1196 14138 1230
rect 14173 1196 14207 1230
rect 14242 1196 14276 1230
rect 14311 1196 14345 1230
rect 14380 1196 14414 1230
rect 14449 1196 14483 1230
rect 14518 1196 14552 1230
rect 14587 1196 14621 1230
rect 14656 1196 14690 1230
rect 14725 1196 14759 1230
rect 14794 1196 14828 1230
rect 14863 1196 14897 1230
rect 14932 1196 14966 1230
rect 15001 1196 15035 1230
rect 15233 1196 15267 1230
rect 15367 1196 15401 1230
rect 15599 1196 15633 1230
rect 15677 1196 15711 1230
rect 15755 1196 15789 1230
rect 15832 1196 15866 1230
rect 15909 1196 15943 1230
rect 5961 866 5995 900
rect 6037 866 6071 900
rect 6112 866 6146 900
rect 6187 866 6221 900
rect 6262 866 6296 900
rect 6337 866 6371 900
rect 6412 866 6446 900
rect 6487 866 6521 900
rect 5961 494 5995 528
rect 6037 494 6071 528
rect 6112 494 6146 528
rect 6187 494 6221 528
rect 6262 494 6296 528
rect 6337 494 6371 528
rect 6412 494 6446 528
rect 6487 494 6521 528
<< locali >>
rect 204 3272 4936 3278
rect 6993 3272 9058 3278
rect 204 3238 278 3272
rect 326 3238 346 3272
rect 408 3238 414 3272
rect 448 3238 456 3272
rect 516 3238 538 3272
rect 584 3238 618 3272
rect 682 3238 686 3272
rect 788 3238 792 3272
rect 856 3238 864 3272
rect 924 3238 936 3272
rect 992 3238 1008 3272
rect 1060 3238 1080 3272
rect 1128 3238 1152 3272
rect 1196 3238 1224 3272
rect 1264 3238 1296 3272
rect 1332 3238 1366 3272
rect 1402 3238 1434 3272
rect 1474 3238 1502 3272
rect 1546 3238 1570 3272
rect 1618 3238 1638 3272
rect 1690 3238 1706 3272
rect 1762 3238 1774 3272
rect 1834 3238 1842 3272
rect 1906 3238 1910 3272
rect 2012 3238 2016 3272
rect 2080 3238 2088 3272
rect 2148 3238 2160 3272
rect 2216 3238 2232 3272
rect 2284 3238 2304 3272
rect 2352 3238 2376 3272
rect 2420 3238 2448 3272
rect 2488 3238 2520 3272
rect 2556 3238 2590 3272
rect 2626 3238 2658 3272
rect 2698 3238 2726 3272
rect 2770 3238 2794 3272
rect 2842 3238 2862 3272
rect 2914 3238 2930 3272
rect 2986 3238 2998 3272
rect 3058 3238 3066 3272
rect 3130 3238 3134 3272
rect 3236 3238 3240 3272
rect 3304 3238 3312 3272
rect 3372 3238 3384 3272
rect 3440 3238 3456 3272
rect 3508 3238 3528 3272
rect 3576 3238 3600 3272
rect 3644 3238 3672 3272
rect 3712 3238 3744 3272
rect 3780 3238 3814 3272
rect 3850 3238 3882 3272
rect 3922 3238 3950 3272
rect 3994 3238 4018 3272
rect 4066 3238 4086 3272
rect 4138 3238 4154 3272
rect 4210 3238 4222 3272
rect 4282 3238 4290 3272
rect 4354 3238 4358 3272
rect 4460 3238 4464 3272
rect 4528 3238 4536 3272
rect 4596 3238 4608 3272
rect 4664 3238 4680 3272
rect 4732 3238 4752 3272
rect 4800 3238 4824 3272
rect 4858 3238 4936 3272
rect 204 3232 4936 3238
rect 204 3200 250 3232
rect 204 3157 210 3200
rect 244 3157 250 3200
rect 204 3123 250 3157
rect 204 3079 210 3123
rect 244 3079 250 3123
rect 204 3055 250 3079
rect 4890 3204 4936 3232
rect 4890 3164 4896 3204
rect 4930 3164 4936 3204
rect 4890 3136 4936 3164
rect 4890 3090 4896 3136
rect 4930 3090 4936 3136
rect 4890 3068 4936 3090
rect 204 2992 210 3055
rect 244 2992 250 3055
rect 204 2987 250 2992
rect 204 2953 210 2987
rect 244 2953 250 2987
rect 204 2939 250 2953
rect 204 2885 210 2939
rect 244 2885 250 2939
rect 204 2858 250 2885
rect 193 2851 250 2858
rect 193 2817 210 2851
rect 244 2817 250 2851
rect 193 2812 250 2817
rect 427 3049 4713 3055
rect 427 3015 501 3049
rect 539 3015 569 3049
rect 611 3015 637 3049
rect 683 3015 705 3049
rect 755 3015 773 3049
rect 828 3015 841 3049
rect 901 3015 909 3049
rect 974 3015 977 3049
rect 1011 3015 1013 3049
rect 1079 3015 1086 3049
rect 1147 3015 1159 3049
rect 1215 3015 1232 3049
rect 1283 3015 1305 3049
rect 1351 3015 1378 3049
rect 1419 3015 1451 3049
rect 1487 3015 1521 3049
rect 1558 3015 1589 3049
rect 1631 3015 1657 3049
rect 1704 3015 1725 3049
rect 1777 3015 1793 3049
rect 1850 3015 1861 3049
rect 1923 3015 1929 3049
rect 1996 3015 1997 3049
rect 2031 3015 2035 3049
rect 2099 3015 2108 3049
rect 2167 3015 2181 3049
rect 2235 3015 2254 3049
rect 2303 3015 2327 3049
rect 2371 3015 2400 3049
rect 2439 3015 2473 3049
rect 2507 3015 2541 3049
rect 2580 3015 2609 3049
rect 2653 3015 2677 3049
rect 2726 3015 2745 3049
rect 2799 3015 2813 3049
rect 2872 3015 2881 3049
rect 2945 3015 2949 3049
rect 2983 3015 2984 3049
rect 3051 3015 3057 3049
rect 3119 3015 3130 3049
rect 3187 3015 3203 3049
rect 3255 3015 3276 3049
rect 3323 3015 3349 3049
rect 3391 3015 3422 3049
rect 3459 3015 3493 3049
rect 3529 3015 3561 3049
rect 3602 3015 3629 3049
rect 3663 3015 3678 3049
rect 3731 3015 3754 3049
rect 3799 3015 3831 3049
rect 3867 3015 3901 3049
rect 3942 3015 3969 3049
rect 4019 3015 4037 3049
rect 4096 3015 4105 3049
rect 4207 3015 4216 3049
rect 4275 3015 4293 3049
rect 4343 3015 4370 3049
rect 4411 3015 4445 3049
rect 4481 3015 4513 3049
rect 4558 3015 4581 3049
rect 4635 3015 4713 3049
rect 427 3009 4713 3015
rect 427 2977 473 3009
rect 427 2943 433 2977
rect 467 2943 473 2977
rect 427 2938 473 2943
rect 427 2904 433 2938
rect 467 2904 473 2938
rect 427 2902 473 2904
rect 427 2836 433 2902
rect 467 2836 473 2902
rect 4667 2981 4713 3009
rect 4667 2941 4673 2981
rect 4707 2941 4713 2981
rect 4667 2913 4713 2941
rect 4667 2867 4673 2913
rect 4707 2867 4713 2913
rect 427 2827 473 2836
rect 193 2783 244 2812
rect 193 2780 210 2783
rect -101 2764 -67 2776
rect -101 2692 -67 2726
rect -101 2624 -67 2650
rect -101 2556 -67 2570
rect -101 2488 -67 2489
rect -101 2442 -67 2454
rect -101 2361 -67 2386
rect -101 2284 -67 2318
rect -101 2234 -67 2246
rect 55 2764 89 2776
rect 55 2692 89 2726
rect 55 2624 89 2650
rect 55 2556 89 2570
rect 55 2488 89 2489
rect 55 2442 89 2454
rect 55 2361 89 2386
rect 55 2284 89 2318
rect 55 2234 89 2246
rect 193 2746 199 2780
rect 233 2746 244 2749
rect 193 2715 244 2746
rect 193 2705 210 2715
rect 193 2671 199 2705
rect 233 2671 244 2681
rect 193 2647 244 2671
rect 193 2630 210 2647
rect 193 2596 199 2630
rect 233 2596 244 2613
rect 193 2579 244 2596
rect 193 2555 210 2579
rect 193 2521 199 2555
rect 233 2521 244 2545
rect 193 2511 244 2521
rect 193 2480 210 2511
rect 193 2446 199 2480
rect 233 2446 244 2477
rect 193 2443 244 2446
rect 193 2409 210 2443
rect 193 2405 244 2409
rect 193 2371 199 2405
rect 233 2375 244 2405
rect 193 2341 210 2371
rect 193 2330 244 2341
rect 193 2296 199 2330
rect 233 2307 244 2330
rect 193 2273 210 2296
rect 193 2255 244 2273
rect 193 2221 199 2255
rect 233 2239 244 2255
rect 193 2205 210 2221
rect -71 2156 -59 2190
rect -21 2156 13 2190
rect 47 2156 63 2190
rect 193 2180 244 2205
rect 193 2146 199 2180
rect 233 2171 244 2180
rect 193 2137 210 2146
rect 193 2106 244 2137
rect 193 2072 199 2106
rect 233 2103 244 2106
rect 193 2069 210 2072
rect 193 2035 244 2069
rect 193 2032 210 2035
rect 193 1998 199 2032
rect 233 1998 244 2001
rect 193 1967 244 1998
rect 193 1958 210 1967
rect 193 1924 199 1958
rect 233 1924 244 1933
rect 193 1899 244 1924
rect 193 1865 210 1899
rect 427 2768 433 2827
rect 467 2768 473 2827
rect 427 2752 473 2768
rect 427 2700 433 2752
rect 467 2700 473 2752
rect 427 2677 473 2700
rect 427 2632 433 2677
rect 467 2632 473 2677
rect 427 2602 473 2632
rect 427 2564 433 2602
rect 467 2564 473 2602
rect 427 2530 473 2564
rect 427 2494 433 2530
rect 467 2494 473 2530
rect 427 2462 473 2494
rect 427 2420 433 2462
rect 467 2420 473 2462
rect 427 2394 473 2420
rect 427 2346 433 2394
rect 467 2346 473 2394
rect 427 2326 473 2346
rect 427 2272 433 2326
rect 467 2272 473 2326
rect 427 2258 473 2272
rect 427 2198 433 2258
rect 467 2198 473 2258
rect 427 2190 473 2198
rect 427 2124 433 2190
rect 467 2124 473 2190
rect 427 2122 473 2124
rect 427 2088 433 2122
rect 467 2088 473 2122
rect 427 2084 473 2088
rect 427 2020 433 2084
rect 467 2020 473 2084
rect 427 2010 473 2020
rect 427 1952 433 2010
rect 467 1952 473 2010
rect 427 1936 473 1952
rect 244 1865 250 1890
rect 193 1844 250 1865
rect 204 1831 250 1844
rect 204 1778 210 1831
rect 244 1778 250 1831
rect 204 1763 250 1778
rect 204 1701 210 1763
rect 244 1701 250 1763
rect 204 1695 250 1701
rect 204 1663 210 1695
rect 244 1663 250 1695
rect 427 1884 433 1936
rect 467 1884 473 1936
rect 720 2788 754 2817
rect 720 2715 754 2749
rect 720 2647 754 2675
rect 720 2579 754 2596
rect 720 2511 754 2517
rect 720 2472 754 2477
rect 720 2393 754 2409
rect 720 2314 754 2341
rect 720 2239 754 2273
rect 720 2171 754 2200
rect 720 2103 754 2120
rect 720 2035 754 2069
rect 720 1967 754 2001
rect 720 1917 754 1933
rect 876 2792 910 2817
rect 876 2717 910 2749
rect 876 2647 910 2681
rect 876 2579 910 2608
rect 876 2511 910 2533
rect 876 2443 910 2458
rect 876 2375 910 2383
rect 876 2307 910 2308
rect 876 2267 910 2273
rect 876 2192 910 2205
rect 876 2117 910 2137
rect 876 2042 910 2069
rect 876 1967 910 2001
rect 876 1917 910 1933
rect 1032 2792 1066 2817
rect 1032 2717 1066 2749
rect 1032 2647 1066 2681
rect 1032 2579 1066 2608
rect 1032 2511 1066 2533
rect 1032 2443 1066 2458
rect 1032 2375 1066 2383
rect 1032 2307 1066 2308
rect 1032 2267 1066 2273
rect 1032 2192 1066 2205
rect 1032 2117 1066 2137
rect 1032 2042 1066 2069
rect 1032 1967 1066 2001
rect 1032 1917 1066 1933
rect 1142 2792 1176 2817
rect 1142 2717 1176 2749
rect 1142 2647 1176 2681
rect 1142 2579 1176 2608
rect 1142 2511 1176 2533
rect 1142 2443 1176 2458
rect 1142 2375 1176 2383
rect 1142 2307 1176 2308
rect 1142 2267 1176 2273
rect 1142 2192 1176 2205
rect 1142 2117 1176 2137
rect 1142 2042 1176 2069
rect 1142 1967 1176 2001
rect 1142 1917 1176 1933
rect 1298 2792 1332 2817
rect 1298 2717 1332 2749
rect 1298 2647 1332 2681
rect 1298 2579 1332 2608
rect 1298 2511 1332 2533
rect 1298 2443 1332 2458
rect 1298 2375 1332 2383
rect 1298 2307 1332 2308
rect 1298 2267 1332 2273
rect 1298 2192 1332 2205
rect 1298 2117 1332 2137
rect 1298 2042 1332 2069
rect 1298 1967 1332 2001
rect 1298 1917 1332 1933
rect 1454 2788 1488 2817
rect 1454 2715 1488 2749
rect 1454 2647 1488 2675
rect 1454 2579 1488 2596
rect 1454 2511 1488 2517
rect 1454 2472 1488 2477
rect 1454 2393 1488 2409
rect 1454 2314 1488 2341
rect 1454 2239 1488 2273
rect 1454 2171 1488 2200
rect 1454 2103 1488 2120
rect 1454 2035 1488 2069
rect 1454 1967 1488 2001
rect 1454 1917 1488 1933
rect 1610 2792 1644 2817
rect 1610 2717 1644 2749
rect 1610 2647 1644 2681
rect 1610 2579 1644 2608
rect 1610 2511 1644 2533
rect 1610 2443 1644 2458
rect 1610 2375 1644 2383
rect 1610 2307 1644 2308
rect 1610 2267 1644 2273
rect 1610 2192 1644 2205
rect 1610 2117 1644 2137
rect 1610 2042 1644 2069
rect 1610 1967 1644 2001
rect 1610 1917 1644 1933
rect 1766 2788 1800 2817
rect 1766 2715 1800 2749
rect 1766 2647 1800 2675
rect 1766 2579 1800 2596
rect 1766 2511 1800 2517
rect 1766 2472 1800 2477
rect 1766 2393 1800 2409
rect 1766 2314 1800 2341
rect 1766 2239 1800 2273
rect 1766 2171 1800 2200
rect 1766 2103 1800 2120
rect 1766 2035 1800 2069
rect 1766 1967 1800 2001
rect 1766 1917 1800 1933
rect 1922 2792 1956 2817
rect 1922 2717 1956 2749
rect 1922 2647 1956 2681
rect 1922 2579 1956 2608
rect 1922 2511 1956 2533
rect 1922 2443 1956 2458
rect 1922 2375 1956 2383
rect 1922 2307 1956 2308
rect 1922 2267 1956 2273
rect 1922 2192 1956 2205
rect 1922 2117 1956 2137
rect 1922 2042 1956 2069
rect 1922 1967 1956 2001
rect 1922 1917 1956 1933
rect 2078 2792 2112 2817
rect 2078 2717 2112 2749
rect 2078 2647 2112 2681
rect 2078 2579 2112 2608
rect 2078 2511 2112 2533
rect 2078 2443 2112 2458
rect 2078 2375 2112 2383
rect 2078 2307 2112 2308
rect 2078 2267 2112 2273
rect 2078 2192 2112 2205
rect 2078 2117 2112 2137
rect 2078 2042 2112 2069
rect 2078 1967 2112 2001
rect 2078 1917 2112 1933
rect 2234 2792 2268 2817
rect 2234 2717 2268 2749
rect 2234 2647 2268 2681
rect 2234 2579 2268 2608
rect 2234 2511 2268 2533
rect 2234 2443 2268 2458
rect 2234 2375 2268 2383
rect 2234 2307 2268 2308
rect 2234 2267 2268 2273
rect 2234 2192 2268 2205
rect 2234 2117 2268 2137
rect 2234 2042 2268 2069
rect 2234 1967 2268 2001
rect 2234 1917 2268 1933
rect 2390 2792 2424 2817
rect 2390 2717 2424 2749
rect 2390 2647 2424 2681
rect 2390 2579 2424 2608
rect 2390 2511 2424 2533
rect 2390 2443 2424 2458
rect 2390 2375 2424 2383
rect 2390 2307 2424 2308
rect 2390 2267 2424 2273
rect 2390 2192 2424 2205
rect 2390 2117 2424 2137
rect 2390 2042 2424 2069
rect 2390 1967 2424 2001
rect 2390 1917 2424 1933
rect 2546 2792 2580 2817
rect 2546 2717 2580 2749
rect 2546 2647 2580 2681
rect 2546 2579 2580 2608
rect 2546 2511 2580 2533
rect 2546 2443 2580 2458
rect 2546 2375 2580 2383
rect 2546 2307 2580 2308
rect 2546 2267 2580 2273
rect 2546 2192 2580 2205
rect 2546 2117 2580 2137
rect 2546 2042 2580 2069
rect 2546 1967 2580 2001
rect 2546 1917 2580 1933
rect 2702 2792 2736 2817
rect 2702 2717 2736 2749
rect 2702 2647 2736 2681
rect 2702 2579 2736 2608
rect 2702 2511 2736 2533
rect 2702 2443 2736 2458
rect 2702 2375 2736 2383
rect 2702 2307 2736 2308
rect 2702 2267 2736 2273
rect 2702 2192 2736 2205
rect 2702 2117 2736 2137
rect 2702 2042 2736 2069
rect 2702 1967 2736 2001
rect 2702 1917 2736 1933
rect 2858 2792 2892 2817
rect 2858 2717 2892 2749
rect 2858 2647 2892 2681
rect 2858 2579 2892 2608
rect 2858 2511 2892 2533
rect 2858 2443 2892 2458
rect 2858 2375 2892 2383
rect 2858 2307 2892 2308
rect 2858 2267 2892 2273
rect 2858 2192 2892 2205
rect 2858 2117 2892 2137
rect 2858 2042 2892 2069
rect 2858 1967 2892 2001
rect 2858 1917 2892 1933
rect 3014 2792 3048 2817
rect 3014 2717 3048 2749
rect 3014 2647 3048 2681
rect 3014 2579 3048 2608
rect 3014 2511 3048 2533
rect 3014 2443 3048 2458
rect 3014 2375 3048 2383
rect 3014 2307 3048 2308
rect 3014 2267 3048 2273
rect 3014 2192 3048 2205
rect 3014 2117 3048 2137
rect 3014 2042 3048 2069
rect 3014 1967 3048 2001
rect 3014 1917 3048 1933
rect 3170 2792 3204 2817
rect 3170 2717 3204 2749
rect 3170 2647 3204 2681
rect 3170 2579 3204 2608
rect 3170 2511 3204 2533
rect 3170 2443 3204 2458
rect 3170 2375 3204 2383
rect 3170 2307 3204 2308
rect 3170 2267 3204 2273
rect 3170 2192 3204 2205
rect 3170 2117 3204 2137
rect 3170 2042 3204 2069
rect 3170 1967 3204 2001
rect 3170 1917 3204 1933
rect 3326 2792 3360 2817
rect 3326 2717 3360 2749
rect 3326 2647 3360 2681
rect 3326 2579 3360 2608
rect 3326 2511 3360 2533
rect 3326 2443 3360 2458
rect 3326 2375 3360 2383
rect 3326 2307 3360 2308
rect 3326 2267 3360 2273
rect 3326 2192 3360 2205
rect 3326 2117 3360 2137
rect 3326 2042 3360 2069
rect 3326 1967 3360 2001
rect 3326 1917 3360 1933
rect 3482 2792 3516 2817
rect 3482 2717 3516 2749
rect 3482 2647 3516 2681
rect 3482 2579 3516 2608
rect 3482 2511 3516 2533
rect 3482 2443 3516 2458
rect 3482 2375 3516 2383
rect 3482 2307 3516 2308
rect 3482 2267 3516 2273
rect 3482 2192 3516 2205
rect 3482 2117 3516 2137
rect 3482 2042 3516 2069
rect 3482 1967 3516 2001
rect 3482 1917 3516 1933
rect 3638 2789 3672 2817
rect 3638 2715 3672 2749
rect 3638 2647 3672 2677
rect 3638 2579 3672 2599
rect 3638 2511 3672 2520
rect 3638 2475 3672 2477
rect 3638 2396 3672 2409
rect 3638 2317 3672 2341
rect 3638 2239 3672 2273
rect 3638 2171 3672 2204
rect 3638 2103 3672 2125
rect 3638 2035 3672 2046
rect 3638 1967 3672 2001
rect 3638 1917 3672 1933
rect 3794 2792 3828 2817
rect 3794 2717 3828 2749
rect 3794 2647 3828 2681
rect 3794 2579 3828 2608
rect 3794 2511 3828 2533
rect 3794 2443 3828 2458
rect 3794 2375 3828 2383
rect 3794 2307 3828 2308
rect 3794 2267 3828 2273
rect 3794 2192 3828 2205
rect 3794 2117 3828 2137
rect 3794 2042 3828 2069
rect 3794 1967 3828 2001
rect 3794 1917 3828 1933
rect 3950 2790 3984 2817
rect 3950 2715 3984 2749
rect 3950 2647 3984 2678
rect 3950 2579 3984 2600
rect 3950 2511 3984 2522
rect 3950 2443 3984 2444
rect 3950 2400 3984 2409
rect 3950 2322 3984 2341
rect 3950 2244 3984 2273
rect 3950 2171 3984 2205
rect 3950 2103 3984 2132
rect 3950 2035 3984 2054
rect 3950 1967 3984 2001
rect 3950 1917 3984 1933
rect 4106 2792 4140 2817
rect 4106 2717 4140 2749
rect 4106 2647 4140 2681
rect 4106 2579 4140 2608
rect 4667 2845 4713 2867
rect 4667 2793 4673 2845
rect 4707 2793 4713 2845
rect 4667 2777 4713 2793
rect 4667 2719 4673 2777
rect 4707 2719 4713 2777
rect 4667 2709 4713 2719
rect 4667 2645 4673 2709
rect 4707 2645 4713 2709
rect 4667 2641 4713 2645
rect 4667 2607 4673 2641
rect 4707 2607 4713 2641
rect 4667 2605 4713 2607
rect 4261 2569 4277 2603
rect 4338 2569 4372 2603
rect 4422 2569 4467 2603
rect 4505 2569 4517 2603
rect 4106 2511 4140 2533
rect 4667 2539 4673 2605
rect 4707 2539 4713 2605
rect 4667 2531 4713 2539
rect 4667 2471 4673 2531
rect 4707 2471 4713 2531
rect 4106 2443 4140 2458
rect 4106 2375 4140 2383
rect 4106 2307 4140 2308
rect 4106 2267 4140 2273
rect 4106 2192 4140 2205
rect 4106 2117 4140 2137
rect 4106 2042 4140 2069
rect 4106 1967 4140 2001
rect 4106 1917 4140 1933
rect 4216 2377 4250 2409
rect 4216 2307 4250 2341
rect 4216 2239 4250 2261
rect 4216 2171 4250 2179
rect 4216 2131 4250 2137
rect 4216 2049 4250 2069
rect 4216 1967 4250 2001
rect 4216 1917 4250 1933
rect 4372 2377 4406 2409
rect 4372 2307 4406 2341
rect 4372 2239 4406 2261
rect 4372 2171 4406 2179
rect 4372 2131 4406 2137
rect 4372 2049 4406 2069
rect 4372 1967 4406 2001
rect 4372 1917 4406 1933
rect 4528 2377 4562 2409
rect 4528 2307 4562 2341
rect 4528 2239 4562 2261
rect 4528 2171 4562 2179
rect 4528 2131 4562 2137
rect 4528 2049 4562 2069
rect 4528 1967 4562 2001
rect 4528 1917 4562 1933
rect 4667 2457 4713 2471
rect 4667 2403 4673 2457
rect 4707 2403 4713 2457
rect 4667 2383 4713 2403
rect 4667 2335 4673 2383
rect 4707 2335 4713 2383
rect 4667 2309 4713 2335
rect 4667 2267 4673 2309
rect 4707 2267 4713 2309
rect 4667 2235 4713 2267
rect 4667 2199 4673 2235
rect 4707 2199 4713 2235
rect 4667 2165 4713 2199
rect 4667 2127 4673 2165
rect 4707 2127 4713 2165
rect 4667 2097 4713 2127
rect 4667 2052 4673 2097
rect 4707 2052 4713 2097
rect 4667 2029 4713 2052
rect 4667 1977 4673 2029
rect 4707 1977 4713 2029
rect 4667 1961 4713 1977
rect 427 1862 473 1884
rect 4667 1902 4673 1961
rect 4707 1902 4713 1961
rect 4667 1893 4713 1902
rect 427 1816 433 1862
rect 467 1816 473 1862
rect 751 1839 781 1873
rect 815 1839 817 1873
rect 851 1839 876 1873
rect 910 1839 917 1873
rect 951 1839 971 1873
rect 1005 1839 1021 1873
rect 1187 1839 1203 1873
rect 1237 1839 1245 1873
rect 1311 1839 1318 1873
rect 1385 1839 1391 1873
rect 1459 1839 1464 1873
rect 1498 1839 1499 1873
rect 1533 1839 1537 1873
rect 1571 1839 1573 1873
rect 1607 1839 1610 1873
rect 1644 1839 1647 1873
rect 1681 1839 1682 1873
rect 1716 1839 1721 1873
rect 1788 1839 1795 1873
rect 1860 1839 1869 1873
rect 1932 1839 1943 1873
rect 2004 1839 2017 1873
rect 2051 1839 2067 1873
rect 2123 1839 2139 1873
rect 2200 1839 2210 1873
rect 2273 1839 2281 1873
rect 2346 1839 2353 1873
rect 2419 1839 2425 1873
rect 2491 1839 2497 1873
rect 2563 1839 2569 1873
rect 2603 1839 2641 1873
rect 2675 1839 2691 1873
rect 2747 1839 2762 1873
rect 2797 1839 2835 1873
rect 2879 1839 2907 1873
rect 2962 1839 2979 1873
rect 3045 1839 3051 1873
rect 3085 1839 3094 1873
rect 3157 1839 3176 1873
rect 3228 1839 3258 1873
rect 3299 1839 3315 1873
rect 3371 1839 3387 1873
rect 3421 1839 3461 1873
rect 3495 1839 3534 1873
rect 3568 1839 3607 1873
rect 3641 1839 3661 1873
rect 3714 1839 3734 1873
rect 3787 1839 3807 1873
rect 3860 1839 3880 1873
rect 3933 1839 3953 1873
rect 4006 1839 4025 1873
rect 4079 1839 4095 1873
rect 427 1788 473 1816
rect 427 1748 433 1788
rect 467 1748 473 1788
rect 427 1720 473 1748
rect 4667 1827 4673 1893
rect 4707 1827 4713 1893
rect 4667 1788 4713 1827
rect 4667 1752 4673 1788
rect 4707 1752 4713 1788
rect 4667 1720 4713 1752
rect 427 1714 516 1720
rect 1029 1714 2207 1720
rect 2358 1714 3506 1720
rect 4135 1714 4713 1720
rect 427 1680 525 1714
rect 559 1680 593 1714
rect 627 1680 661 1714
rect 695 1680 729 1714
rect 763 1680 797 1714
rect 831 1680 865 1714
rect 899 1680 933 1714
rect 967 1680 1001 1714
rect 1035 1680 1067 1714
rect 1103 1680 1137 1714
rect 1178 1680 1205 1714
rect 1255 1680 1273 1714
rect 1332 1680 1341 1714
rect 1443 1680 1451 1714
rect 1511 1680 1527 1714
rect 1579 1680 1603 1714
rect 1647 1680 1679 1714
rect 1715 1680 1749 1714
rect 1789 1680 1817 1714
rect 1865 1680 1885 1714
rect 1941 1680 1953 1714
rect 2017 1680 2021 1714
rect 2055 1680 2059 1714
rect 2123 1680 2135 1714
rect 2191 1680 2225 1714
rect 2259 1680 2293 1714
rect 2327 1680 2361 1714
rect 2395 1680 2396 1714
rect 2463 1680 2476 1714
rect 2531 1680 2556 1714
rect 2599 1680 2633 1714
rect 2670 1680 2701 1714
rect 2750 1680 2769 1714
rect 2829 1680 2837 1714
rect 2871 1680 2874 1714
rect 2939 1680 2973 1714
rect 3018 1680 3041 1714
rect 3093 1680 3109 1714
rect 3168 1680 3177 1714
rect 3243 1680 3245 1714
rect 3279 1680 3284 1714
rect 3347 1680 3359 1714
rect 3415 1680 3434 1714
rect 3483 1680 3517 1714
rect 3551 1680 3585 1714
rect 3619 1680 3653 1714
rect 3687 1680 3721 1714
rect 3755 1680 3789 1714
rect 3823 1680 3857 1714
rect 3891 1680 3925 1714
rect 3959 1680 3993 1714
rect 4027 1680 4061 1714
rect 4095 1680 4129 1714
rect 4163 1680 4173 1714
rect 4231 1680 4257 1714
rect 4299 1680 4333 1714
rect 4375 1680 4401 1714
rect 4458 1680 4469 1714
rect 4503 1680 4507 1714
rect 4571 1680 4590 1714
rect 4639 1680 4713 1714
rect 427 1674 516 1680
rect 1029 1674 2207 1680
rect 2358 1674 3506 1680
rect 4135 1674 4713 1680
rect 4890 3016 4896 3068
rect 4930 3016 4936 3068
rect 4890 3000 4936 3016
rect 4890 2942 4896 3000
rect 4930 2942 4936 3000
rect 4890 2932 4936 2942
rect 4890 2868 4896 2932
rect 4930 2868 4936 2932
rect 4890 2864 4936 2868
rect 4890 2830 4896 2864
rect 4930 2830 4936 2864
rect 4890 2828 4936 2830
rect 4890 2762 4896 2828
rect 4930 2762 4936 2828
rect 4890 2754 4936 2762
rect 4890 2694 4896 2754
rect 4930 2694 4936 2754
rect 4890 2680 4936 2694
rect 4890 2626 4896 2680
rect 4930 2626 4936 2680
rect 4890 2606 4936 2626
rect 4890 2558 4896 2606
rect 4930 2558 4936 2606
rect 4890 2532 4936 2558
rect 4890 2490 4896 2532
rect 4930 2490 4936 2532
rect 4890 2458 4936 2490
rect 4890 2422 4896 2458
rect 4930 2422 4936 2458
rect 4890 2388 4936 2422
rect 4890 2350 4896 2388
rect 4930 2350 4936 2388
rect 4890 2320 4936 2350
rect 4890 2276 4896 2320
rect 4930 2276 4936 2320
rect 4890 2252 4936 2276
rect 4890 2202 4896 2252
rect 4930 2202 4936 2252
rect 4890 2184 4936 2202
rect 4890 2127 4896 2184
rect 4930 2127 4936 2184
rect 4890 2116 4936 2127
rect 4890 2052 4896 2116
rect 4930 2052 4936 2116
rect 4890 2048 4936 2052
rect 4890 2014 4896 2048
rect 4930 2014 4936 2048
rect 4890 2011 4936 2014
rect 4890 1946 4896 2011
rect 4930 1946 4936 2011
rect 4890 1936 4936 1946
rect 4890 1878 4896 1936
rect 4930 1878 4936 1936
rect 4890 1861 4936 1878
rect 4890 1810 4896 1861
rect 4930 1810 4936 1861
rect 4890 1786 4936 1810
rect 4890 1742 4896 1786
rect 4930 1742 4936 1786
rect 4890 1711 4936 1742
rect 4890 1674 4896 1711
rect 4930 1674 4936 1711
rect 210 1627 244 1661
rect 210 1559 244 1593
rect 210 1495 244 1525
rect 4890 1640 4936 1674
rect 4890 1602 4896 1640
rect 4930 1602 4936 1640
rect 4890 1561 4936 1602
rect 4890 1527 4896 1561
rect 4930 1527 4936 1561
rect 4890 1495 4936 1527
rect 210 1491 4936 1495
rect 210 1457 340 1491
rect 374 1457 408 1491
rect 442 1457 476 1491
rect 510 1457 544 1491
rect 578 1457 612 1491
rect 646 1457 680 1491
rect 714 1457 748 1491
rect 782 1457 816 1491
rect 850 1457 884 1491
rect 918 1457 952 1491
rect 986 1490 1020 1491
rect 1054 1490 1088 1491
rect 1122 1490 1156 1491
rect 1190 1490 1224 1491
rect 1258 1490 1292 1491
rect 991 1457 1020 1490
rect 1065 1457 1088 1490
rect 1139 1457 1156 1490
rect 1213 1457 1224 1490
rect 1287 1457 1292 1490
rect 1326 1490 1360 1491
rect 1394 1490 1428 1491
rect 1462 1490 1496 1491
rect 1530 1490 1564 1491
rect 1598 1490 1632 1491
rect 1666 1490 1700 1491
rect 1326 1457 1327 1490
rect 1394 1457 1401 1490
rect 1462 1457 1475 1490
rect 1530 1457 1549 1490
rect 1598 1457 1623 1490
rect 1666 1457 1697 1490
rect 1734 1457 1768 1491
rect 1802 1490 1836 1491
rect 1870 1490 1904 1491
rect 1938 1490 1972 1491
rect 2006 1490 2040 1491
rect 2074 1490 2108 1491
rect 1805 1457 1836 1490
rect 1879 1457 1904 1490
rect 1953 1457 1972 1490
rect 2027 1457 2040 1490
rect 2102 1457 2108 1490
rect 2142 1490 2176 1491
rect 2142 1457 2143 1490
rect 2210 1457 2244 1491
rect 2278 1457 2312 1491
rect 2346 1490 2380 1491
rect 2346 1457 2375 1490
rect 2414 1457 2448 1491
rect 2482 1490 2516 1491
rect 2550 1490 2584 1491
rect 2618 1490 2652 1491
rect 2686 1490 2720 1491
rect 2754 1490 2788 1491
rect 2822 1490 2856 1491
rect 2483 1457 2516 1490
rect 2557 1457 2584 1490
rect 2631 1457 2652 1490
rect 2705 1457 2720 1490
rect 2779 1457 2788 1490
rect 2853 1457 2856 1490
rect 2890 1490 2924 1491
rect 2958 1490 2992 1491
rect 3026 1490 3060 1491
rect 3094 1490 3128 1491
rect 3162 1490 3196 1491
rect 2890 1457 2893 1490
rect 2958 1457 2967 1490
rect 3026 1457 3041 1490
rect 3094 1457 3115 1490
rect 3162 1457 3190 1490
rect 3230 1457 3264 1491
rect 3298 1490 3332 1491
rect 3366 1490 3400 1491
rect 3434 1490 3468 1491
rect 3502 1490 3536 1491
rect 3570 1490 3604 1491
rect 3299 1457 3332 1490
rect 3374 1457 3400 1490
rect 3449 1457 3468 1490
rect 3524 1457 3536 1490
rect 3599 1457 3604 1490
rect 3638 1490 3672 1491
rect 3706 1490 3740 1491
rect 3774 1490 3808 1491
rect 3842 1490 3876 1491
rect 3638 1457 3640 1490
rect 3706 1457 3715 1490
rect 3774 1457 3790 1490
rect 3842 1457 3865 1490
rect 3910 1457 3944 1491
rect 3978 1457 4012 1491
rect 4046 1457 4080 1491
rect 4114 1489 4148 1491
rect 4146 1457 4148 1489
rect 4182 1489 4216 1491
rect 4250 1489 4284 1491
rect 4318 1489 4352 1491
rect 4182 1457 4191 1489
rect 4250 1457 4270 1489
rect 4318 1457 4349 1489
rect 4386 1457 4420 1491
rect 4454 1489 4488 1491
rect 4522 1489 4556 1491
rect 4590 1489 4624 1491
rect 4462 1457 4488 1489
rect 4540 1457 4556 1489
rect 4618 1457 4624 1489
rect 4658 1489 4692 1491
rect 4726 1489 4760 1491
rect 4794 1489 4828 1491
rect 4658 1457 4662 1489
rect 4726 1457 4740 1489
rect 4794 1457 4818 1489
rect 4862 1457 4936 1491
rect 210 1456 957 1457
rect 991 1456 1031 1457
rect 1065 1456 1105 1457
rect 1139 1456 1179 1457
rect 1213 1456 1253 1457
rect 1287 1456 1327 1457
rect 1361 1456 1401 1457
rect 1435 1456 1475 1457
rect 1509 1456 1549 1457
rect 1583 1456 1623 1457
rect 1657 1456 1697 1457
rect 1731 1456 1771 1457
rect 1805 1456 1845 1457
rect 1879 1456 1919 1457
rect 1953 1456 1993 1457
rect 2027 1456 2068 1457
rect 2102 1456 2143 1457
rect 2177 1456 2375 1457
rect 2409 1456 2449 1457
rect 2483 1456 2523 1457
rect 2557 1456 2597 1457
rect 2631 1456 2671 1457
rect 2705 1456 2745 1457
rect 2779 1456 2819 1457
rect 2853 1456 2893 1457
rect 2927 1456 2967 1457
rect 3001 1456 3041 1457
rect 3075 1456 3115 1457
rect 3149 1456 3190 1457
rect 3224 1456 3265 1457
rect 3299 1456 3340 1457
rect 3374 1456 3415 1457
rect 3449 1456 3490 1457
rect 3524 1456 3565 1457
rect 3599 1456 3640 1457
rect 3674 1456 3715 1457
rect 3749 1456 3790 1457
rect 3824 1456 3865 1457
rect 3899 1456 4112 1457
rect 210 1455 4112 1456
rect 4146 1455 4191 1457
rect 4225 1455 4270 1457
rect 4304 1455 4349 1457
rect 4383 1455 4428 1457
rect 4462 1455 4506 1457
rect 4540 1455 4584 1457
rect 4618 1455 4662 1457
rect 4696 1455 4740 1457
rect 4774 1455 4818 1457
rect 4852 1455 4936 1457
rect 210 1449 4936 1455
rect 5098 3238 5170 3272
rect 5211 3238 5245 3272
rect 5279 3238 5313 3272
rect 5354 3238 5381 3272
rect 5429 3238 5449 3272
rect 5504 3238 5517 3272
rect 5579 3238 5585 3272
rect 5687 3238 5693 3272
rect 5755 3238 5767 3272
rect 5823 3238 5841 3272
rect 5891 3238 5915 3272
rect 5959 3238 5989 3272
rect 6027 3238 6061 3272
rect 6097 3238 6129 3272
rect 6171 3238 6197 3272
rect 6245 3238 6265 3272
rect 6319 3238 6333 3272
rect 6393 3238 6401 3272
rect 6467 3238 6469 3272
rect 6503 3238 6507 3272
rect 6571 3238 6581 3272
rect 6639 3238 6655 3272
rect 6707 3238 6729 3272
rect 6775 3238 6803 3272
rect 6843 3238 6911 3272
rect 5098 3204 5133 3238
rect 5098 3198 5099 3204
rect 5132 3164 5133 3170
rect 5098 3136 5133 3164
rect 5098 3124 5099 3136
rect 5132 3090 5133 3102
rect 5098 3068 5133 3090
rect 5098 3050 5099 3068
rect 6877 3200 6911 3238
rect 6877 3126 6911 3157
rect 6877 3055 6911 3089
rect 5132 3016 5133 3034
rect 5098 3000 5133 3016
rect 5098 2976 5099 3000
rect 5132 2942 5133 2966
rect 5098 2932 5133 2942
rect 5098 2902 5099 2932
rect 5132 2868 5133 2898
rect 5098 2864 5133 2868
rect 5098 2830 5099 2864
rect 5098 2828 5133 2830
rect 5132 2796 5133 2828
rect 5098 2762 5099 2794
rect 5098 2754 5133 2762
rect 5132 2728 5133 2754
rect 5098 2694 5099 2720
rect 5098 2680 5133 2694
rect 5132 2660 5133 2680
rect 5098 2626 5099 2646
rect 5098 2606 5133 2626
rect 5132 2592 5133 2606
rect 5098 2558 5099 2572
rect 5098 2532 5133 2558
rect 5132 2524 5133 2532
rect 5098 2490 5099 2498
rect 5098 2458 5133 2490
rect 5132 2456 5133 2458
rect 5098 2422 5099 2424
rect 5098 2388 5133 2422
rect 5098 2384 5099 2388
rect 5132 2350 5133 2354
rect 5098 2320 5133 2350
rect 5098 2310 5099 2320
rect 5132 2276 5133 2286
rect 5098 2252 5133 2276
rect 5098 2236 5099 2252
rect 5132 2202 5133 2218
rect 5098 2184 5133 2202
rect 5098 2162 5099 2184
rect 5132 2128 5133 2150
rect 5098 2116 5133 2128
rect 5098 2088 5099 2116
rect 5132 2054 5133 2082
rect 5098 2048 5133 2054
rect 5098 2014 5099 2048
rect 5098 2013 5133 2014
rect 5132 1980 5133 2013
rect 5098 1946 5099 1979
rect 5098 1938 5133 1946
rect 5132 1912 5133 1938
rect 5098 1878 5099 1904
rect 5098 1863 5133 1878
rect 5132 1844 5133 1863
rect 5098 1810 5099 1829
rect 5098 1788 5133 1810
rect 5132 1776 5133 1788
rect 5098 1742 5099 1754
rect 5098 1713 5133 1742
rect 5132 1708 5133 1713
rect 5098 1674 5099 1679
rect 5351 3049 6697 3055
rect 5351 3015 5433 3049
rect 5477 3015 5501 3049
rect 5564 3015 5569 3049
rect 5603 3015 5637 3049
rect 5674 3015 5705 3049
rect 5746 3015 5773 3049
rect 5818 3015 5841 3049
rect 5890 3015 5909 3049
rect 5962 3015 5977 3049
rect 6035 3015 6045 3049
rect 6108 3015 6113 3049
rect 6215 3015 6220 3049
rect 6283 3015 6293 3049
rect 6351 3015 6366 3049
rect 6419 3015 6439 3049
rect 6487 3015 6512 3049
rect 6555 3015 6585 3049
rect 6623 3015 6697 3049
rect 5351 3009 6697 3015
rect 5351 2981 5397 3009
rect 5351 2943 5357 2981
rect 5391 2943 5397 2981
rect 5351 2913 5397 2943
rect 5351 2868 5357 2913
rect 5391 2868 5397 2913
rect 5351 2845 5397 2868
rect 6651 2975 6697 3009
rect 6651 2941 6657 2975
rect 6691 2941 6697 2975
rect 6651 2938 6697 2941
rect 6651 2904 6657 2938
rect 6691 2904 6697 2938
rect 6651 2901 6697 2904
rect 5351 2793 5357 2845
rect 5391 2793 5397 2845
rect 5351 2777 5397 2793
rect 5351 2718 5357 2777
rect 5391 2718 5397 2777
rect 5351 2709 5397 2718
rect 5351 2643 5357 2709
rect 5391 2643 5397 2709
rect 5351 2641 5397 2643
rect 5351 2607 5357 2641
rect 5391 2607 5397 2641
rect 5351 2602 5397 2607
rect 5351 2539 5357 2602
rect 5391 2539 5397 2602
rect 5351 2528 5397 2539
rect 5351 2471 5357 2528
rect 5391 2471 5397 2528
rect 5351 2454 5397 2471
rect 5351 2403 5357 2454
rect 5391 2403 5397 2454
rect 5351 2380 5397 2403
rect 5351 2335 5357 2380
rect 5391 2335 5397 2380
rect 5351 2306 5397 2335
rect 5351 2267 5357 2306
rect 5391 2267 5397 2306
rect 5351 2233 5397 2267
rect 5351 2198 5357 2233
rect 5391 2198 5397 2233
rect 5351 2165 5397 2198
rect 5351 2124 5357 2165
rect 5391 2124 5397 2165
rect 5351 2097 5397 2124
rect 5351 2050 5357 2097
rect 5391 2050 5397 2097
rect 5351 2029 5397 2050
rect 5351 1976 5357 2029
rect 5391 1976 5397 2029
rect 5351 1961 5397 1976
rect 5351 1902 5357 1961
rect 5391 1902 5397 1961
rect 5502 2792 5536 2817
rect 5502 2717 5536 2749
rect 5502 2647 5536 2681
rect 5502 2579 5536 2608
rect 5502 2511 5536 2533
rect 5502 2443 5536 2458
rect 5502 2375 5536 2383
rect 5502 2307 5536 2308
rect 5502 2267 5536 2273
rect 5502 2192 5536 2205
rect 5502 2117 5536 2137
rect 5502 2042 5536 2069
rect 5502 1967 5536 2001
rect 5502 1917 5536 1933
rect 5658 2788 5692 2817
rect 5658 2715 5692 2749
rect 5658 2647 5692 2675
rect 5658 2579 5692 2596
rect 5658 2511 5692 2517
rect 5658 2472 5692 2477
rect 5658 2393 5692 2409
rect 5658 2314 5692 2341
rect 5658 2239 5692 2273
rect 5658 2171 5692 2200
rect 5658 2103 5692 2120
rect 5658 2035 5692 2069
rect 5658 1967 5692 2001
rect 5846 2851 5848 2867
rect 5812 2817 5814 2833
rect 5812 2792 5848 2817
rect 5846 2783 5848 2792
rect 5812 2749 5814 2758
rect 5812 2717 5848 2749
rect 5846 2715 5848 2717
rect 5812 2681 5814 2683
rect 5812 2647 5848 2681
rect 5812 2642 5814 2647
rect 5846 2608 5848 2613
rect 5812 2579 5848 2608
rect 5812 2567 5814 2579
rect 5846 2533 5848 2545
rect 5812 2511 5848 2533
rect 5812 2492 5814 2511
rect 5846 2458 5848 2477
rect 5812 2443 5848 2458
rect 5812 2417 5814 2443
rect 5846 2383 5848 2409
rect 5812 2375 5848 2383
rect 5812 2342 5814 2375
rect 5846 2308 5848 2341
rect 5812 2307 5848 2308
rect 5812 2273 5814 2307
rect 5812 2267 5848 2273
rect 5846 2239 5848 2267
rect 5812 2205 5814 2233
rect 5812 2192 5848 2205
rect 5846 2171 5848 2192
rect 5812 2137 5814 2158
rect 5812 2117 5848 2137
rect 5846 2103 5848 2117
rect 5812 2069 5814 2083
rect 5812 2042 5848 2069
rect 5846 2035 5848 2042
rect 5812 2001 5814 2008
rect 5812 1967 5848 2001
rect 5658 1917 5692 1933
rect 5814 1917 5848 1933
rect 6030 2792 6064 2817
rect 6030 2717 6064 2749
rect 6030 2647 6064 2681
rect 6030 2579 6064 2608
rect 6030 2511 6064 2533
rect 6030 2443 6064 2458
rect 6030 2375 6064 2383
rect 6030 2307 6064 2308
rect 6030 2267 6064 2273
rect 6030 2192 6064 2205
rect 6030 2117 6064 2137
rect 6030 2042 6064 2069
rect 6030 1967 6064 2001
rect 6030 1917 6064 1933
rect 6246 2792 6280 2817
rect 6246 2717 6280 2749
rect 6246 2647 6280 2681
rect 6246 2579 6280 2608
rect 6246 2511 6280 2533
rect 6512 2788 6546 2833
rect 6512 2709 6546 2754
rect 6512 2629 6546 2675
rect 6512 2549 6546 2595
rect 6246 2443 6280 2458
rect 6246 2375 6280 2383
rect 6356 2509 6390 2519
rect 6356 2435 6390 2469
rect 6356 2389 6390 2401
rect 6356 2317 6390 2333
rect 6512 2503 6546 2515
rect 6512 2389 6546 2401
rect 6512 2317 6546 2333
rect 6651 2836 6657 2901
rect 6691 2836 6697 2901
rect 6651 2827 6697 2836
rect 6651 2768 6657 2827
rect 6691 2768 6697 2827
rect 6651 2753 6697 2768
rect 6651 2700 6657 2753
rect 6691 2700 6697 2753
rect 6651 2679 6697 2700
rect 6651 2632 6657 2679
rect 6691 2632 6697 2679
rect 6651 2605 6697 2632
rect 6651 2564 6657 2605
rect 6691 2564 6697 2605
rect 6651 2531 6697 2564
rect 6651 2496 6657 2531
rect 6691 2496 6697 2531
rect 6651 2462 6697 2496
rect 6651 2423 6657 2462
rect 6691 2423 6697 2462
rect 6651 2394 6697 2423
rect 6651 2349 6657 2394
rect 6691 2349 6697 2394
rect 6651 2326 6697 2349
rect 6246 2307 6280 2308
rect 6651 2275 6657 2326
rect 6691 2275 6697 2326
rect 6246 2267 6280 2273
rect 6401 2239 6417 2273
rect 6470 2239 6485 2273
rect 6651 2258 6697 2275
rect 6246 2192 6280 2205
rect 6246 2117 6280 2137
rect 6246 2042 6280 2069
rect 6246 1967 6280 2001
rect 6246 1917 6280 1933
rect 6651 2201 6657 2258
rect 6691 2201 6697 2258
rect 6651 2190 6697 2201
rect 6651 2127 6657 2190
rect 6691 2127 6697 2190
rect 6651 2122 6697 2127
rect 6651 2088 6657 2122
rect 6691 2088 6697 2122
rect 6651 2086 6697 2088
rect 6651 2020 6657 2086
rect 6691 2020 6697 2086
rect 6651 2011 6697 2020
rect 6651 1952 6657 2011
rect 6691 1952 6697 2011
rect 6651 1936 6697 1952
rect 5351 1893 5397 1902
rect 5351 1828 5357 1893
rect 5391 1828 5397 1893
rect 6651 1884 6657 1936
rect 6691 1884 6697 1936
rect 5547 1839 5563 1873
rect 5597 1839 5648 1873
rect 5692 1839 5733 1873
rect 5787 1839 5803 1873
rect 5859 1839 5875 1873
rect 5913 1839 5953 1873
rect 5990 1839 6031 1873
rect 6067 1839 6108 1873
rect 6144 1839 6185 1873
rect 6220 1839 6235 1873
rect 6651 1861 6697 1884
rect 5351 1788 5397 1828
rect 5351 1754 5357 1788
rect 5391 1754 5397 1788
rect 5351 1720 5397 1754
rect 6651 1816 6657 1861
rect 6691 1816 6697 1861
rect 6651 1786 6697 1816
rect 6651 1748 6657 1786
rect 6691 1748 6697 1786
rect 6651 1720 6697 1748
rect 5351 1714 5826 1720
rect 6509 1714 6697 1720
rect 5351 1680 5425 1714
rect 5463 1680 5493 1714
rect 5545 1680 5561 1714
rect 5626 1680 5629 1714
rect 5663 1680 5673 1714
rect 5731 1680 5754 1714
rect 5799 1680 5833 1714
rect 5867 1680 5901 1714
rect 5935 1680 5969 1714
rect 6003 1680 6037 1714
rect 6071 1680 6105 1714
rect 6139 1680 6173 1714
rect 6207 1680 6241 1714
rect 6275 1680 6309 1714
rect 6343 1680 6377 1714
rect 6411 1680 6445 1714
rect 6479 1680 6513 1714
rect 6547 1680 6566 1714
rect 6615 1680 6697 1714
rect 5351 1674 5826 1680
rect 6509 1674 6697 1680
rect 6877 2987 6911 3018
rect 6877 2919 6911 2944
rect 6877 2851 6911 2870
rect 6877 2783 6911 2796
rect 6877 2715 6911 2723
rect 6877 2647 6911 2650
rect 6877 2611 6911 2613
rect 6877 2538 6911 2545
rect 6877 2465 6911 2477
rect 6877 2392 6911 2409
rect 6877 2319 6911 2341
rect 6877 2246 6911 2273
rect 6877 2173 6911 2205
rect 6877 2103 6911 2137
rect 6877 2035 6911 2066
rect 6877 1967 6911 1993
rect 6877 1899 6911 1920
rect 6877 1831 6911 1847
rect 6877 1763 6911 1774
rect 6877 1695 6911 1701
rect 5098 1640 5133 1674
rect 5098 1638 5099 1640
rect 5132 1604 5133 1606
rect 5098 1563 5133 1604
rect 5132 1529 5133 1563
rect 5098 1491 5133 1529
rect 6877 1627 6911 1628
rect 6877 1589 6911 1593
rect 6877 1492 6911 1525
rect 6163 1491 6241 1492
rect 6275 1491 6319 1492
rect 6353 1491 6397 1492
rect 6431 1491 6476 1492
rect 6510 1491 6555 1492
rect 6589 1491 6634 1492
rect 6668 1491 6713 1492
rect 6747 1491 6792 1492
rect 6826 1491 6871 1492
rect 5098 1457 5167 1491
rect 5204 1457 5235 1491
rect 5276 1457 5303 1491
rect 5348 1457 5371 1491
rect 5420 1457 5439 1491
rect 5492 1457 5507 1491
rect 5564 1457 5575 1491
rect 5636 1457 5643 1491
rect 5709 1457 5711 1491
rect 5745 1457 5748 1491
rect 5813 1457 5847 1491
rect 5881 1457 5915 1491
rect 5949 1457 5983 1491
rect 6017 1457 6051 1491
rect 6085 1457 6119 1491
rect 6153 1457 6187 1491
rect 6221 1458 6241 1491
rect 6289 1458 6319 1491
rect 6221 1457 6255 1458
rect 6289 1457 6323 1458
rect 6357 1457 6391 1491
rect 6431 1458 6459 1491
rect 6510 1458 6527 1491
rect 6589 1458 6595 1491
rect 6425 1457 6459 1458
rect 6493 1457 6527 1458
rect 6561 1457 6595 1458
rect 6629 1458 6634 1491
rect 6697 1458 6713 1491
rect 6765 1458 6792 1491
rect 6833 1458 6871 1491
rect 6905 1491 6911 1492
rect 6993 3238 7077 3272
rect 7111 3238 7114 3272
rect 7148 3238 7155 3272
rect 7216 3238 7233 3272
rect 7284 3238 7311 3272
rect 7352 3238 7386 3272
rect 7424 3238 7454 3272
rect 7503 3238 7522 3272
rect 7582 3238 7590 3272
rect 7624 3238 7627 3272
rect 7692 3238 7726 3272
rect 7771 3238 7794 3272
rect 7846 3238 7862 3272
rect 7921 3238 7930 3272
rect 7996 3238 7998 3272
rect 8032 3238 8037 3272
rect 8100 3238 8112 3272
rect 8168 3238 8187 3272
rect 8236 3238 8262 3272
rect 8304 3238 8338 3272
rect 8372 3238 8406 3272
rect 8448 3238 8474 3272
rect 8524 3238 8542 3272
rect 8600 3238 8610 3272
rect 8676 3238 8678 3272
rect 8712 3238 8718 3272
rect 8780 3238 8794 3272
rect 8848 3238 8870 3272
rect 8916 3238 8946 3272
rect 8984 3238 9058 3272
rect 6993 3232 9058 3238
rect 6993 3204 7039 3232
rect 6993 3166 6999 3204
rect 7033 3166 7039 3204
rect 6993 3136 7039 3166
rect 6993 3093 6999 3136
rect 7033 3093 7039 3136
rect 6993 3068 7039 3093
rect 6993 3020 6999 3068
rect 7033 3020 7039 3068
rect 9012 3198 9058 3232
rect 9012 3157 9018 3198
rect 9052 3157 9058 3198
rect 9012 3124 9058 3157
rect 9012 3089 9018 3124
rect 9052 3089 9058 3124
rect 9012 3055 9058 3089
rect 6993 3000 7039 3020
rect 6993 2947 6999 3000
rect 7033 2947 7039 3000
rect 6993 2932 7039 2947
rect 6993 2874 6999 2932
rect 7033 2874 7039 2932
rect 6993 2864 7039 2874
rect 6993 2801 6999 2864
rect 7033 2801 7039 2864
rect 6993 2796 7039 2801
rect 6993 2694 6999 2796
rect 7033 2694 7039 2796
rect 6993 2689 7039 2694
rect 6993 2626 6999 2689
rect 7033 2626 7039 2689
rect 6993 2616 7039 2626
rect 6993 2558 6999 2616
rect 7033 2558 7039 2616
rect 6993 2543 7039 2558
rect 6993 2490 6999 2543
rect 7033 2490 7039 2543
rect 6993 2470 7039 2490
rect 6993 2422 6999 2470
rect 7033 2422 7039 2470
rect 6993 2397 7039 2422
rect 6993 2354 6999 2397
rect 7033 2354 7039 2397
rect 6993 2324 7039 2354
rect 6993 2286 6999 2324
rect 7033 2286 7039 2324
rect 6993 2252 7039 2286
rect 6993 2217 6999 2252
rect 7033 2217 7039 2252
rect 6993 2184 7039 2217
rect 6993 2144 6999 2184
rect 7033 2144 7039 2184
rect 6993 2116 7039 2144
rect 6993 2071 6999 2116
rect 7033 2071 7039 2116
rect 6993 2048 7039 2071
rect 6993 1998 6999 2048
rect 7033 1998 7039 2048
rect 6993 1980 7039 1998
rect 6993 1926 6999 1980
rect 7033 1926 7039 1980
rect 6993 1912 7039 1926
rect 6993 1854 6999 1912
rect 7033 1854 7039 1912
rect 6993 1844 7039 1854
rect 6993 1782 6999 1844
rect 7033 1782 7039 1844
rect 6993 1776 7039 1782
rect 6993 1710 6999 1776
rect 7033 1710 7039 1776
rect 6993 1708 7039 1710
rect 6993 1674 6999 1708
rect 7033 1674 7039 1708
rect 7219 3049 8835 3055
rect 7219 3015 7299 3049
rect 7336 3015 7367 3049
rect 7414 3015 7435 3049
rect 7492 3015 7503 3049
rect 7570 3015 7571 3049
rect 7605 3015 7639 3049
rect 7680 3015 7707 3049
rect 7756 3015 7775 3049
rect 7833 3015 7843 3049
rect 7910 3015 7911 3049
rect 7945 3015 7953 3049
rect 8013 3015 8030 3049
rect 8081 3015 8107 3049
rect 8149 3015 8183 3049
rect 8218 3015 8251 3049
rect 8295 3015 8319 3049
rect 8372 3015 8387 3049
rect 8449 3015 8455 3049
rect 8489 3015 8492 3049
rect 8557 3015 8569 3049
rect 8625 3015 8646 3049
rect 8693 3015 8723 3049
rect 8761 3015 8835 3049
rect 7219 3009 8835 3015
rect 7219 2981 7265 3009
rect 7219 2943 7225 2981
rect 7259 2943 7265 2981
rect 7219 2913 7265 2943
rect 7219 2869 7225 2913
rect 7259 2869 7265 2913
rect 8789 2975 8835 3009
rect 8789 2941 8795 2975
rect 8829 2941 8835 2975
rect 8789 2938 8835 2941
rect 7219 2845 7265 2869
rect 7219 2795 7225 2845
rect 7259 2795 7265 2845
rect 7219 2777 7265 2795
rect 7219 2721 7225 2777
rect 7259 2721 7265 2777
rect 7219 2709 7265 2721
rect 7219 2648 7225 2709
rect 7259 2648 7265 2709
rect 7219 2641 7265 2648
rect 7219 2575 7225 2641
rect 7259 2575 7265 2641
rect 7219 2573 7265 2575
rect 7219 2539 7225 2573
rect 7259 2539 7265 2573
rect 7219 2536 7265 2539
rect 7219 2471 7225 2536
rect 7259 2471 7265 2536
rect 7219 2463 7265 2471
rect 7219 2403 7225 2463
rect 7259 2403 7265 2463
rect 7219 2390 7265 2403
rect 7219 2335 7225 2390
rect 7259 2335 7265 2390
rect 7219 2317 7265 2335
rect 7219 2267 7225 2317
rect 7259 2267 7265 2317
rect 7219 2244 7265 2267
rect 7219 2199 7225 2244
rect 7259 2199 7265 2244
rect 7219 2171 7265 2199
rect 7219 2131 7225 2171
rect 7259 2131 7265 2171
rect 7219 2098 7265 2131
rect 7219 2063 7225 2098
rect 7259 2063 7265 2098
rect 7219 2029 7265 2063
rect 7219 1991 7225 2029
rect 7259 1991 7265 2029
rect 7219 1961 7265 1991
rect 7219 1918 7225 1961
rect 7259 1918 7265 1961
rect 7219 1893 7265 1918
rect 7370 2792 7404 2817
rect 7370 2717 7404 2749
rect 7370 2647 7404 2681
rect 7370 2579 7404 2608
rect 7370 2511 7404 2533
rect 7370 2443 7404 2458
rect 7370 2375 7404 2383
rect 7370 2307 7404 2308
rect 7370 2267 7404 2273
rect 7370 2192 7404 2205
rect 7370 2117 7404 2137
rect 7370 2042 7404 2069
rect 7370 1967 7404 2001
rect 7370 1917 7404 1933
rect 7586 2792 7620 2817
rect 7586 2717 7620 2749
rect 7586 2647 7620 2681
rect 7586 2579 7620 2608
rect 7586 2511 7620 2533
rect 7586 2443 7620 2458
rect 7586 2375 7620 2383
rect 7586 2307 7620 2308
rect 7586 2267 7620 2273
rect 7586 2192 7620 2205
rect 7586 2117 7620 2137
rect 7586 2042 7620 2069
rect 7586 1967 7620 2001
rect 7586 1917 7620 1933
rect 7802 2792 7836 2817
rect 7802 2717 7836 2749
rect 7802 2647 7836 2681
rect 7802 2579 7836 2608
rect 7802 2511 7836 2533
rect 7802 2443 7836 2458
rect 7802 2375 7836 2383
rect 7802 2307 7836 2308
rect 7802 2267 7836 2273
rect 7802 2192 7836 2205
rect 7802 2117 7836 2137
rect 7802 2042 7836 2069
rect 7802 1967 7836 2001
rect 7802 1917 7836 1933
rect 8018 2851 8052 2878
rect 8789 2904 8795 2938
rect 8829 2904 8835 2938
rect 8789 2901 8835 2904
rect 8018 2783 8052 2806
rect 8018 2715 8052 2734
rect 8018 2647 8052 2662
rect 8018 2579 8052 2590
rect 8018 2511 8052 2517
rect 8018 2443 8052 2444
rect 8018 2405 8052 2409
rect 8018 2332 8052 2341
rect 8018 2259 8052 2273
rect 8018 2186 8052 2205
rect 8018 2113 8052 2137
rect 8018 2040 8052 2069
rect 8018 1967 8052 2001
rect 8018 1917 8052 1933
rect 8174 2788 8208 2817
rect 8174 2715 8208 2749
rect 8174 2647 8208 2675
rect 8174 2579 8208 2596
rect 8174 2511 8208 2517
rect 8174 2472 8208 2477
rect 8174 2393 8208 2409
rect 8174 2314 8208 2341
rect 8174 2239 8208 2273
rect 8174 2171 8208 2200
rect 8174 2103 8208 2120
rect 8174 2035 8208 2069
rect 8174 1967 8208 2001
rect 8174 1917 8208 1933
rect 8330 2792 8364 2817
rect 8330 2717 8364 2749
rect 8330 2647 8364 2681
rect 8330 2579 8364 2608
rect 8330 2511 8364 2533
rect 8330 2443 8364 2458
rect 8330 2375 8364 2383
rect 8330 2307 8364 2308
rect 8330 2267 8364 2273
rect 8330 2192 8364 2205
rect 8330 2117 8364 2137
rect 8330 2042 8364 2069
rect 8330 1967 8364 2001
rect 8330 1917 8364 1933
rect 8486 2788 8520 2817
rect 8486 2715 8520 2749
rect 8486 2647 8520 2675
rect 8486 2579 8520 2596
rect 8486 2511 8520 2517
rect 8486 2472 8520 2477
rect 8486 2393 8520 2409
rect 8486 2314 8520 2341
rect 8486 2239 8520 2273
rect 8486 2171 8520 2200
rect 8486 2103 8520 2120
rect 8486 2035 8520 2069
rect 8486 1967 8520 2001
rect 8486 1917 8520 1933
rect 8642 2792 8676 2817
rect 8642 2717 8676 2749
rect 8642 2647 8676 2681
rect 8642 2579 8676 2608
rect 8642 2511 8676 2533
rect 8642 2443 8676 2458
rect 8642 2375 8676 2383
rect 8642 2307 8676 2308
rect 8642 2267 8676 2273
rect 8642 2192 8676 2205
rect 8642 2117 8676 2137
rect 8642 2042 8676 2069
rect 8642 1967 8676 2001
rect 8642 1917 8676 1933
rect 8789 2836 8795 2901
rect 8829 2836 8835 2901
rect 8789 2827 8835 2836
rect 8789 2768 8795 2827
rect 8829 2768 8835 2827
rect 8789 2753 8835 2768
rect 8789 2700 8795 2753
rect 8829 2700 8835 2753
rect 8789 2679 8835 2700
rect 8789 2632 8795 2679
rect 8829 2632 8835 2679
rect 8789 2605 8835 2632
rect 8789 2564 8795 2605
rect 8829 2564 8835 2605
rect 8789 2531 8835 2564
rect 8789 2496 8795 2531
rect 8829 2496 8835 2531
rect 8789 2462 8835 2496
rect 8789 2423 8795 2462
rect 8829 2423 8835 2462
rect 8789 2394 8835 2423
rect 8789 2349 8795 2394
rect 8829 2349 8835 2394
rect 8789 2326 8835 2349
rect 8789 2275 8795 2326
rect 8829 2275 8835 2326
rect 8789 2258 8835 2275
rect 8789 2201 8795 2258
rect 8829 2201 8835 2258
rect 8789 2190 8835 2201
rect 8789 2127 8795 2190
rect 8829 2127 8835 2190
rect 8789 2122 8835 2127
rect 8789 2088 8795 2122
rect 8829 2088 8835 2122
rect 8789 2086 8835 2088
rect 8789 2020 8795 2086
rect 8829 2020 8835 2086
rect 8789 2011 8835 2020
rect 8789 1952 8795 2011
rect 8829 1952 8835 2011
rect 8789 1936 8835 1952
rect 7219 1845 7225 1893
rect 7259 1845 7265 1893
rect 8789 1884 8795 1936
rect 8829 1884 8835 1936
rect 7219 1806 7265 1845
rect 7415 1839 7431 1873
rect 7485 1839 7507 1873
rect 7563 1839 7582 1873
rect 7640 1839 7657 1873
rect 7717 1839 7732 1873
rect 7794 1839 7807 1873
rect 7871 1839 7882 1873
rect 7948 1839 7957 1873
rect 7991 1839 8007 1873
rect 8063 1839 8079 1873
rect 8135 1839 8151 1873
rect 8213 1839 8223 1873
rect 8291 1839 8295 1873
rect 8329 1839 8335 1873
rect 8401 1839 8413 1873
rect 8473 1839 8490 1873
rect 8544 1839 8567 1873
rect 8615 1839 8631 1873
rect 8789 1861 8835 1884
rect 7219 1754 7225 1806
rect 7259 1754 7265 1806
rect 7219 1714 7265 1754
rect 8789 1816 8795 1861
rect 8829 1816 8835 1861
rect 8789 1786 8835 1816
rect 8789 1748 8795 1786
rect 8829 1748 8835 1786
rect 8789 1720 8835 1748
rect 7742 1714 8835 1720
rect 7219 1680 7293 1714
rect 7327 1680 7361 1714
rect 7395 1680 7429 1714
rect 7463 1680 7497 1714
rect 7531 1680 7565 1714
rect 7599 1680 7633 1714
rect 7667 1680 7701 1714
rect 7735 1680 7769 1714
rect 7814 1680 7837 1714
rect 7887 1680 7905 1714
rect 7960 1680 7973 1714
rect 8033 1680 8041 1714
rect 8106 1680 8109 1714
rect 8143 1680 8145 1714
rect 8211 1680 8218 1714
rect 8279 1680 8291 1714
rect 8347 1680 8363 1714
rect 8415 1680 8435 1714
rect 8483 1680 8507 1714
rect 8551 1680 8579 1714
rect 8619 1680 8651 1714
rect 8687 1680 8721 1714
rect 8757 1680 8835 1714
rect 7742 1674 8835 1680
rect 9012 3016 9018 3055
rect 9052 3016 9058 3055
rect 9012 2987 9058 3016
rect 9012 2942 9018 2987
rect 9052 2942 9058 2987
rect 9012 2919 9058 2942
rect 9012 2868 9018 2919
rect 9052 2868 9058 2919
rect 9012 2851 9058 2868
rect 9012 2794 9018 2851
rect 9052 2794 9058 2851
rect 9012 2783 9058 2794
rect 9012 2720 9018 2783
rect 9052 2720 9058 2783
rect 9012 2715 9058 2720
rect 9012 2681 9018 2715
rect 9052 2681 9058 2715
rect 9012 2680 9058 2681
rect 9012 2613 9018 2680
rect 9052 2613 9058 2680
rect 9012 2606 9058 2613
rect 9012 2545 9018 2606
rect 9052 2545 9058 2606
rect 9012 2532 9058 2545
rect 9012 2477 9018 2532
rect 9052 2477 9058 2532
rect 9012 2458 9058 2477
rect 9012 2409 9018 2458
rect 9052 2409 9058 2458
rect 9012 2384 9058 2409
rect 9012 2341 9018 2384
rect 9052 2341 9058 2384
rect 9012 2310 9058 2341
rect 9012 2273 9018 2310
rect 9052 2273 9058 2310
rect 9012 2239 9058 2273
rect 9012 2202 9018 2239
rect 9052 2202 9058 2239
rect 9012 2171 9058 2202
rect 9012 2128 9018 2171
rect 9052 2128 9058 2171
rect 9012 2103 9058 2128
rect 9012 2054 9018 2103
rect 9052 2054 9058 2103
rect 9012 2035 9058 2054
rect 9012 1979 9018 2035
rect 9052 1979 9058 2035
rect 9012 1967 9058 1979
rect 9012 1904 9018 1967
rect 9052 1904 9058 1967
rect 9012 1899 9058 1904
rect 9012 1865 9018 1899
rect 9052 1865 9058 1899
rect 9012 1863 9058 1865
rect 9012 1797 9018 1863
rect 9052 1797 9058 1863
rect 9012 1788 9058 1797
rect 9012 1729 9018 1788
rect 9052 1729 9058 1788
rect 9012 1713 9058 1729
rect 6993 1672 7039 1674
rect 6993 1606 6999 1672
rect 7033 1606 7039 1672
rect 6993 1600 7039 1606
rect 6993 1566 6999 1600
rect 7033 1566 7039 1600
rect 6993 1528 7039 1566
rect 6993 1494 6999 1528
rect 7033 1494 7039 1528
rect 9012 1661 9018 1713
rect 9052 1661 9058 1713
rect 9497 3088 11735 3094
rect 9497 3054 9588 3088
rect 9622 3054 9673 3088
rect 9707 3054 9759 3088
rect 9793 3054 9845 3088
rect 9879 3054 9931 3088
rect 9965 3054 10041 3088
rect 10075 3054 10116 3088
rect 10150 3054 10191 3088
rect 10225 3054 10266 3088
rect 10300 3054 10341 3088
rect 10375 3054 10416 3088
rect 10450 3054 10491 3088
rect 10525 3054 10566 3088
rect 10600 3054 10641 3088
rect 10675 3054 10716 3088
rect 10750 3054 10791 3088
rect 10825 3054 10866 3088
rect 10900 3054 10941 3088
rect 10975 3054 11016 3088
rect 11050 3054 11091 3088
rect 11125 3054 11167 3088
rect 11201 3054 11243 3088
rect 11277 3054 11319 3088
rect 11353 3054 11395 3088
rect 11429 3054 11471 3088
rect 11505 3054 11547 3088
rect 11581 3054 11623 3088
rect 11657 3054 11735 3088
rect 9497 3049 11735 3054
rect 9497 3016 9571 3049
rect 9497 2982 9503 3016
rect 9537 3015 9571 3016
rect 9605 3015 9639 3049
rect 9673 3015 9707 3049
rect 9741 3015 9775 3049
rect 9809 3015 9843 3049
rect 9877 3015 9911 3049
rect 9945 3015 9979 3049
rect 10013 3015 10047 3049
rect 10081 3015 10115 3049
rect 10149 3015 10183 3049
rect 10217 3015 10251 3049
rect 10285 3015 10319 3049
rect 10353 3015 10387 3049
rect 10421 3015 10455 3049
rect 10489 3015 10523 3049
rect 10557 3015 10591 3049
rect 10625 3015 10659 3049
rect 10693 3015 10727 3049
rect 10761 3015 10795 3049
rect 10829 3015 10863 3049
rect 10897 3015 10931 3049
rect 10965 3015 10999 3049
rect 11033 3015 11067 3049
rect 11101 3015 11135 3049
rect 11169 3015 11203 3049
rect 11237 3015 11271 3049
rect 11305 3015 11339 3049
rect 11373 3015 11407 3049
rect 11441 3015 11475 3049
rect 11509 3015 11543 3049
rect 11577 3015 11611 3049
rect 11645 3016 11735 3049
rect 11645 3015 11695 3016
rect 9537 2982 9543 3015
rect 9497 2943 9543 2982
rect 9497 2904 9503 2943
rect 9537 2904 9543 2943
rect 11689 2982 11695 3015
rect 11729 2982 11735 3016
rect 11689 2981 11735 2982
rect 11689 2947 11695 2981
rect 11729 2947 11735 2981
rect 11689 2944 11735 2947
rect 9497 2870 9543 2904
rect 9497 2836 9503 2870
rect 9537 2836 9543 2870
rect 9497 2802 9543 2836
rect 9497 2763 9503 2802
rect 9537 2763 9543 2802
rect 9497 2734 9543 2763
rect 9497 2690 9503 2734
rect 9537 2690 9543 2734
rect 9497 2666 9543 2690
rect 9497 2617 9503 2666
rect 9537 2617 9543 2666
rect 9497 2598 9543 2617
rect 9497 2544 9503 2598
rect 9537 2544 9543 2598
rect 9497 2530 9543 2544
rect 9497 2472 9503 2530
rect 9537 2472 9543 2530
rect 9497 2462 9543 2472
rect 9497 2400 9503 2462
rect 9537 2400 9543 2462
rect 9497 2394 9543 2400
rect 9497 2328 9503 2394
rect 9537 2328 9543 2394
rect 9497 2326 9543 2328
rect 9497 2292 9503 2326
rect 9537 2292 9543 2326
rect 9497 2290 9543 2292
rect 9497 2224 9503 2290
rect 9537 2224 9543 2290
rect 9497 2218 9543 2224
rect 9497 2156 9503 2218
rect 9537 2156 9543 2218
rect 9497 2146 9543 2156
rect 9497 2088 9503 2146
rect 9537 2088 9543 2146
rect 9497 2074 9543 2088
rect 9497 2020 9503 2074
rect 9537 2020 9543 2074
rect 9497 2002 9543 2020
rect 9497 1952 9503 2002
rect 9537 1952 9543 2002
rect 9497 1930 9543 1952
rect 9497 1884 9503 1930
rect 9537 1884 9543 1930
rect 9648 2851 9682 2875
rect 9648 2783 9682 2803
rect 9804 2851 9838 2867
rect 9804 2783 9838 2817
rect 9648 2715 9682 2731
rect 9648 2647 9682 2659
rect 9648 2579 9682 2587
rect 9648 2511 9682 2515
rect 9648 2405 9682 2409
rect 9648 2332 9682 2341
rect 9648 2259 9682 2273
rect 9648 2186 9682 2205
rect 9648 2113 9682 2137
rect 9648 2040 9682 2069
rect 9648 1967 9682 2001
rect 9837 2748 9838 2749
rect 9803 2715 9838 2748
rect 9803 2708 9804 2715
rect 9837 2674 9838 2681
rect 9803 2647 9838 2674
rect 9803 2634 9804 2647
rect 9837 2600 9838 2613
rect 9803 2579 9838 2600
rect 9803 2560 9804 2579
rect 9837 2526 9838 2545
rect 9803 2511 9838 2526
rect 9803 2486 9804 2511
rect 9837 2452 9838 2477
rect 9803 2443 9838 2452
rect 9803 2412 9804 2443
rect 9837 2378 9838 2409
rect 9803 2375 9838 2378
rect 9803 2341 9804 2375
rect 9803 2338 9838 2341
rect 9837 2307 9838 2338
rect 9803 2273 9804 2304
rect 9803 2264 9838 2273
rect 9837 2239 9838 2264
rect 9803 2205 9804 2230
rect 9803 2190 9838 2205
rect 9837 2171 9838 2190
rect 9803 2137 9804 2156
rect 9803 2116 9838 2137
rect 9837 2103 9838 2116
rect 9803 2069 9804 2082
rect 9803 2042 9838 2069
rect 9837 2035 9838 2042
rect 9803 2001 9804 2008
rect 9803 1967 9838 2001
rect 9648 1917 9682 1933
rect 9804 1917 9838 1933
rect 9960 2851 9994 2875
rect 9960 2783 9994 2803
rect 9960 2715 9994 2731
rect 9960 2647 9994 2659
rect 9960 2579 9994 2587
rect 9960 2511 9994 2515
rect 9960 2405 9994 2409
rect 9960 2332 9994 2341
rect 9960 2259 9994 2273
rect 9960 2186 9994 2205
rect 9960 2113 9994 2137
rect 9960 2040 9994 2069
rect 9960 1967 9994 2001
rect 9960 1917 9994 1933
rect 10116 2851 10150 2867
rect 10116 2783 10150 2817
rect 10116 2715 10150 2748
rect 10116 2647 10150 2671
rect 10116 2579 10150 2594
rect 10116 2511 10150 2517
rect 10116 2474 10150 2477
rect 10116 2397 10150 2409
rect 10116 2320 10150 2341
rect 10116 2243 10150 2273
rect 10116 2171 10150 2205
rect 10116 2103 10150 2132
rect 10116 2035 10150 2054
rect 10116 1967 10150 2001
rect 10116 1917 10150 1933
rect 10272 2851 10306 2875
rect 10272 2783 10306 2803
rect 10272 2715 10306 2731
rect 10272 2647 10306 2659
rect 10272 2579 10306 2587
rect 10272 2511 10306 2515
rect 10272 2405 10306 2409
rect 10272 2332 10306 2341
rect 10272 2259 10306 2273
rect 10272 2186 10306 2205
rect 10272 2113 10306 2137
rect 10272 2040 10306 2069
rect 10272 1967 10306 2001
rect 10272 1917 10306 1933
rect 10428 2851 10462 2867
rect 10428 2783 10462 2817
rect 10428 2715 10462 2748
rect 10428 2647 10462 2671
rect 10428 2579 10462 2594
rect 10428 2511 10462 2517
rect 10428 2474 10462 2477
rect 10428 2397 10462 2409
rect 10428 2320 10462 2341
rect 10428 2243 10462 2273
rect 10428 2171 10462 2205
rect 10428 2103 10462 2132
rect 10428 2035 10462 2054
rect 10428 1967 10462 2001
rect 10428 1917 10462 1933
rect 10584 2851 10618 2875
rect 10584 2783 10618 2803
rect 10584 2715 10618 2731
rect 10584 2647 10618 2659
rect 10584 2579 10618 2587
rect 10584 2511 10618 2515
rect 10584 2405 10618 2409
rect 10584 2332 10618 2341
rect 10584 2259 10618 2273
rect 10584 2186 10618 2205
rect 10584 2113 10618 2137
rect 10584 2040 10618 2069
rect 10584 1967 10618 2001
rect 10584 1917 10618 1933
rect 10740 2851 10774 2867
rect 10740 2810 10774 2817
rect 10740 2731 10774 2749
rect 10740 2651 10774 2681
rect 10740 2579 10774 2613
rect 10740 2511 10774 2537
rect 10740 2443 10774 2457
rect 10740 2375 10774 2377
rect 10740 2331 10774 2341
rect 10740 2251 10774 2273
rect 10740 2171 10774 2205
rect 10740 2103 10774 2137
rect 10740 2035 10774 2057
rect 10740 1967 10774 2001
rect 10740 1917 10774 1933
rect 10896 2851 10930 2875
rect 10896 2783 10930 2803
rect 10896 2715 10930 2731
rect 10896 2647 10930 2659
rect 10896 2579 10930 2587
rect 10896 2511 10930 2515
rect 10896 2405 10930 2409
rect 10896 2332 10930 2341
rect 10896 2259 10930 2273
rect 10896 2186 10930 2205
rect 10896 2113 10930 2137
rect 10896 2040 10930 2069
rect 10896 1967 10930 2001
rect 10896 1917 10930 1933
rect 11052 2851 11086 2867
rect 11052 2810 11086 2817
rect 11052 2734 11086 2749
rect 11052 2658 11086 2681
rect 11052 2582 11086 2613
rect 11052 2511 11086 2545
rect 11052 2443 11086 2472
rect 11052 2375 11086 2395
rect 11052 2307 11086 2318
rect 11052 2239 11086 2241
rect 11052 2198 11086 2205
rect 11052 2121 11086 2137
rect 11052 2044 11086 2069
rect 11052 1967 11086 2001
rect 11052 1917 11086 1933
rect 11208 2851 11242 2875
rect 11208 2783 11242 2803
rect 11208 2715 11242 2731
rect 11208 2647 11242 2659
rect 11208 2579 11242 2587
rect 11208 2511 11242 2515
rect 11208 2405 11242 2409
rect 11208 2332 11242 2341
rect 11208 2259 11242 2273
rect 11208 2186 11242 2205
rect 11208 2113 11242 2137
rect 11208 2040 11242 2069
rect 11208 1967 11242 2001
rect 11208 1917 11242 1933
rect 11364 2851 11398 2867
rect 11364 2783 11398 2817
rect 11364 2715 11398 2748
rect 11364 2647 11398 2674
rect 11364 2579 11398 2600
rect 11364 2511 11398 2526
rect 11364 2443 11398 2452
rect 11364 2375 11398 2378
rect 11364 2338 11398 2341
rect 11364 2264 11398 2273
rect 11364 2190 11398 2205
rect 11364 2116 11398 2137
rect 11364 2042 11398 2069
rect 11364 1967 11398 2001
rect 11364 1917 11398 1933
rect 11520 2851 11554 2875
rect 11520 2783 11554 2803
rect 11520 2715 11554 2731
rect 11520 2647 11554 2659
rect 11520 2579 11554 2587
rect 11520 2511 11554 2515
rect 11520 2405 11554 2409
rect 11520 2332 11554 2341
rect 11520 2259 11554 2273
rect 11520 2186 11554 2205
rect 11520 2113 11554 2137
rect 11520 2040 11554 2069
rect 11520 1967 11554 2001
rect 11520 1917 11554 1933
rect 11689 2879 11695 2944
rect 11729 2879 11735 2944
rect 11689 2872 11735 2879
rect 11689 2811 11695 2872
rect 11729 2811 11735 2872
rect 11689 2800 11735 2811
rect 11689 2743 11695 2800
rect 11729 2743 11735 2800
rect 11689 2728 11735 2743
rect 11689 2675 11695 2728
rect 11729 2675 11735 2728
rect 11689 2656 11735 2675
rect 11689 2607 11695 2656
rect 11729 2607 11735 2656
rect 11689 2584 11735 2607
rect 11689 2539 11695 2584
rect 11729 2539 11735 2584
rect 11689 2512 11735 2539
rect 11689 2471 11695 2512
rect 11729 2471 11735 2512
rect 11689 2440 11735 2471
rect 11689 2403 11695 2440
rect 11729 2403 11735 2440
rect 11689 2369 11735 2403
rect 11689 2334 11695 2369
rect 11729 2334 11735 2369
rect 11689 2301 11735 2334
rect 11689 2262 11695 2301
rect 11729 2262 11735 2301
rect 11689 2233 11735 2262
rect 11689 2190 11695 2233
rect 11729 2190 11735 2233
rect 11689 2165 11735 2190
rect 11689 2117 11695 2165
rect 11729 2117 11735 2165
rect 11689 2097 11735 2117
rect 11689 2044 11695 2097
rect 11729 2044 11735 2097
rect 11689 2029 11735 2044
rect 11689 1971 11695 2029
rect 11729 1971 11735 2029
rect 11689 1932 11735 1971
rect 9497 1858 9543 1884
rect 11689 1898 11695 1932
rect 11729 1898 11735 1932
rect 9497 1816 9503 1858
rect 9537 1816 9543 1858
rect 9693 1839 9709 1873
rect 9745 1839 9796 1873
rect 9838 1839 9881 1873
rect 9933 1839 9949 1873
rect 10005 1839 10021 1873
rect 10055 1839 10096 1873
rect 10130 1839 10170 1873
rect 10204 1839 10244 1873
rect 10278 1839 10286 1873
rect 10352 1839 10362 1873
rect 10426 1839 10437 1873
rect 10500 1839 10512 1873
rect 10574 1839 10587 1873
rect 10648 1839 10662 1873
rect 10722 1839 10737 1873
rect 10796 1839 10812 1873
rect 10870 1839 10886 1873
rect 10941 1839 10954 1873
rect 10991 1839 11047 1873
rect 11086 1839 11140 1873
rect 11181 1839 11197 1873
rect 11253 1839 11269 1873
rect 11305 1839 11364 1873
rect 11398 1839 11457 1873
rect 11493 1839 11509 1873
rect 11689 1862 11735 1898
rect 9497 1786 9543 1816
rect 9497 1748 9503 1786
rect 9537 1748 9543 1786
rect 9497 1720 9543 1748
rect 11689 1825 11695 1862
rect 11729 1825 11735 1862
rect 11689 1794 11735 1825
rect 11689 1752 11695 1794
rect 11729 1752 11735 1794
rect 11689 1720 11735 1752
rect 9497 1714 9604 1720
rect 10240 1714 11735 1720
rect 9497 1680 9517 1714
rect 9551 1680 9587 1714
rect 9621 1680 9655 1714
rect 9689 1680 9723 1714
rect 9757 1680 9791 1714
rect 9825 1680 9859 1714
rect 9893 1680 9927 1714
rect 9961 1680 9995 1714
rect 10029 1680 10063 1714
rect 10097 1680 10131 1714
rect 10165 1680 10199 1714
rect 10233 1680 10267 1714
rect 10312 1680 10335 1714
rect 10387 1680 10403 1714
rect 10462 1680 10471 1714
rect 10537 1680 10539 1714
rect 10573 1680 10578 1714
rect 10641 1680 10653 1714
rect 10709 1680 10728 1714
rect 10777 1680 10803 1714
rect 10845 1680 10878 1714
rect 10913 1680 10947 1714
rect 10987 1680 11015 1714
rect 11062 1680 11083 1714
rect 11137 1680 11151 1714
rect 11211 1680 11219 1714
rect 11285 1680 11287 1714
rect 11321 1680 11325 1714
rect 11389 1680 11399 1714
rect 11457 1680 11473 1714
rect 11525 1680 11547 1714
rect 11593 1680 11621 1714
rect 11661 1680 11735 1714
rect 9497 1674 9604 1680
rect 10240 1674 11735 1680
rect 11916 3064 17128 3070
rect 11916 3030 11994 3064
rect 12028 3030 12056 3064
rect 12100 3030 12124 3064
rect 12172 3030 12192 3064
rect 12244 3030 12260 3064
rect 12316 3030 12328 3064
rect 12388 3030 12396 3064
rect 12460 3030 12464 3064
rect 12566 3030 12570 3064
rect 12634 3030 12642 3064
rect 12702 3030 12714 3064
rect 12770 3030 12786 3064
rect 12838 3030 12858 3064
rect 12906 3030 12930 3064
rect 12974 3030 13002 3064
rect 13042 3030 13074 3064
rect 13110 3030 13144 3064
rect 13180 3030 13212 3064
rect 13252 3030 13280 3064
rect 13324 3030 13348 3064
rect 13396 3030 13416 3064
rect 13468 3030 13484 3064
rect 13540 3030 13552 3064
rect 13612 3030 13620 3064
rect 13684 3030 13688 3064
rect 13790 3030 13794 3064
rect 13858 3030 13866 3064
rect 13926 3030 13938 3064
rect 13994 3030 14010 3064
rect 14062 3030 14082 3064
rect 14130 3030 14154 3064
rect 14198 3030 14226 3064
rect 14266 3030 14298 3064
rect 14334 3030 14368 3064
rect 14404 3030 14436 3064
rect 14476 3030 14504 3064
rect 14548 3030 14572 3064
rect 14620 3030 14640 3064
rect 14692 3030 14708 3064
rect 14764 3030 14776 3064
rect 14836 3030 14844 3064
rect 14908 3030 14912 3064
rect 15014 3030 15018 3064
rect 15082 3030 15090 3064
rect 15150 3030 15162 3064
rect 15218 3030 15234 3064
rect 15286 3030 15306 3064
rect 15354 3030 15378 3064
rect 15422 3030 15450 3064
rect 15490 3030 15522 3064
rect 15558 3030 15592 3064
rect 15628 3030 15660 3064
rect 15700 3030 15728 3064
rect 15772 3030 15796 3064
rect 15844 3030 15864 3064
rect 15916 3030 15932 3064
rect 15988 3030 16000 3064
rect 16060 3030 16068 3064
rect 16132 3030 16136 3064
rect 16238 3030 16243 3064
rect 16306 3030 16316 3064
rect 16374 3030 16389 3064
rect 16442 3030 16462 3064
rect 16510 3030 16544 3064
rect 16606 3030 16612 3064
rect 16714 3030 16720 3064
rect 16782 3030 16794 3064
rect 16850 3030 16868 3064
rect 16918 3030 16942 3064
rect 16986 3030 17016 3064
rect 17054 3030 17128 3064
rect 11916 3024 17128 3030
rect 11916 2996 11962 3024
rect 11916 2958 11922 2996
rect 11956 2958 11962 2996
rect 11916 2928 11962 2958
rect 11916 2885 11922 2928
rect 11956 2885 11962 2928
rect 11916 2860 11962 2885
rect 11916 2812 11922 2860
rect 11956 2812 11962 2860
rect 11916 2792 11962 2812
rect 11916 2739 11922 2792
rect 11956 2739 11962 2792
rect 14529 2996 14575 3024
rect 14529 2962 14535 2996
rect 14569 2962 14575 2996
rect 14529 2961 14575 2962
rect 14529 2927 14535 2961
rect 14569 2927 14575 2961
rect 14529 2926 14575 2927
rect 14529 2892 14535 2926
rect 14569 2892 14575 2926
rect 14529 2887 14575 2892
rect 14529 2822 14535 2887
rect 14569 2822 14575 2887
rect 14529 2813 14575 2822
rect 12266 2744 12281 2778
rect 12336 2744 12354 2778
rect 12406 2744 12427 2778
rect 12476 2744 12500 2778
rect 12546 2744 12573 2778
rect 12616 2744 12646 2778
rect 12685 2744 12719 2778
rect 12754 2744 12789 2778
rect 12826 2744 12858 2778
rect 12899 2744 12927 2778
rect 12972 2744 12996 2778
rect 13045 2744 13065 2778
rect 13118 2744 13134 2778
rect 13191 2744 13203 2778
rect 13264 2744 13272 2778
rect 13337 2744 13341 2778
rect 13375 2744 13376 2778
rect 13444 2744 13449 2778
rect 13513 2744 13522 2778
rect 13582 2744 13595 2778
rect 13651 2744 13668 2778
rect 13720 2744 13741 2778
rect 13789 2744 13814 2778
rect 13858 2744 13887 2778
rect 13927 2744 13960 2778
rect 13996 2744 14031 2778
rect 14066 2744 14100 2778
rect 14138 2744 14169 2778
rect 14210 2744 14227 2778
rect 14529 2753 14535 2813
rect 14569 2753 14575 2813
rect 17082 2992 17128 3024
rect 17082 2942 17088 2992
rect 17122 2942 17128 2992
rect 17082 2920 17128 2942
rect 17082 2874 17088 2920
rect 17122 2874 17128 2920
rect 17082 2848 17128 2874
rect 17082 2806 17088 2848
rect 17122 2806 17128 2848
rect 11916 2724 11962 2739
rect 11916 2666 11922 2724
rect 11956 2666 11962 2724
rect 11916 2656 11962 2666
rect 14529 2739 14575 2753
rect 14853 2744 14877 2778
rect 14930 2744 14947 2778
rect 15004 2744 15017 2778
rect 15078 2744 15087 2778
rect 15152 2744 15157 2778
rect 15191 2744 15192 2778
rect 15226 2744 15227 2778
rect 15261 2744 15266 2778
rect 15330 2744 15340 2778
rect 15399 2744 15414 2778
rect 15468 2744 15488 2778
rect 15537 2744 15562 2778
rect 15606 2744 15636 2778
rect 15675 2744 15710 2778
rect 15744 2744 15779 2778
rect 15818 2744 15848 2778
rect 15892 2744 15917 2778
rect 15966 2744 15986 2778
rect 16040 2744 16055 2778
rect 16114 2744 16124 2778
rect 16188 2744 16193 2778
rect 16227 2744 16228 2778
rect 16296 2744 16302 2778
rect 16365 2744 16376 2778
rect 16434 2744 16450 2778
rect 16503 2744 16524 2778
rect 16572 2744 16598 2778
rect 16641 2744 16672 2778
rect 16710 2744 16745 2778
rect 16779 2744 16814 2778
rect 16848 2744 16872 2778
rect 17082 2776 17128 2806
rect 14529 2684 14535 2739
rect 14569 2684 14575 2739
rect 14529 2665 14575 2684
rect 11916 2593 11922 2656
rect 11956 2593 11962 2656
rect 12302 2626 12326 2660
rect 12370 2626 12400 2660
rect 12438 2626 12472 2660
rect 12508 2626 12540 2660
rect 12582 2626 12608 2660
rect 12656 2626 12676 2660
rect 12730 2626 12744 2660
rect 12804 2626 12812 2660
rect 12878 2626 12880 2660
rect 12914 2626 12918 2660
rect 12982 2626 12992 2660
rect 13050 2626 13066 2660
rect 13118 2626 13140 2660
rect 13186 2626 13214 2660
rect 13254 2626 13288 2660
rect 13322 2626 13356 2660
rect 13396 2626 13424 2660
rect 13470 2626 13492 2660
rect 13544 2626 13560 2660
rect 13618 2626 13628 2660
rect 13692 2626 13696 2660
rect 13730 2626 13732 2660
rect 13798 2626 13806 2660
rect 13866 2626 13880 2660
rect 13934 2626 13954 2660
rect 14002 2626 14028 2660
rect 14070 2626 14102 2660
rect 14138 2626 14172 2660
rect 14210 2626 14222 2660
rect 14529 2615 14535 2665
rect 14569 2615 14575 2665
rect 17082 2738 17088 2776
rect 17122 2738 17128 2776
rect 17082 2704 17128 2738
rect 17082 2670 17088 2704
rect 17122 2670 17128 2704
rect 14896 2626 14912 2660
rect 14946 2626 14980 2660
rect 15014 2626 15048 2660
rect 15082 2626 15116 2660
rect 15179 2626 15184 2660
rect 15286 2626 15291 2660
rect 15354 2626 15364 2660
rect 15422 2626 15437 2660
rect 15490 2626 15510 2660
rect 15558 2626 15583 2660
rect 15626 2626 15656 2660
rect 15694 2626 15728 2660
rect 15763 2626 15796 2660
rect 15836 2626 15864 2660
rect 15909 2626 15932 2660
rect 15982 2626 16000 2660
rect 16055 2626 16068 2660
rect 16128 2626 16136 2660
rect 16201 2626 16204 2660
rect 16238 2626 16240 2660
rect 16306 2626 16313 2660
rect 16374 2626 16386 2660
rect 16442 2626 16459 2660
rect 16510 2626 16532 2660
rect 16578 2626 16604 2660
rect 16646 2626 16676 2660
rect 16714 2626 16748 2660
rect 16782 2626 16816 2660
rect 16854 2626 16866 2660
rect 17082 2636 17128 2670
rect 11916 2588 11962 2593
rect 11916 2486 11922 2588
rect 11956 2486 11962 2588
rect 11916 2481 11962 2486
rect 11916 2418 11922 2481
rect 11956 2418 11962 2481
rect 14266 2599 14300 2615
rect 14266 2526 14300 2554
rect 14266 2453 14300 2474
rect 11916 2408 11962 2418
rect 11916 2350 11922 2408
rect 11956 2350 11962 2408
rect 12302 2390 12325 2424
rect 12370 2390 12398 2424
rect 12438 2390 12471 2424
rect 12506 2390 12540 2424
rect 12578 2390 12608 2424
rect 12651 2390 12676 2424
rect 12724 2390 12744 2424
rect 12797 2390 12812 2424
rect 12870 2390 12880 2424
rect 12943 2390 12948 2424
rect 13050 2390 13055 2424
rect 13118 2390 13128 2424
rect 13186 2390 13200 2424
rect 13254 2390 13272 2424
rect 13322 2390 13344 2424
rect 13390 2390 13416 2424
rect 13458 2390 13488 2424
rect 13526 2390 13560 2424
rect 13594 2390 13628 2424
rect 13666 2390 13696 2424
rect 13738 2390 13764 2424
rect 13810 2390 13832 2424
rect 13882 2390 13900 2424
rect 13954 2390 13968 2424
rect 14002 2390 14036 2424
rect 14070 2390 14104 2424
rect 14138 2390 14172 2424
rect 14206 2390 14222 2424
rect 11916 2335 11962 2350
rect 11916 2282 11922 2335
rect 11956 2282 11962 2335
rect 11916 2262 11962 2282
rect 11916 2214 11922 2262
rect 11956 2214 11962 2262
rect 11916 2189 11962 2214
rect 11916 2146 11922 2189
rect 11956 2146 11962 2189
rect 14266 2380 14300 2393
rect 14266 2307 14300 2312
rect 14266 2265 14300 2273
rect 12252 2154 12268 2188
rect 12302 2154 12336 2188
rect 12370 2154 12404 2188
rect 12454 2154 12472 2188
rect 12528 2154 12540 2188
rect 12602 2154 12608 2188
rect 12710 2154 12716 2188
rect 12778 2154 12789 2188
rect 12846 2154 12862 2188
rect 12914 2154 12935 2188
rect 12982 2154 13008 2188
rect 13050 2154 13081 2188
rect 13118 2154 13152 2188
rect 13188 2154 13220 2188
rect 13261 2154 13288 2188
rect 13334 2154 13356 2188
rect 13407 2154 13424 2188
rect 13480 2154 13492 2188
rect 13553 2154 13560 2188
rect 13626 2154 13628 2188
rect 13662 2154 13665 2188
rect 13730 2154 13738 2188
rect 13798 2154 13811 2188
rect 13866 2154 13884 2188
rect 13934 2154 13957 2188
rect 14002 2154 14030 2188
rect 14070 2154 14103 2188
rect 14138 2154 14172 2188
rect 14210 2154 14222 2188
rect 14266 2184 14300 2200
rect 11916 2116 11962 2146
rect 11916 2078 11922 2116
rect 11956 2078 11962 2116
rect 11916 2044 11962 2078
rect 11916 2010 11922 2044
rect 11956 2010 11962 2044
rect 11916 1976 11962 2010
rect 11916 1938 11922 1976
rect 11956 1938 11962 1976
rect 14266 2103 14300 2127
rect 14266 2022 14300 2053
rect 14266 1963 14300 1979
rect 14529 2591 14575 2615
rect 14529 2546 14535 2591
rect 14569 2546 14575 2591
rect 14529 2517 14575 2546
rect 14529 2477 14535 2517
rect 14569 2477 14575 2517
rect 14529 2443 14575 2477
rect 14529 2408 14535 2443
rect 14569 2408 14575 2443
rect 14529 2373 14575 2408
rect 14529 2335 14535 2373
rect 14569 2335 14575 2373
rect 14529 2304 14575 2335
rect 14529 2261 14535 2304
rect 14569 2261 14575 2304
rect 14529 2235 14575 2261
rect 14529 2187 14535 2235
rect 14569 2187 14575 2235
rect 14529 2166 14575 2187
rect 14529 2113 14535 2166
rect 14569 2113 14575 2166
rect 14529 2097 14575 2113
rect 14529 2039 14535 2097
rect 14569 2039 14575 2097
rect 14529 2028 14575 2039
rect 14529 1964 14535 2028
rect 14569 1964 14575 2028
rect 14529 1959 14575 1964
rect 14780 2599 14814 2615
rect 14780 2526 14814 2554
rect 14780 2453 14814 2474
rect 17082 2598 17088 2636
rect 17122 2598 17128 2636
rect 17082 2568 17128 2598
rect 17082 2525 17088 2568
rect 17122 2525 17128 2568
rect 17082 2500 17128 2525
rect 17082 2452 17088 2500
rect 17122 2452 17128 2500
rect 17082 2432 17128 2452
rect 14780 2380 14814 2393
rect 14946 2390 14971 2424
rect 15014 2390 15046 2424
rect 15082 2390 15116 2424
rect 15155 2390 15184 2424
rect 15230 2390 15252 2424
rect 15305 2390 15320 2424
rect 15380 2390 15388 2424
rect 15454 2390 15456 2424
rect 15490 2390 15494 2424
rect 15558 2390 15568 2424
rect 15626 2390 15642 2424
rect 15694 2390 15716 2424
rect 15762 2390 15790 2424
rect 15830 2390 15864 2424
rect 15898 2390 15932 2424
rect 15972 2390 16000 2424
rect 16046 2390 16068 2424
rect 16120 2390 16136 2424
rect 16194 2390 16204 2424
rect 16268 2390 16272 2424
rect 16306 2390 16308 2424
rect 16374 2390 16382 2424
rect 16442 2390 16456 2424
rect 16510 2390 16530 2424
rect 16578 2390 16604 2424
rect 16646 2390 16680 2424
rect 16714 2390 16748 2424
rect 16782 2390 16816 2424
rect 16850 2390 16866 2424
rect 14780 2307 14814 2312
rect 14780 2265 14814 2273
rect 14780 2184 14814 2200
rect 17082 2379 17088 2432
rect 17122 2379 17128 2432
rect 17082 2364 17128 2379
rect 17082 2306 17088 2364
rect 17122 2306 17128 2364
rect 17082 2296 17128 2306
rect 17082 2233 17088 2296
rect 17122 2233 17128 2296
rect 17082 2228 17128 2233
rect 14896 2154 14912 2188
rect 14946 2154 14980 2188
rect 15014 2154 15048 2188
rect 15098 2154 15116 2188
rect 15172 2154 15184 2188
rect 15246 2154 15252 2188
rect 15354 2154 15360 2188
rect 15422 2154 15433 2188
rect 15490 2154 15506 2188
rect 15558 2154 15579 2188
rect 15626 2154 15652 2188
rect 15694 2154 15725 2188
rect 15762 2154 15796 2188
rect 15832 2154 15864 2188
rect 15905 2154 15932 2188
rect 15978 2154 16000 2188
rect 16051 2154 16068 2188
rect 16124 2154 16136 2188
rect 16197 2154 16204 2188
rect 16270 2154 16272 2188
rect 16306 2154 16309 2188
rect 16374 2154 16382 2188
rect 16442 2154 16455 2188
rect 16510 2154 16528 2188
rect 16578 2154 16601 2188
rect 16646 2154 16674 2188
rect 16714 2154 16747 2188
rect 16782 2154 16816 2188
rect 16854 2154 16866 2188
rect 14780 2103 14814 2127
rect 14780 2022 14814 2053
rect 14780 1963 14814 1979
rect 17082 2126 17088 2228
rect 17122 2126 17128 2228
rect 17082 2121 17128 2126
rect 17082 2058 17088 2121
rect 17122 2058 17128 2121
rect 17082 2048 17128 2058
rect 17082 1990 17088 2048
rect 17122 1990 17128 2048
rect 17082 1975 17128 1990
rect 11916 1908 11962 1938
rect 12302 1918 12325 1952
rect 12370 1918 12398 1952
rect 12438 1918 12471 1952
rect 12506 1918 12540 1952
rect 12578 1918 12608 1952
rect 12651 1918 12676 1952
rect 12724 1918 12744 1952
rect 12797 1918 12812 1952
rect 12870 1918 12880 1952
rect 12943 1918 12948 1952
rect 13050 1918 13055 1952
rect 13118 1918 13128 1952
rect 13186 1918 13200 1952
rect 13254 1918 13272 1952
rect 13322 1918 13344 1952
rect 13390 1918 13416 1952
rect 13458 1918 13488 1952
rect 13526 1918 13560 1952
rect 13594 1918 13628 1952
rect 13666 1918 13696 1952
rect 13738 1918 13764 1952
rect 13810 1918 13832 1952
rect 13882 1918 13900 1952
rect 13954 1918 13968 1952
rect 14002 1918 14036 1952
rect 14070 1918 14104 1952
rect 14138 1918 14172 1952
rect 14206 1918 14222 1952
rect 14529 1925 14535 1959
rect 14569 1925 14575 1959
rect 14529 1923 14575 1925
rect 11916 1866 11922 1908
rect 11956 1866 11962 1908
rect 11916 1828 11962 1866
rect 11916 1794 11922 1828
rect 11956 1794 11962 1828
rect 11916 1776 11962 1794
rect 11916 1722 11922 1776
rect 11956 1722 11962 1776
rect 11916 1690 11962 1722
rect 14529 1856 14535 1923
rect 14569 1856 14575 1923
rect 14946 1918 14971 1952
rect 15014 1918 15046 1952
rect 15082 1918 15116 1952
rect 15155 1918 15184 1952
rect 15230 1918 15252 1952
rect 15305 1918 15320 1952
rect 15380 1918 15388 1952
rect 15454 1918 15456 1952
rect 15490 1918 15494 1952
rect 15558 1918 15568 1952
rect 15626 1918 15642 1952
rect 15694 1918 15716 1952
rect 15762 1918 15790 1952
rect 15830 1918 15864 1952
rect 15898 1918 15932 1952
rect 15972 1918 16000 1952
rect 16046 1918 16068 1952
rect 16120 1918 16136 1952
rect 16194 1918 16204 1952
rect 16268 1918 16272 1952
rect 16306 1918 16308 1952
rect 16374 1918 16382 1952
rect 16442 1918 16456 1952
rect 16510 1918 16530 1952
rect 16578 1918 16604 1952
rect 16646 1918 16680 1952
rect 16714 1918 16748 1952
rect 16782 1918 16816 1952
rect 16850 1918 16866 1952
rect 17082 1922 17088 1975
rect 17122 1922 17128 1975
rect 14529 1848 14575 1856
rect 14529 1787 14535 1848
rect 14569 1787 14575 1848
rect 14529 1773 14575 1787
rect 14529 1718 14535 1773
rect 14569 1718 14575 1773
rect 14529 1690 14575 1718
rect 17082 1902 17128 1922
rect 17082 1854 17088 1902
rect 17122 1854 17128 1902
rect 17082 1829 17128 1854
rect 17082 1786 17088 1829
rect 17122 1786 17128 1829
rect 17082 1756 17128 1786
rect 17082 1718 17088 1756
rect 17122 1718 17128 1756
rect 17082 1690 17128 1718
rect 11916 1684 15661 1690
rect 15817 1684 17128 1690
rect 9012 1638 9058 1661
rect 11916 1650 11990 1684
rect 12028 1650 12058 1684
rect 12102 1650 12126 1684
rect 12176 1650 12194 1684
rect 12250 1650 12262 1684
rect 12324 1650 12330 1684
rect 12432 1650 12438 1684
rect 12500 1650 12512 1684
rect 12568 1650 12586 1684
rect 12636 1650 12660 1684
rect 12704 1650 12734 1684
rect 12772 1650 12806 1684
rect 12842 1650 12874 1684
rect 12916 1650 12942 1684
rect 12990 1650 13010 1684
rect 13064 1650 13078 1684
rect 13138 1650 13146 1684
rect 13212 1650 13214 1684
rect 13248 1650 13252 1684
rect 13316 1650 13326 1684
rect 13384 1650 13399 1684
rect 13452 1650 13472 1684
rect 13520 1650 13545 1684
rect 13588 1650 13618 1684
rect 13656 1650 13690 1684
rect 13725 1650 13758 1684
rect 13798 1650 13826 1684
rect 13871 1650 13894 1684
rect 13944 1650 13962 1684
rect 14017 1650 14030 1684
rect 14090 1650 14098 1684
rect 14163 1650 14166 1684
rect 14200 1650 14202 1684
rect 14268 1650 14275 1684
rect 14336 1650 14348 1684
rect 14404 1650 14421 1684
rect 14472 1650 14494 1684
rect 14540 1650 14567 1684
rect 14608 1650 14640 1684
rect 14676 1650 14710 1684
rect 14747 1650 14778 1684
rect 14820 1650 14846 1684
rect 14893 1650 14914 1684
rect 14966 1650 14982 1684
rect 15039 1650 15050 1684
rect 15112 1650 15118 1684
rect 15185 1650 15186 1684
rect 15220 1650 15224 1684
rect 15288 1650 15297 1684
rect 15356 1650 15370 1684
rect 15424 1650 15443 1684
rect 15492 1650 15516 1684
rect 15560 1650 15589 1684
rect 15628 1650 15662 1684
rect 15696 1650 15730 1684
rect 15764 1650 15798 1684
rect 15832 1650 15855 1684
rect 15900 1650 15929 1684
rect 15968 1650 16002 1684
rect 16037 1650 16070 1684
rect 16111 1650 16138 1684
rect 16185 1650 16206 1684
rect 16259 1650 16274 1684
rect 16333 1650 16342 1684
rect 16407 1650 16410 1684
rect 16444 1650 16447 1684
rect 16512 1650 16521 1684
rect 16580 1650 16595 1684
rect 16648 1650 16668 1684
rect 16716 1650 16741 1684
rect 16784 1650 16814 1684
rect 16852 1650 16886 1684
rect 16921 1650 16954 1684
rect 16994 1650 17128 1684
rect 11916 1644 15661 1650
rect 15817 1644 17128 1650
rect 9012 1593 9018 1638
rect 9052 1593 9058 1638
rect 9012 1563 9058 1593
rect 9012 1525 9018 1563
rect 9052 1525 9058 1563
rect 9012 1497 9058 1525
rect 6993 1491 7039 1494
rect 7761 1491 9058 1497
rect 6905 1458 7067 1491
rect 6629 1457 6663 1458
rect 6697 1457 6731 1458
rect 6765 1457 6799 1458
rect 6833 1457 7067 1458
rect 7101 1457 7135 1491
rect 7169 1457 7203 1491
rect 7237 1457 7271 1491
rect 7305 1457 7339 1491
rect 7373 1457 7407 1491
rect 7441 1457 7475 1491
rect 7509 1457 7543 1491
rect 7577 1457 7611 1491
rect 7645 1457 7679 1491
rect 7713 1457 7747 1491
rect 7781 1457 7799 1491
rect 7849 1457 7876 1491
rect 7917 1457 7951 1491
rect 7987 1457 8019 1491
rect 8064 1457 8087 1491
rect 8140 1457 8155 1491
rect 8216 1457 8223 1491
rect 8257 1457 8258 1491
rect 8325 1457 8334 1491
rect 8393 1457 8410 1491
rect 8461 1457 8486 1491
rect 8529 1457 8562 1491
rect 8597 1457 8631 1491
rect 8672 1457 8699 1491
rect 8748 1457 8767 1491
rect 8824 1457 8835 1491
rect 8900 1457 8903 1491
rect 8937 1457 8942 1491
rect 8976 1457 9058 1491
rect 210 1400 4935 1449
rect 5098 1421 9058 1457
rect 5098 1387 5910 1421
rect 5944 1387 6000 1421
rect 6034 1387 6091 1421
rect 6125 1387 9058 1421
rect 3987 1196 4003 1230
rect 4037 1196 4072 1230
rect 4106 1196 4141 1230
rect 4175 1196 4210 1230
rect 4244 1196 4279 1230
rect 4313 1196 4348 1230
rect 4382 1196 4417 1230
rect 4451 1196 4486 1230
rect 4520 1196 4555 1230
rect 4589 1196 4624 1230
rect 4658 1196 4693 1230
rect 4727 1196 4761 1230
rect 4795 1196 4829 1230
rect 4863 1196 4897 1230
rect 4931 1196 4965 1230
rect 4999 1196 5033 1230
rect 5067 1196 5101 1230
rect 5135 1196 5169 1230
rect 5203 1196 5237 1230
rect 5271 1196 5305 1230
rect 5339 1196 5373 1230
rect 5407 1196 5441 1230
rect 5475 1196 5509 1230
rect 5543 1196 5577 1230
rect 5611 1196 5627 1230
rect 6703 1196 6719 1230
rect 6772 1196 6810 1230
rect 6848 1196 6909 1230
rect 6943 1196 6959 1230
rect 7015 1196 7029 1230
rect 7065 1196 7099 1230
rect 7135 1196 7149 1230
rect 7255 1196 7293 1230
rect 7331 1196 7365 1230
rect 7399 1196 7415 1230
rect 7547 1196 7563 1230
rect 7626 1196 7631 1230
rect 7665 1196 7668 1230
rect 7733 1196 7744 1230
rect 7801 1196 7820 1230
rect 7869 1196 7896 1230
rect 7937 1196 7971 1230
rect 8006 1196 8039 1230
rect 8082 1196 8107 1230
rect 8158 1196 8176 1230
rect 8234 1196 8245 1230
rect 8310 1196 8314 1230
rect 8348 1196 8383 1230
rect 8417 1196 8452 1230
rect 8486 1196 8521 1230
rect 8555 1196 8571 1230
rect 8627 1196 8643 1230
rect 8677 1196 8711 1230
rect 8745 1196 8779 1230
rect 8813 1196 8847 1230
rect 8881 1196 8915 1230
rect 8949 1196 8983 1230
rect 9017 1196 9051 1230
rect 9085 1196 9119 1230
rect 9153 1196 9187 1230
rect 9221 1196 9255 1230
rect 9289 1196 9323 1230
rect 9357 1196 9391 1230
rect 9425 1196 9459 1230
rect 9493 1196 9527 1230
rect 9561 1196 9595 1230
rect 9629 1196 9664 1230
rect 9698 1196 9705 1230
rect 9767 1196 9780 1230
rect 9836 1196 9855 1230
rect 9905 1196 9930 1230
rect 9974 1196 10005 1230
rect 10043 1196 10078 1230
rect 10114 1196 10147 1230
rect 10189 1196 10216 1230
rect 10264 1196 10285 1230
rect 10339 1196 10354 1230
rect 10414 1196 10423 1230
rect 10489 1196 10492 1230
rect 10526 1196 10530 1230
rect 10595 1196 10605 1230
rect 10664 1196 10680 1230
rect 10733 1196 10755 1230
rect 10802 1196 10830 1230
rect 10871 1196 10905 1230
rect 10940 1196 10975 1230
rect 11014 1196 11044 1230
rect 11089 1196 11113 1230
rect 11147 1196 11163 1230
rect 11219 1196 11235 1230
rect 11291 1196 11303 1230
rect 11364 1196 11371 1230
rect 11437 1196 11439 1230
rect 11473 1196 11476 1230
rect 11541 1196 11549 1230
rect 11609 1196 11622 1230
rect 11677 1196 11695 1230
rect 11745 1196 11768 1230
rect 11813 1196 11841 1230
rect 11881 1196 11914 1230
rect 11949 1196 11983 1230
rect 12021 1196 12051 1230
rect 12094 1196 12119 1230
rect 12167 1196 12187 1230
rect 12240 1196 12255 1230
rect 12313 1196 12323 1230
rect 12386 1196 12391 1230
rect 12493 1196 12498 1230
rect 12561 1196 12571 1230
rect 12629 1196 12644 1230
rect 12697 1196 12717 1230
rect 12765 1196 12790 1230
rect 12833 1196 12863 1230
rect 12901 1196 12935 1230
rect 12970 1196 13003 1230
rect 13043 1196 13071 1230
rect 13116 1196 13139 1230
rect 13189 1196 13207 1230
rect 13262 1196 13276 1230
rect 13335 1196 13345 1230
rect 13408 1196 13414 1230
rect 13481 1196 13483 1230
rect 13517 1196 13520 1230
rect 13586 1196 13593 1230
rect 13655 1196 13666 1230
rect 13724 1196 13739 1230
rect 13793 1196 13812 1230
rect 13862 1196 13885 1230
rect 13931 1196 13958 1230
rect 14000 1196 14031 1230
rect 14069 1196 14104 1230
rect 14138 1196 14173 1230
rect 14211 1196 14242 1230
rect 14284 1196 14311 1230
rect 14357 1196 14380 1230
rect 14430 1196 14449 1230
rect 14503 1196 14518 1230
rect 14576 1196 14587 1230
rect 14649 1196 14656 1230
rect 14722 1196 14725 1230
rect 14759 1196 14761 1230
rect 14828 1196 14833 1230
rect 14897 1196 14905 1230
rect 14966 1196 14977 1230
rect 15035 1196 15051 1230
rect 15217 1196 15233 1230
rect 15286 1196 15367 1230
rect 15403 1196 15417 1230
rect 15583 1196 15599 1230
rect 15633 1196 15677 1230
rect 15711 1196 15755 1230
rect 15789 1196 15829 1230
rect 15866 1196 15909 1230
rect 15947 1196 15959 1230
rect 5900 1130 5934 1146
rect 3942 1078 3976 1094
rect 1524 1032 1588 1066
rect 1647 1032 1656 1066
rect 1723 1032 1724 1066
rect 1758 1032 1765 1066
rect 1826 1032 1841 1066
rect 1894 1032 1917 1066
rect 1962 1032 1993 1066
rect 2030 1032 2064 1066
rect 2103 1032 2132 1066
rect 2179 1032 2200 1066
rect 2255 1032 2268 1066
rect 2330 1032 2336 1066
rect 2954 1034 2966 1066
rect 3000 1066 3049 1068
rect 3083 1066 3132 1068
rect 3166 1066 3215 1068
rect 3249 1066 3299 1068
rect 3333 1066 3383 1068
rect 3000 1034 3023 1066
rect 3083 1034 3091 1066
rect 2954 1032 3023 1034
rect 3057 1032 3091 1034
rect 3125 1034 3132 1066
rect 3193 1034 3215 1066
rect 3125 1032 3159 1034
rect 3193 1032 3227 1034
rect 3261 1032 3295 1066
rect 3333 1034 3363 1066
rect 3417 1034 3431 1066
rect 3329 1032 3363 1034
rect 3397 1032 3431 1034
rect 3942 1019 3976 1044
rect 3942 946 3976 976
rect 3942 874 3976 908
rect 2260 754 2294 792
rect 3172 759 3206 797
rect 3942 806 3976 839
rect 3942 738 3976 766
rect 3942 670 3976 693
rect 3942 602 3976 620
rect 3942 534 3976 547
rect 3942 466 3976 473
rect 1685 376 1719 414
rect 1789 327 1823 365
rect 1895 383 1929 422
rect 2151 377 2185 415
rect 3085 383 3119 421
rect 3257 386 3291 424
rect 3942 398 3976 399
rect 3942 359 3976 364
rect 3942 285 3976 296
rect 3942 194 3976 228
rect 3942 144 3976 160
rect 4048 1082 4082 1094
rect 4048 1010 4082 1044
rect 4048 942 4082 976
rect 4048 874 4082 904
rect 4048 806 4082 832
rect 4048 738 4082 760
rect 4048 670 4082 688
rect 4048 602 4082 616
rect 4048 534 4082 543
rect 4048 466 4082 470
rect 4048 431 4082 432
rect 4048 358 4082 364
rect 4048 285 4082 296
rect 4048 194 4082 228
rect 4048 144 4082 160
rect 4154 1082 4188 1094
rect 4154 1010 4188 1044
rect 4154 942 4188 976
rect 4154 874 4188 904
rect 4154 806 4188 832
rect 4154 738 4188 760
rect 4154 670 4188 688
rect 4154 602 4188 616
rect 4154 534 4188 543
rect 4154 466 4188 470
rect 4154 431 4188 432
rect 4154 358 4188 364
rect 4154 285 4188 296
rect 4154 194 4188 228
rect 4154 144 4188 160
rect 4260 1082 4294 1094
rect 4260 1010 4294 1044
rect 4260 942 4294 976
rect 4260 874 4294 904
rect 4260 806 4294 832
rect 4260 738 4294 760
rect 4260 670 4294 688
rect 4260 602 4294 616
rect 4260 534 4294 543
rect 4260 466 4294 470
rect 4260 431 4294 432
rect 4260 358 4294 364
rect 4260 285 4294 296
rect 4260 194 4294 228
rect 4260 144 4294 160
rect 4366 1082 4400 1094
rect 4366 1010 4400 1044
rect 4366 942 4400 976
rect 4366 874 4400 904
rect 4366 806 4400 832
rect 4366 738 4400 760
rect 4366 670 4400 688
rect 4366 602 4400 616
rect 4366 534 4400 543
rect 4366 466 4400 470
rect 4366 431 4400 432
rect 4366 358 4400 364
rect 4366 285 4400 296
rect 4366 194 4400 228
rect 4366 144 4400 160
rect 4472 1082 4506 1094
rect 4472 1010 4506 1044
rect 4472 942 4506 976
rect 4472 874 4506 904
rect 4472 806 4506 832
rect 4472 738 4506 760
rect 4472 670 4506 688
rect 4472 602 4506 616
rect 4472 534 4506 543
rect 4472 466 4506 470
rect 4472 431 4506 432
rect 4472 358 4506 364
rect 4472 285 4506 296
rect 4472 194 4506 228
rect 4472 144 4506 160
rect 4578 1082 4612 1094
rect 4578 1010 4612 1044
rect 4578 942 4612 976
rect 4578 874 4612 904
rect 4578 806 4612 832
rect 4578 738 4612 760
rect 4578 670 4612 688
rect 4578 602 4612 616
rect 4578 534 4612 543
rect 4578 466 4612 470
rect 4578 431 4612 432
rect 4578 358 4612 364
rect 4578 285 4612 296
rect 4578 194 4612 228
rect 4578 144 4612 160
rect 4684 1082 4718 1094
rect 4684 1010 4718 1044
rect 4684 942 4718 976
rect 4684 874 4718 904
rect 4684 806 4718 832
rect 4684 738 4718 760
rect 4684 670 4718 688
rect 4684 602 4718 616
rect 4684 534 4718 543
rect 4684 466 4718 470
rect 4684 431 4718 432
rect 4684 358 4718 364
rect 4684 285 4718 296
rect 4684 194 4718 228
rect 4684 144 4718 160
rect 4790 1082 4824 1094
rect 4790 1010 4824 1044
rect 4790 942 4824 976
rect 4790 874 4824 904
rect 4790 806 4824 832
rect 4790 738 4824 760
rect 4790 670 4824 688
rect 4790 602 4824 616
rect 4790 534 4824 543
rect 4790 466 4824 470
rect 4790 431 4824 432
rect 4790 358 4824 364
rect 4790 285 4824 296
rect 4790 194 4824 228
rect 4790 144 4824 160
rect 4896 1082 4930 1094
rect 4896 1010 4930 1044
rect 4896 942 4930 976
rect 4896 874 4930 904
rect 4896 806 4930 832
rect 4896 738 4930 760
rect 4896 670 4930 688
rect 4896 602 4930 616
rect 4896 534 4930 543
rect 4896 466 4930 470
rect 4896 431 4930 432
rect 4896 358 4930 364
rect 4896 285 4930 296
rect 4896 194 4930 228
rect 4896 144 4930 160
rect 5002 1082 5036 1094
rect 5002 1010 5036 1044
rect 5002 942 5036 976
rect 5002 874 5036 904
rect 5002 806 5036 832
rect 5002 738 5036 760
rect 5002 670 5036 688
rect 5002 602 5036 616
rect 5002 534 5036 543
rect 5002 466 5036 470
rect 5002 431 5036 432
rect 5002 358 5036 364
rect 5002 285 5036 296
rect 5002 194 5036 228
rect 5002 144 5036 160
rect 5108 1082 5142 1094
rect 5108 1010 5142 1044
rect 5108 942 5142 976
rect 5108 874 5142 904
rect 5108 806 5142 832
rect 5108 738 5142 760
rect 5108 670 5142 688
rect 5108 602 5142 616
rect 5108 534 5142 543
rect 5108 466 5142 470
rect 5108 431 5142 432
rect 5108 358 5142 364
rect 5108 285 5142 296
rect 5108 194 5142 228
rect 5108 144 5142 160
rect 5214 1082 5248 1094
rect 5214 1010 5248 1044
rect 5214 942 5248 976
rect 5214 874 5248 904
rect 5214 806 5248 832
rect 5214 738 5248 760
rect 5214 670 5248 688
rect 5214 602 5248 616
rect 5214 534 5248 543
rect 5214 466 5248 470
rect 5214 431 5248 432
rect 5214 358 5248 364
rect 5214 285 5248 296
rect 5214 194 5248 228
rect 5214 144 5248 160
rect 5320 1082 5354 1094
rect 5320 1010 5354 1044
rect 5320 942 5354 976
rect 5320 874 5354 904
rect 5320 806 5354 832
rect 5320 738 5354 760
rect 5320 670 5354 688
rect 5320 602 5354 616
rect 5320 534 5354 543
rect 5320 466 5354 470
rect 5320 431 5354 432
rect 5320 358 5354 364
rect 5320 285 5354 296
rect 5320 194 5354 228
rect 5320 144 5354 160
rect 5426 1082 5460 1094
rect 5426 1010 5460 1044
rect 5426 942 5460 976
rect 5426 874 5460 904
rect 5426 806 5460 832
rect 5426 738 5460 760
rect 5426 670 5460 688
rect 5426 602 5460 616
rect 5426 534 5460 543
rect 5426 466 5460 470
rect 5426 431 5460 432
rect 5426 358 5460 364
rect 5426 285 5460 296
rect 5426 194 5460 228
rect 5426 144 5460 160
rect 5532 1082 5566 1094
rect 5532 1010 5566 1044
rect 5532 942 5566 976
rect 5532 874 5566 904
rect 5532 806 5566 832
rect 5532 738 5566 760
rect 5532 670 5566 688
rect 5532 602 5566 616
rect 5532 534 5566 543
rect 5532 466 5566 470
rect 5532 431 5566 432
rect 5532 358 5566 364
rect 5532 285 5566 296
rect 5532 194 5566 228
rect 5532 144 5566 160
rect 5638 1082 5672 1094
rect 5638 1010 5672 1044
rect 5638 942 5672 976
rect 5900 1062 5934 1096
rect 5900 994 5934 1020
rect 5900 944 5934 948
rect 6116 1074 6150 1096
rect 6116 994 6150 1028
rect 6116 944 6150 960
rect 6332 1130 6366 1146
rect 6332 1062 6366 1096
rect 6548 1074 6582 1096
rect 6332 1020 6333 1028
rect 6332 994 6367 1020
rect 6366 982 6367 994
rect 6332 948 6333 960
rect 6548 994 6582 1028
rect 6332 944 6366 948
rect 6548 944 6582 960
rect 6658 1027 6692 1036
rect 6658 954 6692 968
rect 5638 874 5672 904
rect 5945 866 5957 900
rect 5995 866 6037 900
rect 6074 866 6112 900
rect 6157 866 6187 900
rect 6240 866 6262 900
rect 6323 866 6337 900
rect 6371 866 6372 900
rect 6406 866 6412 900
rect 6446 866 6455 900
rect 6521 866 6537 900
rect 6658 880 6692 900
rect 5638 806 5672 832
rect 5638 738 5672 760
rect 5638 670 5672 688
rect 5638 602 5672 616
rect 5900 804 5934 816
rect 5900 732 5934 766
rect 5900 664 5934 698
rect 5900 614 5934 630
rect 6116 800 6150 816
rect 6116 732 6150 766
rect 6116 664 6150 678
rect 6332 804 6366 816
rect 6332 800 6333 804
rect 6366 766 6367 770
rect 6332 732 6367 766
rect 6548 800 6582 816
rect 6548 732 6582 766
rect 6332 664 6366 698
rect 6332 614 6366 630
rect 6548 664 6582 678
rect 6658 806 6692 832
rect 6658 732 6692 764
rect 6658 662 6692 696
rect 5638 534 5672 543
rect 6658 594 6692 624
rect 5945 494 5957 528
rect 5995 494 6037 528
rect 6074 494 6112 528
rect 6157 494 6187 528
rect 6240 494 6262 528
rect 6323 494 6337 528
rect 6371 494 6372 528
rect 6406 494 6412 528
rect 6446 494 6455 528
rect 6521 494 6537 528
rect 6658 510 6692 550
rect 6814 1020 6848 1036
rect 6814 940 6848 968
rect 6814 866 6848 900
rect 6814 798 6848 825
rect 6814 730 6848 744
rect 6814 662 6848 663
rect 6814 616 6848 628
rect 6814 544 6848 560
rect 6970 1070 7004 1086
rect 6970 1002 7004 1036
rect 6970 934 7004 952
rect 6970 866 7004 874
rect 6970 830 7004 832
rect 6970 752 7004 764
rect 6970 674 7004 696
rect 6970 595 7004 628
rect 5638 466 5672 470
rect 5638 431 5672 432
rect 5638 358 5672 364
rect 5638 285 5672 296
rect 5900 378 5934 400
rect 5900 298 5934 332
rect 5900 248 5934 264
rect 6116 434 6150 450
rect 6116 366 6150 400
rect 6116 298 6150 324
rect 6116 248 6150 252
rect 6332 378 6366 400
rect 6332 298 6366 332
rect 6332 248 6366 264
rect 6548 434 6582 450
rect 6658 436 6692 476
rect 6970 516 7004 560
rect 7126 1020 7160 1036
rect 7126 940 7160 968
rect 7126 866 7160 900
rect 7126 798 7160 825
rect 7126 730 7160 744
rect 7126 662 7160 663
rect 7126 616 7160 628
rect 7126 544 7160 560
rect 7236 1078 7270 1094
rect 7236 1010 7270 1044
rect 7236 942 7270 952
rect 7236 874 7270 878
rect 7236 838 7270 840
rect 7236 764 7270 772
rect 7236 690 7270 704
rect 7236 616 7270 636
rect 6970 437 7004 482
rect 7236 541 7270 568
rect 7236 466 7270 500
rect 6548 366 6582 400
rect 6548 298 6582 324
rect 6548 248 6582 252
rect 7236 398 7270 432
rect 7236 330 7270 357
rect 7236 262 7270 282
rect 5638 194 5672 228
rect 5638 144 5672 160
rect 7236 194 7270 207
rect 7392 1082 7426 1094
rect 7392 1010 7426 1044
rect 7392 942 7426 970
rect 7392 874 7426 892
rect 7392 806 7426 814
rect 7392 770 7426 772
rect 7392 692 7426 704
rect 7392 614 7426 636
rect 7392 536 7426 568
rect 7392 466 7426 500
rect 7392 398 7426 424
rect 7392 330 7426 346
rect 7392 262 7426 267
rect 7392 222 7426 228
rect 7392 144 7426 160
rect 7502 1019 7536 1044
rect 7502 944 7536 976
rect 7502 874 7536 908
rect 7502 806 7536 835
rect 7502 738 7536 760
rect 7502 670 7536 685
rect 7502 602 7536 610
rect 7502 534 7536 535
rect 7502 494 7536 500
rect 7502 419 7536 432
rect 7502 344 7536 364
rect 7502 269 7536 296
rect 7502 194 7536 228
rect 7502 144 7536 160
rect 7718 1078 7752 1094
rect 7718 1010 7752 1044
rect 7718 942 7752 974
rect 7718 874 7752 900
rect 7718 806 7752 826
rect 7718 738 7752 752
rect 7718 670 7752 678
rect 7718 602 7752 604
rect 7718 564 7752 568
rect 7718 490 7752 500
rect 7718 416 7752 432
rect 7718 342 7752 364
rect 7718 268 7752 296
rect 7718 194 7752 228
rect 7718 144 7752 160
rect 7934 1019 7968 1044
rect 7934 944 7968 976
rect 7934 874 7968 908
rect 7934 806 7968 835
rect 7934 738 7968 760
rect 7934 670 7968 685
rect 7934 602 7968 610
rect 7934 534 7968 535
rect 7934 494 7968 500
rect 7934 419 7968 432
rect 7934 344 7968 364
rect 7934 269 7968 296
rect 7934 194 7968 228
rect 7934 144 7968 160
rect 8150 1078 8184 1094
rect 8150 1010 8184 1044
rect 8150 942 8184 976
rect 8150 886 8184 908
rect 8150 810 8184 840
rect 8150 738 8184 772
rect 8150 670 8184 699
rect 8150 602 8184 622
rect 8150 534 8184 545
rect 8150 466 8184 468
rect 8150 425 8184 432
rect 8150 348 8184 364
rect 8150 271 8184 296
rect 8150 194 8184 228
rect 8150 144 8184 160
rect 8366 1019 8400 1044
rect 8366 944 8400 976
rect 8366 874 8400 908
rect 8366 806 8400 835
rect 8366 738 8400 760
rect 8366 670 8400 685
rect 8366 602 8400 610
rect 8366 534 8400 535
rect 8366 494 8400 500
rect 8366 419 8400 432
rect 8366 344 8400 364
rect 8366 269 8400 296
rect 8366 194 8400 228
rect 8366 144 8400 160
rect 8582 1078 8616 1094
rect 8582 1010 8616 1044
rect 8582 942 8616 974
rect 8582 874 8616 900
rect 8582 806 8616 826
rect 8582 738 8616 752
rect 8582 670 8616 678
rect 8582 602 8616 604
rect 8582 564 8616 568
rect 8582 490 8616 500
rect 8582 416 8616 432
rect 8582 342 8616 364
rect 8582 268 8616 296
rect 8582 194 8616 228
rect 8582 144 8616 160
rect 8798 1078 8832 1094
rect 8798 1010 8832 1044
rect 8798 942 8832 974
rect 8798 874 8832 900
rect 8798 806 8832 826
rect 8798 738 8832 752
rect 8798 670 8832 678
rect 8798 602 8832 604
rect 8798 564 8832 568
rect 8798 490 8832 500
rect 8798 416 8832 432
rect 8798 342 8832 364
rect 8798 268 8832 296
rect 8798 194 8832 228
rect 8798 144 8832 160
rect 9014 1078 9048 1094
rect 9014 1010 9048 1044
rect 9014 942 9048 974
rect 9014 874 9048 900
rect 9014 806 9048 826
rect 9014 738 9048 752
rect 9014 670 9048 678
rect 9014 602 9048 604
rect 9014 564 9048 568
rect 9014 490 9048 500
rect 9014 416 9048 432
rect 9014 342 9048 364
rect 9014 268 9048 296
rect 9014 194 9048 228
rect 9014 144 9048 160
rect 9230 1078 9264 1094
rect 9230 1010 9264 1044
rect 9230 942 9264 974
rect 9230 874 9264 900
rect 9230 806 9264 826
rect 9230 738 9264 752
rect 9230 670 9264 678
rect 9230 602 9264 604
rect 9230 564 9264 568
rect 9230 490 9264 500
rect 9230 416 9264 432
rect 9230 342 9264 364
rect 9230 268 9264 296
rect 9230 194 9264 228
rect 9230 144 9264 160
rect 9446 1078 9480 1094
rect 9446 1010 9480 1044
rect 9446 942 9480 974
rect 9446 874 9480 900
rect 9446 806 9480 826
rect 9446 738 9480 752
rect 9446 670 9480 678
rect 9446 602 9480 604
rect 9446 564 9480 568
rect 9446 490 9480 500
rect 9446 416 9480 432
rect 9446 342 9480 364
rect 9446 268 9480 296
rect 9446 194 9480 228
rect 9446 144 9480 160
rect 9662 1078 9696 1094
rect 9662 1010 9696 1044
rect 9662 942 9696 974
rect 9662 874 9696 900
rect 9662 806 9696 826
rect 9662 738 9696 752
rect 9662 670 9696 678
rect 9662 602 9696 604
rect 9662 564 9696 568
rect 9662 490 9696 500
rect 9662 416 9696 432
rect 9662 342 9696 364
rect 9662 268 9696 296
rect 9662 194 9696 228
rect 9662 144 9696 160
rect 9878 1019 9912 1044
rect 9878 944 9912 976
rect 9878 874 9912 908
rect 9878 806 9912 835
rect 9878 738 9912 760
rect 9878 670 9912 685
rect 9878 602 9912 610
rect 9878 534 9912 535
rect 9878 494 9912 500
rect 9878 419 9912 432
rect 9878 344 9912 364
rect 9878 269 9912 296
rect 9878 194 9912 228
rect 9878 144 9912 160
rect 10094 1019 10128 1044
rect 10094 944 10128 976
rect 10094 874 10128 908
rect 10094 806 10128 835
rect 10094 738 10128 760
rect 10094 670 10128 685
rect 10094 602 10128 610
rect 10094 534 10128 535
rect 10094 494 10128 500
rect 10094 419 10128 432
rect 10094 344 10128 364
rect 10094 269 10128 296
rect 10094 194 10128 228
rect 10094 144 10128 160
rect 10310 1078 10344 1094
rect 10310 1010 10344 1044
rect 10310 942 10344 974
rect 10310 874 10344 900
rect 10310 806 10344 826
rect 10310 738 10344 752
rect 10310 670 10344 678
rect 10310 602 10344 604
rect 10310 564 10344 568
rect 10310 490 10344 500
rect 10310 416 10344 432
rect 10310 342 10344 364
rect 10310 268 10344 296
rect 10310 194 10344 228
rect 10310 144 10344 160
rect 10526 1019 10560 1044
rect 10526 944 10560 976
rect 10526 874 10560 908
rect 10526 806 10560 835
rect 10526 738 10560 760
rect 10526 670 10560 685
rect 10526 602 10560 610
rect 10526 534 10560 535
rect 10526 494 10560 500
rect 10526 419 10560 432
rect 10526 344 10560 364
rect 10526 269 10560 296
rect 10526 194 10560 228
rect 10526 144 10560 160
rect 10742 1078 10776 1094
rect 10742 1010 10776 1044
rect 10742 942 10776 974
rect 10742 874 10776 900
rect 10742 806 10776 826
rect 10742 738 10776 752
rect 10742 670 10776 678
rect 10742 602 10776 604
rect 10742 564 10776 568
rect 10742 490 10776 500
rect 10742 416 10776 432
rect 10742 342 10776 364
rect 10742 268 10776 296
rect 10742 194 10776 228
rect 10742 144 10776 160
rect 10958 1019 10992 1044
rect 10958 944 10992 976
rect 10958 874 10992 908
rect 10958 806 10992 835
rect 10958 738 10992 760
rect 10958 670 10992 685
rect 10958 602 10992 610
rect 10958 534 10992 535
rect 10958 494 10992 500
rect 10958 419 10992 432
rect 10958 344 10992 364
rect 10958 269 10992 296
rect 10958 194 10992 228
rect 10958 144 10992 160
rect 11174 1078 11208 1094
rect 11174 1010 11208 1044
rect 11174 942 11208 974
rect 11174 874 11208 900
rect 11174 806 11208 826
rect 11174 738 11208 752
rect 11174 670 11208 678
rect 11174 602 11208 604
rect 11174 564 11208 568
rect 11174 490 11208 500
rect 11174 416 11208 432
rect 11174 342 11208 364
rect 11174 268 11208 296
rect 11174 194 11208 228
rect 11174 144 11208 160
rect 11390 1019 11424 1044
rect 11390 944 11424 976
rect 11390 874 11424 908
rect 11390 806 11424 835
rect 11390 738 11424 760
rect 11390 670 11424 685
rect 11390 602 11424 610
rect 11390 534 11424 535
rect 11390 494 11424 500
rect 11390 419 11424 432
rect 11390 344 11424 364
rect 11390 269 11424 296
rect 11390 194 11424 228
rect 11390 144 11424 160
rect 11606 1078 11640 1094
rect 11606 1010 11640 1044
rect 11606 942 11640 974
rect 11606 874 11640 900
rect 11606 806 11640 826
rect 11606 738 11640 752
rect 11606 670 11640 678
rect 11606 602 11640 604
rect 11606 564 11640 568
rect 11606 490 11640 500
rect 11606 416 11640 432
rect 11606 342 11640 364
rect 11606 268 11640 296
rect 11606 194 11640 228
rect 11606 144 11640 160
rect 11822 1078 11823 1094
rect 11856 1044 11857 1060
rect 11822 1019 11857 1044
rect 11822 1010 11823 1019
rect 11856 976 11857 985
rect 11822 944 11857 976
rect 11822 942 11823 944
rect 11856 908 11857 910
rect 11822 874 11857 908
rect 11856 869 11857 874
rect 11822 835 11823 840
rect 11822 806 11857 835
rect 11856 794 11857 806
rect 11822 760 11823 772
rect 11822 738 11857 760
rect 11856 719 11857 738
rect 11822 685 11823 704
rect 11822 670 11857 685
rect 11856 644 11857 670
rect 11822 610 11823 636
rect 11822 602 11857 610
rect 11856 569 11857 602
rect 11822 535 11823 568
rect 11822 534 11857 535
rect 11856 500 11857 534
rect 11822 494 11857 500
rect 11822 466 11823 494
rect 11856 432 11857 460
rect 11822 419 11857 432
rect 11822 398 11823 419
rect 11856 364 11857 385
rect 11822 344 11857 364
rect 11822 330 11823 344
rect 11856 296 11857 310
rect 11822 269 11857 296
rect 11822 262 11823 269
rect 11856 228 11857 235
rect 11822 194 11857 228
rect 12038 1078 12072 1094
rect 12038 1010 12072 1044
rect 12038 942 12072 974
rect 12038 874 12072 900
rect 12038 806 12072 826
rect 12038 738 12072 752
rect 12038 670 12072 678
rect 12038 602 12072 604
rect 12038 564 12072 568
rect 12038 490 12072 500
rect 12038 416 12072 432
rect 12038 342 12072 364
rect 12038 268 12072 296
rect 12038 194 12072 228
rect 11822 144 11856 160
rect 12038 144 12072 160
rect 12254 1019 12288 1044
rect 12254 944 12288 976
rect 12254 874 12288 908
rect 12254 806 12288 835
rect 12254 738 12288 760
rect 12254 670 12288 685
rect 12254 602 12288 610
rect 12254 534 12288 535
rect 12254 494 12288 500
rect 12254 419 12288 432
rect 12254 344 12288 364
rect 12254 269 12288 296
rect 12254 194 12288 228
rect 12254 144 12288 160
rect 12470 1078 12504 1094
rect 12470 1010 12504 1044
rect 12470 942 12504 974
rect 12470 874 12504 900
rect 12470 806 12504 826
rect 12470 738 12504 752
rect 12470 670 12504 678
rect 12470 602 12504 604
rect 12470 564 12504 568
rect 12470 490 12504 500
rect 12470 416 12504 432
rect 12470 342 12504 364
rect 12470 268 12504 296
rect 12470 194 12504 228
rect 12470 144 12504 160
rect 12686 1078 12720 1094
rect 12686 1010 12720 1044
rect 12686 942 12720 974
rect 12686 874 12720 900
rect 12686 806 12720 826
rect 12686 738 12720 752
rect 12686 670 12720 678
rect 12686 602 12720 604
rect 12686 564 12720 568
rect 12686 490 12720 500
rect 12686 416 12720 432
rect 12686 342 12720 364
rect 12686 268 12720 296
rect 12686 194 12720 228
rect 12686 144 12720 160
rect 12902 1078 12936 1094
rect 12902 1010 12936 1044
rect 12902 942 12936 974
rect 12902 874 12936 900
rect 12902 806 12936 826
rect 12902 738 12936 752
rect 12902 670 12936 678
rect 12902 602 12936 604
rect 12902 564 12936 568
rect 12902 490 12936 500
rect 12902 416 12936 432
rect 12902 342 12936 364
rect 12902 268 12936 296
rect 12902 194 12936 228
rect 12902 144 12936 160
rect 13118 1078 13152 1094
rect 13118 1010 13152 1044
rect 13118 942 13152 974
rect 13118 874 13152 900
rect 13118 806 13152 826
rect 13118 738 13152 752
rect 13118 670 13152 678
rect 13118 602 13152 604
rect 13118 564 13152 568
rect 13118 490 13152 500
rect 13118 416 13152 432
rect 13118 342 13152 364
rect 13118 268 13152 296
rect 13118 194 13152 228
rect 13118 144 13152 160
rect 13334 1078 13368 1094
rect 13334 1010 13368 1044
rect 13334 942 13368 974
rect 13334 874 13368 900
rect 13334 806 13368 826
rect 13334 738 13368 752
rect 13334 670 13368 678
rect 13334 602 13368 604
rect 13334 564 13368 568
rect 13334 490 13368 500
rect 13334 416 13368 432
rect 13334 342 13368 364
rect 13334 268 13368 296
rect 13334 194 13368 228
rect 13334 144 13368 160
rect 13550 1078 13584 1094
rect 13550 1010 13584 1044
rect 13550 942 13584 974
rect 13550 874 13584 900
rect 13550 806 13584 826
rect 13550 738 13584 752
rect 13550 670 13584 678
rect 13550 602 13584 604
rect 13550 564 13584 568
rect 13550 490 13584 500
rect 13550 416 13584 432
rect 13550 342 13584 364
rect 13550 268 13584 296
rect 13550 194 13584 228
rect 13550 144 13584 160
rect 13766 1078 13800 1094
rect 13766 1010 13800 1044
rect 13766 942 13800 974
rect 13766 874 13800 900
rect 13766 806 13800 826
rect 13766 738 13800 752
rect 13766 670 13800 678
rect 13766 602 13800 604
rect 13766 564 13800 568
rect 13766 490 13800 500
rect 13766 416 13800 432
rect 13766 342 13800 364
rect 13766 268 13800 296
rect 13766 194 13800 228
rect 13766 144 13800 160
rect 13982 1078 14016 1094
rect 13982 1010 14016 1044
rect 13982 942 14016 974
rect 13982 874 14016 900
rect 13982 806 14016 826
rect 13982 738 14016 752
rect 13982 670 14016 678
rect 13982 602 14016 604
rect 13982 564 14016 568
rect 13982 490 14016 500
rect 13982 416 14016 432
rect 13982 342 14016 364
rect 13982 268 14016 296
rect 13982 194 14016 228
rect 13982 144 14016 160
rect 14198 1078 14232 1094
rect 14198 1010 14232 1044
rect 14198 942 14232 974
rect 14198 874 14232 900
rect 14198 806 14232 826
rect 14198 738 14232 752
rect 14198 670 14232 678
rect 14198 602 14232 604
rect 14198 564 14232 568
rect 14198 490 14232 500
rect 14198 416 14232 432
rect 14198 342 14232 364
rect 14198 268 14232 296
rect 14198 194 14232 228
rect 14198 144 14232 160
rect 14414 1078 14448 1094
rect 14414 1010 14448 1044
rect 14414 942 14448 974
rect 14414 874 14448 900
rect 14414 806 14448 826
rect 14414 738 14448 752
rect 14414 670 14448 678
rect 14414 602 14448 604
rect 14414 564 14448 568
rect 14414 490 14448 500
rect 14414 416 14448 432
rect 14414 342 14448 364
rect 14414 268 14448 296
rect 14414 194 14448 228
rect 14414 144 14448 160
rect 14630 1078 14664 1094
rect 14630 1010 14664 1044
rect 14630 942 14664 974
rect 14630 874 14664 900
rect 14630 806 14664 826
rect 14630 738 14664 752
rect 14630 670 14664 678
rect 14630 602 14664 604
rect 14630 564 14664 568
rect 14630 490 14664 500
rect 14630 416 14664 432
rect 14630 342 14664 364
rect 14630 268 14664 296
rect 14630 194 14664 228
rect 14630 144 14664 160
rect 14846 1078 14880 1094
rect 14846 1010 14880 1044
rect 14846 942 14880 974
rect 14846 874 14880 900
rect 14846 806 14880 826
rect 14846 738 14880 752
rect 14846 670 14880 678
rect 14846 602 14880 604
rect 14846 564 14880 568
rect 14846 490 14880 500
rect 14846 416 14880 432
rect 14846 342 14880 364
rect 14846 268 14880 296
rect 14846 194 14880 228
rect 14846 144 14880 160
rect 15062 1078 15096 1094
rect 15062 1010 15096 1044
rect 15062 942 15096 974
rect 15062 874 15096 900
rect 15062 806 15096 826
rect 15062 738 15096 752
rect 15062 670 15096 678
rect 15062 602 15096 604
rect 15062 564 15096 568
rect 15172 1012 15206 1036
rect 15172 934 15206 968
rect 15172 866 15206 897
rect 15172 798 15206 816
rect 15172 730 15206 734
rect 15172 686 15206 696
rect 15172 604 15206 628
rect 15172 544 15206 560
rect 15428 1012 15462 1036
rect 15428 934 15462 968
rect 15428 866 15462 897
rect 15428 798 15462 816
rect 15428 730 15462 734
rect 15428 686 15462 696
rect 15428 604 15462 628
rect 15428 544 15462 560
rect 15538 1019 15572 1044
rect 15538 944 15572 976
rect 15538 874 15572 908
rect 15538 806 15572 835
rect 15538 738 15572 760
rect 15538 670 15572 685
rect 15538 602 15572 610
rect 15062 490 15096 500
rect 15062 416 15096 432
rect 15062 342 15096 364
rect 15062 268 15096 296
rect 15062 194 15096 228
rect 15062 144 15096 160
rect 15538 534 15572 535
rect 15538 494 15572 500
rect 15538 419 15572 432
rect 15538 344 15572 364
rect 15538 269 15572 296
rect 15538 194 15572 228
rect 15538 144 15572 160
rect 15754 1019 15788 1044
rect 15754 944 15788 976
rect 15754 874 15788 908
rect 15754 806 15788 835
rect 15754 738 15788 760
rect 15754 670 15788 685
rect 15754 602 15788 610
rect 15754 534 15788 535
rect 15754 494 15788 500
rect 15754 419 15788 432
rect 15754 344 15788 364
rect 15754 269 15788 296
rect 15754 194 15788 228
rect 15754 144 15788 160
rect 15970 1019 16004 1044
rect 15970 944 16004 976
rect 15970 874 16004 908
rect 15970 806 16004 835
rect 15970 738 16004 760
rect 15970 670 16004 685
rect 15970 602 16004 610
rect 15970 534 16004 535
rect 15970 494 16004 500
rect 15970 419 16004 432
rect 15970 344 16004 364
rect 15970 269 16004 296
rect 15970 194 16004 228
rect 15970 144 16004 160
rect 1499 48 1523 82
rect 1557 48 1597 82
rect 1656 48 1671 82
rect 1730 48 1745 82
rect 1804 48 1819 82
rect 1878 48 1893 82
rect 1952 48 1967 82
rect 2026 48 2040 82
rect 2100 48 2113 82
rect 2174 48 2186 82
rect 2248 48 2259 82
rect 2979 48 2991 82
rect 3037 48 3065 82
rect 3106 48 3139 82
rect 3175 48 3210 82
rect 3247 48 3279 82
rect 3322 48 3348 82
rect 3397 48 3406 82
rect 3934 40 3946 74
rect 3992 40 4020 74
rect 4062 40 4094 74
rect 4132 40 4168 74
rect 4202 40 4238 74
rect 4276 40 4308 74
rect 4350 40 4378 74
rect 4424 40 4448 74
rect 4498 40 4518 74
rect 4572 40 4587 74
rect 4646 40 4656 74
rect 4719 40 4725 74
rect 4792 40 4794 74
rect 4828 40 4831 74
rect 4897 40 4904 74
rect 4966 40 4977 74
rect 5035 40 5050 74
rect 5104 40 5123 74
rect 5173 40 5196 74
rect 5242 40 5269 74
rect 5311 40 5342 74
rect 5380 40 5415 74
rect 5449 40 5484 74
rect 5522 40 5553 74
rect 5595 40 5622 74
rect 5668 40 5680 74
rect 5923 74 5962 78
rect 5996 74 6035 78
rect 6069 74 6108 78
rect 6142 74 6181 78
rect 5923 44 5940 74
rect 5996 44 6009 74
rect 6069 44 6078 74
rect 6142 44 6147 74
rect 5916 40 5940 44
rect 5974 40 6009 44
rect 6043 40 6078 44
rect 6112 40 6147 44
rect 6215 74 6254 78
rect 6288 74 6327 78
rect 6361 74 6400 78
rect 6434 74 6473 78
rect 6507 74 6546 78
rect 6580 74 6619 78
rect 6653 74 6692 78
rect 6726 74 6765 78
rect 6799 74 6838 78
rect 6872 74 6911 78
rect 6945 74 6984 78
rect 7018 74 7057 78
rect 7091 74 7130 78
rect 7164 74 7203 78
rect 7237 74 7276 78
rect 7310 74 7349 78
rect 7383 74 7422 78
rect 7456 74 7495 78
rect 7529 74 7568 78
rect 7602 74 7641 78
rect 7675 74 7714 78
rect 7748 74 7787 78
rect 7821 74 7860 78
rect 7894 74 7933 78
rect 7967 74 8006 78
rect 8040 74 8079 78
rect 8113 74 8152 78
rect 8186 74 8225 78
rect 8259 74 8298 78
rect 8332 74 8371 78
rect 8405 74 8444 78
rect 8478 74 8517 78
rect 8551 74 8590 78
rect 8624 74 8663 78
rect 8697 74 8736 78
rect 8770 74 8809 78
rect 8843 74 8882 78
rect 8916 74 8955 78
rect 8989 74 9028 78
rect 9062 74 9101 78
rect 9135 74 9174 78
rect 6215 44 6216 74
rect 6181 40 6216 44
rect 6250 44 6254 74
rect 6318 44 6327 74
rect 6386 44 6400 74
rect 6454 44 6473 74
rect 6522 44 6546 74
rect 6590 44 6619 74
rect 6250 40 6284 44
rect 6318 40 6352 44
rect 6386 40 6420 44
rect 6454 40 6488 44
rect 6522 40 6556 44
rect 6590 40 6624 44
rect 6658 40 6692 74
rect 6726 40 6760 74
rect 6799 44 6828 74
rect 6872 44 6896 74
rect 6945 44 6964 74
rect 7018 44 7032 74
rect 7091 44 7100 74
rect 7164 44 7168 74
rect 6794 40 6828 44
rect 6862 40 6896 44
rect 6930 40 6964 44
rect 6998 40 7032 44
rect 7066 40 7100 44
rect 7134 40 7168 44
rect 7202 44 7203 74
rect 7270 44 7276 74
rect 7338 44 7349 74
rect 7406 44 7422 74
rect 7474 44 7495 74
rect 7542 44 7568 74
rect 7610 44 7641 74
rect 7202 40 7236 44
rect 7270 40 7304 44
rect 7338 40 7372 44
rect 7406 40 7440 44
rect 7474 40 7508 44
rect 7542 40 7576 44
rect 7610 40 7644 44
rect 7678 40 7712 74
rect 7748 44 7780 74
rect 7821 44 7848 74
rect 7894 44 7916 74
rect 7967 44 7984 74
rect 8040 44 8052 74
rect 8113 44 8120 74
rect 8186 44 8188 74
rect 7746 40 7780 44
rect 7814 40 7848 44
rect 7882 40 7916 44
rect 7950 40 7984 44
rect 8018 40 8052 44
rect 8086 40 8120 44
rect 8154 40 8188 44
rect 8222 44 8225 74
rect 8290 44 8298 74
rect 8358 44 8371 74
rect 8426 44 8444 74
rect 8494 44 8517 74
rect 8562 44 8590 74
rect 8630 44 8663 74
rect 8222 40 8256 44
rect 8290 40 8324 44
rect 8358 40 8392 44
rect 8426 40 8460 44
rect 8494 40 8528 44
rect 8562 40 8596 44
rect 8630 40 8664 44
rect 8698 40 8732 74
rect 8770 44 8800 74
rect 8843 44 8868 74
rect 8916 44 8936 74
rect 8989 44 9004 74
rect 9062 44 9072 74
rect 9135 44 9140 74
rect 8766 40 8800 44
rect 8834 40 8868 44
rect 8902 40 8936 44
rect 8970 40 9004 44
rect 9038 40 9072 44
rect 9106 40 9140 44
rect 9208 74 9247 78
rect 9281 74 9320 78
rect 9354 74 9393 78
rect 9427 74 9466 78
rect 9500 74 9539 78
rect 9573 74 9612 78
rect 9646 74 9685 78
rect 9719 74 9758 78
rect 9792 74 9831 78
rect 9865 74 9903 78
rect 9937 74 9975 78
rect 10009 74 10047 78
rect 10081 74 10119 78
rect 10153 74 10191 78
rect 10225 74 10263 78
rect 10297 74 10335 78
rect 10369 74 10407 78
rect 10441 74 10479 78
rect 10513 74 10551 78
rect 10585 74 10623 78
rect 10657 74 10695 78
rect 10729 74 10767 78
rect 10801 74 10839 78
rect 10873 74 10911 78
rect 10945 74 10983 78
rect 11017 74 11055 78
rect 11089 74 11127 78
rect 11161 74 11199 78
rect 11233 74 11271 78
rect 11305 74 11343 78
rect 11377 74 11415 78
rect 11449 74 11487 78
rect 11521 74 11559 78
rect 11593 74 11631 78
rect 11665 74 11703 78
rect 11737 74 11775 78
rect 11809 74 11847 78
rect 11881 74 11919 78
rect 11953 74 11991 78
rect 12025 74 12063 78
rect 12097 74 12135 78
rect 12169 74 12207 78
rect 12241 74 12279 78
rect 12313 74 12351 78
rect 12385 74 12423 78
rect 12457 74 12495 78
rect 12529 74 12567 78
rect 12601 74 12639 78
rect 12673 74 12711 78
rect 12745 74 12783 78
rect 12817 74 12855 78
rect 12889 74 12927 78
rect 12961 74 12999 78
rect 13033 74 13071 78
rect 13105 74 13143 78
rect 13177 74 13215 78
rect 13249 74 13287 78
rect 13321 74 13359 78
rect 13393 74 13431 78
rect 13465 74 13503 78
rect 13537 74 13575 78
rect 13609 74 13647 78
rect 13681 74 13719 78
rect 13753 74 13791 78
rect 13825 74 13863 78
rect 13897 74 13935 78
rect 13969 74 14007 78
rect 14041 74 14079 78
rect 14113 74 14151 78
rect 14185 74 14223 78
rect 14257 74 14295 78
rect 14329 74 14367 78
rect 14401 74 14439 78
rect 14473 74 14511 78
rect 14545 74 14583 78
rect 14617 74 14655 78
rect 14689 74 14727 78
rect 14761 74 14799 78
rect 14833 74 14871 78
rect 14905 74 14943 78
rect 14977 74 15015 78
rect 15049 74 15087 78
rect 15121 74 15159 78
rect 15193 74 15231 78
rect 15265 74 15303 78
rect 15337 74 15375 78
rect 15409 74 15447 78
rect 15481 74 15519 78
rect 15553 74 15591 78
rect 15625 74 15663 78
rect 15697 74 15735 78
rect 15769 74 15807 78
rect 15841 74 15879 78
rect 15913 74 15951 78
rect 9174 40 9208 44
rect 9242 44 9247 74
rect 9310 44 9320 74
rect 9378 44 9393 74
rect 9446 44 9466 74
rect 9514 44 9539 74
rect 9582 44 9612 74
rect 9242 40 9276 44
rect 9310 40 9344 44
rect 9378 40 9412 44
rect 9446 40 9480 44
rect 9514 40 9548 44
rect 9582 40 9616 44
rect 9650 40 9684 74
rect 9719 44 9752 74
rect 9792 44 9820 74
rect 9865 44 9888 74
rect 9937 44 9956 74
rect 10009 44 10024 74
rect 10081 44 10092 74
rect 10153 44 10160 74
rect 10225 44 10228 74
rect 9718 40 9752 44
rect 9786 40 9820 44
rect 9854 40 9888 44
rect 9922 40 9956 44
rect 9990 40 10024 44
rect 10058 40 10092 44
rect 10126 40 10160 44
rect 10194 40 10228 44
rect 10262 44 10263 74
rect 10330 44 10335 74
rect 10398 44 10407 74
rect 10466 44 10479 74
rect 10534 44 10551 74
rect 10602 44 10623 74
rect 10670 44 10695 74
rect 10738 44 10767 74
rect 10806 44 10839 74
rect 10262 40 10296 44
rect 10330 40 10364 44
rect 10398 40 10432 44
rect 10466 40 10500 44
rect 10534 40 10568 44
rect 10602 40 10636 44
rect 10670 40 10704 44
rect 10738 40 10772 44
rect 10806 40 10840 44
rect 10874 40 10908 74
rect 10945 44 10976 74
rect 11017 44 11044 74
rect 11089 44 11112 74
rect 11161 44 11180 74
rect 11233 44 11248 74
rect 11305 44 11316 74
rect 11377 44 11384 74
rect 11449 44 11452 74
rect 10942 40 10976 44
rect 11010 40 11044 44
rect 11078 40 11112 44
rect 11146 40 11180 44
rect 11214 40 11248 44
rect 11282 40 11316 44
rect 11350 40 11384 44
rect 11418 40 11452 44
rect 11486 44 11487 74
rect 11554 44 11559 74
rect 11622 44 11631 74
rect 11690 44 11703 74
rect 11758 44 11775 74
rect 11826 44 11847 74
rect 11894 44 11919 74
rect 11962 44 11991 74
rect 12030 44 12063 74
rect 11486 40 11520 44
rect 11554 40 11588 44
rect 11622 40 11656 44
rect 11690 40 11724 44
rect 11758 40 11792 44
rect 11826 40 11860 44
rect 11894 40 11928 44
rect 11962 40 11996 44
rect 12030 40 12064 44
rect 12098 40 12132 74
rect 12169 44 12200 74
rect 12241 44 12268 74
rect 12313 44 12336 74
rect 12385 44 12404 74
rect 12457 44 12472 74
rect 12529 44 12540 74
rect 12601 44 12608 74
rect 12673 44 12676 74
rect 12166 40 12200 44
rect 12234 40 12268 44
rect 12302 40 12336 44
rect 12370 40 12404 44
rect 12438 40 12472 44
rect 12506 40 12540 44
rect 12574 40 12608 44
rect 12642 40 12676 44
rect 12710 44 12711 74
rect 12778 44 12783 74
rect 12846 44 12855 74
rect 12914 44 12927 74
rect 12982 44 12999 74
rect 13050 44 13071 74
rect 13118 44 13143 74
rect 13186 44 13215 74
rect 13254 44 13287 74
rect 12710 40 12744 44
rect 12778 40 12812 44
rect 12846 40 12880 44
rect 12914 40 12948 44
rect 12982 40 13016 44
rect 13050 40 13084 44
rect 13118 40 13152 44
rect 13186 40 13220 44
rect 13254 40 13288 44
rect 13322 40 13356 74
rect 13393 44 13424 74
rect 13465 44 13492 74
rect 13537 44 13560 74
rect 13609 44 13628 74
rect 13681 44 13696 74
rect 13753 44 13764 74
rect 13825 44 13832 74
rect 13897 44 13900 74
rect 13390 40 13424 44
rect 13458 40 13492 44
rect 13526 40 13560 44
rect 13594 40 13628 44
rect 13662 40 13696 44
rect 13730 40 13764 44
rect 13798 40 13832 44
rect 13866 40 13900 44
rect 13934 44 13935 74
rect 14002 44 14007 74
rect 14070 44 14079 74
rect 14138 44 14151 74
rect 14206 44 14223 74
rect 14274 44 14295 74
rect 14342 44 14367 74
rect 14410 44 14439 74
rect 14478 44 14511 74
rect 13934 40 13968 44
rect 14002 40 14036 44
rect 14070 40 14104 44
rect 14138 40 14172 44
rect 14206 40 14240 44
rect 14274 40 14308 44
rect 14342 40 14376 44
rect 14410 40 14444 44
rect 14478 40 14512 44
rect 14546 40 14580 74
rect 14617 44 14648 74
rect 14689 44 14716 74
rect 14761 44 14784 74
rect 14833 44 14852 74
rect 14905 44 14920 74
rect 14977 44 14988 74
rect 15049 44 15056 74
rect 15121 44 15124 74
rect 14614 40 14648 44
rect 14682 40 14716 44
rect 14750 40 14784 44
rect 14818 40 14852 44
rect 14886 40 14920 44
rect 14954 40 14988 44
rect 15022 40 15056 44
rect 15090 40 15124 44
rect 15158 44 15159 74
rect 15226 44 15231 74
rect 15294 44 15303 74
rect 15362 44 15375 74
rect 15430 44 15447 74
rect 15498 44 15519 74
rect 15566 44 15591 74
rect 15634 44 15663 74
rect 15702 44 15735 74
rect 15158 40 15192 44
rect 15226 40 15260 44
rect 15294 40 15328 44
rect 15362 40 15396 44
rect 15430 40 15464 44
rect 15498 40 15532 44
rect 15566 40 15600 44
rect 15634 40 15668 44
rect 15702 40 15736 44
rect 15770 40 15804 74
rect 15841 44 15872 74
rect 15913 44 15940 74
rect 15985 44 15998 74
rect 15838 40 15872 44
rect 15906 40 15940 44
rect 15974 40 15998 44
<< viali >>
rect 292 3238 312 3272
rect 312 3238 326 3272
rect 374 3238 380 3272
rect 380 3238 408 3272
rect 456 3238 482 3272
rect 482 3238 490 3272
rect 538 3238 550 3272
rect 550 3238 572 3272
rect 648 3238 652 3272
rect 652 3238 682 3272
rect 720 3238 754 3272
rect 792 3238 822 3272
rect 822 3238 826 3272
rect 864 3238 890 3272
rect 890 3238 898 3272
rect 936 3238 958 3272
rect 958 3238 970 3272
rect 1008 3238 1026 3272
rect 1026 3238 1042 3272
rect 1080 3238 1094 3272
rect 1094 3238 1114 3272
rect 1152 3238 1162 3272
rect 1162 3238 1186 3272
rect 1224 3238 1230 3272
rect 1230 3238 1258 3272
rect 1296 3238 1298 3272
rect 1298 3238 1330 3272
rect 1368 3238 1400 3272
rect 1400 3238 1402 3272
rect 1440 3238 1468 3272
rect 1468 3238 1474 3272
rect 1512 3238 1536 3272
rect 1536 3238 1546 3272
rect 1584 3238 1604 3272
rect 1604 3238 1618 3272
rect 1656 3238 1672 3272
rect 1672 3238 1690 3272
rect 1728 3238 1740 3272
rect 1740 3238 1762 3272
rect 1800 3238 1808 3272
rect 1808 3238 1834 3272
rect 1872 3238 1876 3272
rect 1876 3238 1906 3272
rect 1944 3238 1978 3272
rect 2016 3238 2046 3272
rect 2046 3238 2050 3272
rect 2088 3238 2114 3272
rect 2114 3238 2122 3272
rect 2160 3238 2182 3272
rect 2182 3238 2194 3272
rect 2232 3238 2250 3272
rect 2250 3238 2266 3272
rect 2304 3238 2318 3272
rect 2318 3238 2338 3272
rect 2376 3238 2386 3272
rect 2386 3238 2410 3272
rect 2448 3238 2454 3272
rect 2454 3238 2482 3272
rect 2520 3238 2522 3272
rect 2522 3238 2554 3272
rect 2592 3238 2624 3272
rect 2624 3238 2626 3272
rect 2664 3238 2692 3272
rect 2692 3238 2698 3272
rect 2736 3238 2760 3272
rect 2760 3238 2770 3272
rect 2808 3238 2828 3272
rect 2828 3238 2842 3272
rect 2880 3238 2896 3272
rect 2896 3238 2914 3272
rect 2952 3238 2964 3272
rect 2964 3238 2986 3272
rect 3024 3238 3032 3272
rect 3032 3238 3058 3272
rect 3096 3238 3100 3272
rect 3100 3238 3130 3272
rect 3168 3238 3202 3272
rect 3240 3238 3270 3272
rect 3270 3238 3274 3272
rect 3312 3238 3338 3272
rect 3338 3238 3346 3272
rect 3384 3238 3406 3272
rect 3406 3238 3418 3272
rect 3456 3238 3474 3272
rect 3474 3238 3490 3272
rect 3528 3238 3542 3272
rect 3542 3238 3562 3272
rect 3600 3238 3610 3272
rect 3610 3238 3634 3272
rect 3672 3238 3678 3272
rect 3678 3238 3706 3272
rect 3744 3238 3746 3272
rect 3746 3238 3778 3272
rect 3816 3238 3848 3272
rect 3848 3238 3850 3272
rect 3888 3238 3916 3272
rect 3916 3238 3922 3272
rect 3960 3238 3984 3272
rect 3984 3238 3994 3272
rect 4032 3238 4052 3272
rect 4052 3238 4066 3272
rect 4104 3238 4120 3272
rect 4120 3238 4138 3272
rect 4176 3238 4188 3272
rect 4188 3238 4210 3272
rect 4248 3238 4256 3272
rect 4256 3238 4282 3272
rect 4320 3238 4324 3272
rect 4324 3238 4354 3272
rect 4392 3238 4426 3272
rect 4464 3238 4494 3272
rect 4494 3238 4498 3272
rect 4536 3238 4562 3272
rect 4562 3238 4570 3272
rect 4608 3238 4630 3272
rect 4630 3238 4642 3272
rect 4680 3238 4698 3272
rect 4698 3238 4714 3272
rect 4752 3238 4766 3272
rect 4766 3238 4786 3272
rect 4824 3238 4858 3272
rect 210 3191 244 3200
rect 210 3166 244 3191
rect 210 3089 244 3113
rect 210 3079 244 3089
rect 4896 3170 4930 3198
rect 4896 3164 4930 3170
rect 4896 3102 4930 3124
rect 4896 3090 4930 3102
rect 210 3021 244 3026
rect 210 2992 244 3021
rect 210 2919 244 2939
rect 210 2905 244 2919
rect 505 3015 535 3049
rect 535 3015 539 3049
rect 577 3015 603 3049
rect 603 3015 611 3049
rect 649 3015 671 3049
rect 671 3015 683 3049
rect 721 3015 739 3049
rect 739 3015 755 3049
rect 794 3015 807 3049
rect 807 3015 828 3049
rect 867 3015 875 3049
rect 875 3015 901 3049
rect 940 3015 943 3049
rect 943 3015 974 3049
rect 1013 3015 1045 3049
rect 1045 3015 1047 3049
rect 1086 3015 1113 3049
rect 1113 3015 1120 3049
rect 1159 3015 1181 3049
rect 1181 3015 1193 3049
rect 1232 3015 1249 3049
rect 1249 3015 1266 3049
rect 1305 3015 1317 3049
rect 1317 3015 1339 3049
rect 1378 3015 1385 3049
rect 1385 3015 1412 3049
rect 1451 3015 1453 3049
rect 1453 3015 1485 3049
rect 1524 3015 1555 3049
rect 1555 3015 1558 3049
rect 1597 3015 1623 3049
rect 1623 3015 1631 3049
rect 1670 3015 1691 3049
rect 1691 3015 1704 3049
rect 1743 3015 1759 3049
rect 1759 3015 1777 3049
rect 1816 3015 1827 3049
rect 1827 3015 1850 3049
rect 1889 3015 1895 3049
rect 1895 3015 1923 3049
rect 1962 3015 1963 3049
rect 1963 3015 1996 3049
rect 2035 3015 2065 3049
rect 2065 3015 2069 3049
rect 2108 3015 2133 3049
rect 2133 3015 2142 3049
rect 2181 3015 2201 3049
rect 2201 3015 2215 3049
rect 2254 3015 2269 3049
rect 2269 3015 2288 3049
rect 2327 3015 2337 3049
rect 2337 3015 2361 3049
rect 2400 3015 2405 3049
rect 2405 3015 2434 3049
rect 2473 3015 2507 3049
rect 2546 3015 2575 3049
rect 2575 3015 2580 3049
rect 2619 3015 2643 3049
rect 2643 3015 2653 3049
rect 2692 3015 2711 3049
rect 2711 3015 2726 3049
rect 2765 3015 2779 3049
rect 2779 3015 2799 3049
rect 2838 3015 2847 3049
rect 2847 3015 2872 3049
rect 2911 3015 2915 3049
rect 2915 3015 2945 3049
rect 2984 3015 3017 3049
rect 3017 3015 3018 3049
rect 3057 3015 3085 3049
rect 3085 3015 3091 3049
rect 3130 3015 3153 3049
rect 3153 3015 3164 3049
rect 3203 3015 3221 3049
rect 3221 3015 3237 3049
rect 3276 3015 3289 3049
rect 3289 3015 3310 3049
rect 3349 3015 3357 3049
rect 3357 3015 3383 3049
rect 3422 3015 3425 3049
rect 3425 3015 3456 3049
rect 3495 3015 3527 3049
rect 3527 3015 3529 3049
rect 3568 3015 3595 3049
rect 3595 3015 3602 3049
rect 3678 3015 3697 3049
rect 3697 3015 3712 3049
rect 3754 3015 3765 3049
rect 3765 3015 3788 3049
rect 3831 3015 3833 3049
rect 3833 3015 3865 3049
rect 3908 3015 3935 3049
rect 3935 3015 3942 3049
rect 3985 3015 4003 3049
rect 4003 3015 4019 3049
rect 4062 3015 4071 3049
rect 4071 3015 4096 3049
rect 4139 3015 4173 3049
rect 4216 3015 4241 3049
rect 4241 3015 4250 3049
rect 4293 3015 4309 3049
rect 4309 3015 4327 3049
rect 4370 3015 4377 3049
rect 4377 3015 4404 3049
rect 4447 3015 4479 3049
rect 4479 3015 4481 3049
rect 4524 3015 4547 3049
rect 4547 3015 4558 3049
rect 4601 3015 4615 3049
rect 4615 3015 4635 3049
rect 433 2943 467 2977
rect 433 2870 467 2902
rect 433 2868 467 2870
rect 4673 2947 4707 2975
rect 4673 2941 4707 2947
rect 4673 2879 4707 2901
rect 4673 2867 4707 2879
rect -101 2760 -67 2764
rect -101 2730 -67 2760
rect -101 2658 -67 2684
rect -101 2650 -67 2658
rect -101 2590 -67 2604
rect -101 2570 -67 2590
rect -101 2522 -67 2523
rect -101 2489 -67 2522
rect -101 2420 -67 2442
rect -101 2408 -67 2420
rect -101 2352 -67 2361
rect -101 2327 -67 2352
rect -101 2250 -67 2280
rect -101 2246 -67 2250
rect 55 2760 89 2764
rect 55 2730 89 2760
rect 55 2658 89 2684
rect 55 2650 89 2658
rect 55 2590 89 2604
rect 55 2570 89 2590
rect 55 2522 89 2523
rect 55 2489 89 2522
rect 55 2420 89 2442
rect 55 2408 89 2420
rect 55 2352 89 2361
rect 55 2327 89 2352
rect 55 2250 89 2280
rect 55 2246 89 2250
rect 199 2749 210 2780
rect 210 2749 233 2780
rect 199 2746 233 2749
rect 199 2681 210 2705
rect 210 2681 233 2705
rect 199 2671 233 2681
rect 199 2613 210 2630
rect 210 2613 233 2630
rect 199 2596 233 2613
rect 199 2545 210 2555
rect 210 2545 233 2555
rect 199 2521 233 2545
rect 199 2477 210 2480
rect 210 2477 233 2480
rect 199 2446 233 2477
rect 199 2375 233 2405
rect 199 2371 210 2375
rect 210 2371 233 2375
rect 199 2307 233 2330
rect 199 2296 210 2307
rect 210 2296 233 2307
rect 199 2239 233 2255
rect 199 2221 210 2239
rect 210 2221 233 2239
rect -59 2156 -55 2190
rect -55 2156 -25 2190
rect 13 2156 47 2190
rect 199 2171 233 2180
rect 199 2146 210 2171
rect 210 2146 233 2171
rect 199 2103 233 2106
rect 199 2072 210 2103
rect 210 2072 233 2103
rect 199 2001 210 2032
rect 210 2001 233 2032
rect 199 1998 233 2001
rect 199 1933 210 1958
rect 210 1933 233 1958
rect 199 1924 233 1933
rect 433 2802 467 2827
rect 433 2793 467 2802
rect 433 2734 467 2752
rect 433 2718 467 2734
rect 433 2666 467 2677
rect 433 2643 467 2666
rect 433 2598 467 2602
rect 433 2568 467 2598
rect 433 2496 467 2528
rect 433 2494 467 2496
rect 433 2428 467 2454
rect 433 2420 467 2428
rect 433 2360 467 2380
rect 433 2346 467 2360
rect 433 2292 467 2306
rect 433 2272 467 2292
rect 433 2224 467 2232
rect 433 2198 467 2224
rect 433 2156 467 2158
rect 433 2124 467 2156
rect 433 2054 467 2084
rect 433 2050 467 2054
rect 433 1986 467 2010
rect 433 1976 467 1986
rect 210 1797 244 1812
rect 210 1778 244 1797
rect 210 1729 244 1735
rect 210 1701 244 1729
rect 433 1918 467 1936
rect 433 1902 467 1918
rect 720 2851 754 2867
rect 720 2833 754 2851
rect 720 2783 754 2788
rect 720 2754 754 2783
rect 720 2681 754 2709
rect 720 2675 754 2681
rect 720 2613 754 2630
rect 720 2596 754 2613
rect 720 2545 754 2551
rect 720 2517 754 2545
rect 720 2443 754 2472
rect 720 2438 754 2443
rect 720 2375 754 2393
rect 720 2359 754 2375
rect 720 2307 754 2314
rect 720 2280 754 2307
rect 720 2205 754 2234
rect 720 2200 754 2205
rect 720 2137 754 2154
rect 720 2120 754 2137
rect 876 2851 910 2867
rect 876 2833 910 2851
rect 876 2783 910 2792
rect 876 2758 910 2783
rect 876 2715 910 2717
rect 876 2683 910 2715
rect 876 2613 910 2642
rect 876 2608 910 2613
rect 876 2545 910 2567
rect 876 2533 910 2545
rect 876 2477 910 2492
rect 876 2458 910 2477
rect 876 2409 910 2417
rect 876 2383 910 2409
rect 876 2341 910 2342
rect 876 2308 910 2341
rect 876 2239 910 2267
rect 876 2233 910 2239
rect 876 2171 910 2192
rect 876 2158 910 2171
rect 876 2103 910 2117
rect 876 2083 910 2103
rect 876 2035 910 2042
rect 876 2008 910 2035
rect 876 1933 910 1967
rect 1032 2851 1066 2867
rect 1032 2833 1066 2851
rect 1032 2783 1066 2792
rect 1032 2758 1066 2783
rect 1032 2715 1066 2717
rect 1032 2683 1066 2715
rect 1032 2613 1066 2642
rect 1032 2608 1066 2613
rect 1032 2545 1066 2567
rect 1032 2533 1066 2545
rect 1032 2477 1066 2492
rect 1032 2458 1066 2477
rect 1032 2409 1066 2417
rect 1032 2383 1066 2409
rect 1032 2341 1066 2342
rect 1032 2308 1066 2341
rect 1032 2239 1066 2267
rect 1032 2233 1066 2239
rect 1032 2171 1066 2192
rect 1032 2158 1066 2171
rect 1032 2103 1066 2117
rect 1032 2083 1066 2103
rect 1032 2035 1066 2042
rect 1032 2008 1066 2035
rect 1032 1933 1066 1967
rect 1142 2851 1176 2867
rect 1142 2833 1176 2851
rect 1142 2783 1176 2792
rect 1142 2758 1176 2783
rect 1142 2715 1176 2717
rect 1142 2683 1176 2715
rect 1142 2613 1176 2642
rect 1142 2608 1176 2613
rect 1142 2545 1176 2567
rect 1142 2533 1176 2545
rect 1142 2477 1176 2492
rect 1142 2458 1176 2477
rect 1142 2409 1176 2417
rect 1142 2383 1176 2409
rect 1142 2341 1176 2342
rect 1142 2308 1176 2341
rect 1142 2239 1176 2267
rect 1142 2233 1176 2239
rect 1142 2171 1176 2192
rect 1142 2158 1176 2171
rect 1142 2103 1176 2117
rect 1142 2083 1176 2103
rect 1142 2035 1176 2042
rect 1142 2008 1176 2035
rect 1142 1933 1176 1967
rect 1298 2851 1332 2867
rect 1298 2833 1332 2851
rect 1298 2783 1332 2792
rect 1298 2758 1332 2783
rect 1298 2715 1332 2717
rect 1298 2683 1332 2715
rect 1298 2613 1332 2642
rect 1298 2608 1332 2613
rect 1298 2545 1332 2567
rect 1298 2533 1332 2545
rect 1298 2477 1332 2492
rect 1298 2458 1332 2477
rect 1298 2409 1332 2417
rect 1298 2383 1332 2409
rect 1298 2341 1332 2342
rect 1298 2308 1332 2341
rect 1298 2239 1332 2267
rect 1298 2233 1332 2239
rect 1298 2171 1332 2192
rect 1298 2158 1332 2171
rect 1298 2103 1332 2117
rect 1298 2083 1332 2103
rect 1298 2035 1332 2042
rect 1298 2008 1332 2035
rect 1298 1933 1332 1967
rect 1454 2851 1488 2867
rect 1454 2833 1488 2851
rect 1454 2783 1488 2788
rect 1454 2754 1488 2783
rect 1454 2681 1488 2709
rect 1454 2675 1488 2681
rect 1454 2613 1488 2630
rect 1454 2596 1488 2613
rect 1454 2545 1488 2551
rect 1454 2517 1488 2545
rect 1454 2443 1488 2472
rect 1454 2438 1488 2443
rect 1454 2375 1488 2393
rect 1454 2359 1488 2375
rect 1454 2307 1488 2314
rect 1454 2280 1488 2307
rect 1454 2205 1488 2234
rect 1454 2200 1488 2205
rect 1454 2137 1488 2154
rect 1454 2120 1488 2137
rect 1610 2851 1644 2867
rect 1610 2833 1644 2851
rect 1610 2783 1644 2792
rect 1610 2758 1644 2783
rect 1610 2715 1644 2717
rect 1610 2683 1644 2715
rect 1610 2613 1644 2642
rect 1610 2608 1644 2613
rect 1610 2545 1644 2567
rect 1610 2533 1644 2545
rect 1610 2477 1644 2492
rect 1610 2458 1644 2477
rect 1610 2409 1644 2417
rect 1610 2383 1644 2409
rect 1610 2341 1644 2342
rect 1610 2308 1644 2341
rect 1610 2239 1644 2267
rect 1610 2233 1644 2239
rect 1610 2171 1644 2192
rect 1610 2158 1644 2171
rect 1610 2103 1644 2117
rect 1610 2083 1644 2103
rect 1610 2035 1644 2042
rect 1610 2008 1644 2035
rect 1610 1933 1644 1967
rect 1766 2851 1800 2867
rect 1766 2833 1800 2851
rect 1766 2783 1800 2788
rect 1766 2754 1800 2783
rect 1766 2681 1800 2709
rect 1766 2675 1800 2681
rect 1766 2613 1800 2630
rect 1766 2596 1800 2613
rect 1766 2545 1800 2551
rect 1766 2517 1800 2545
rect 1766 2443 1800 2472
rect 1766 2438 1800 2443
rect 1766 2375 1800 2393
rect 1766 2359 1800 2375
rect 1766 2307 1800 2314
rect 1766 2280 1800 2307
rect 1766 2205 1800 2234
rect 1766 2200 1800 2205
rect 1766 2137 1800 2154
rect 1766 2120 1800 2137
rect 1922 2851 1956 2867
rect 1922 2833 1956 2851
rect 1922 2783 1956 2792
rect 1922 2758 1956 2783
rect 1922 2715 1956 2717
rect 1922 2683 1956 2715
rect 1922 2613 1956 2642
rect 1922 2608 1956 2613
rect 1922 2545 1956 2567
rect 1922 2533 1956 2545
rect 1922 2477 1956 2492
rect 1922 2458 1956 2477
rect 1922 2409 1956 2417
rect 1922 2383 1956 2409
rect 1922 2341 1956 2342
rect 1922 2308 1956 2341
rect 1922 2239 1956 2267
rect 1922 2233 1956 2239
rect 1922 2171 1956 2192
rect 1922 2158 1956 2171
rect 1922 2103 1956 2117
rect 1922 2083 1956 2103
rect 1922 2035 1956 2042
rect 1922 2008 1956 2035
rect 1922 1933 1956 1967
rect 2078 2851 2112 2867
rect 2078 2833 2112 2851
rect 2078 2783 2112 2792
rect 2078 2758 2112 2783
rect 2078 2715 2112 2717
rect 2078 2683 2112 2715
rect 2078 2613 2112 2642
rect 2078 2608 2112 2613
rect 2078 2545 2112 2567
rect 2078 2533 2112 2545
rect 2078 2477 2112 2492
rect 2078 2458 2112 2477
rect 2078 2409 2112 2417
rect 2078 2383 2112 2409
rect 2078 2341 2112 2342
rect 2078 2308 2112 2341
rect 2078 2239 2112 2267
rect 2078 2233 2112 2239
rect 2078 2171 2112 2192
rect 2078 2158 2112 2171
rect 2078 2103 2112 2117
rect 2078 2083 2112 2103
rect 2078 2035 2112 2042
rect 2078 2008 2112 2035
rect 2078 1933 2112 1967
rect 2234 2851 2268 2867
rect 2234 2833 2268 2851
rect 2234 2783 2268 2792
rect 2234 2758 2268 2783
rect 2234 2715 2268 2717
rect 2234 2683 2268 2715
rect 2234 2613 2268 2642
rect 2234 2608 2268 2613
rect 2234 2545 2268 2567
rect 2234 2533 2268 2545
rect 2234 2477 2268 2492
rect 2234 2458 2268 2477
rect 2234 2409 2268 2417
rect 2234 2383 2268 2409
rect 2234 2341 2268 2342
rect 2234 2308 2268 2341
rect 2234 2239 2268 2267
rect 2234 2233 2268 2239
rect 2234 2171 2268 2192
rect 2234 2158 2268 2171
rect 2234 2103 2268 2117
rect 2234 2083 2268 2103
rect 2234 2035 2268 2042
rect 2234 2008 2268 2035
rect 2234 1933 2268 1967
rect 2390 2851 2424 2867
rect 2390 2833 2424 2851
rect 2390 2783 2424 2792
rect 2390 2758 2424 2783
rect 2390 2715 2424 2717
rect 2390 2683 2424 2715
rect 2390 2613 2424 2642
rect 2390 2608 2424 2613
rect 2390 2545 2424 2567
rect 2390 2533 2424 2545
rect 2390 2477 2424 2492
rect 2390 2458 2424 2477
rect 2390 2409 2424 2417
rect 2390 2383 2424 2409
rect 2390 2341 2424 2342
rect 2390 2308 2424 2341
rect 2390 2239 2424 2267
rect 2390 2233 2424 2239
rect 2390 2171 2424 2192
rect 2390 2158 2424 2171
rect 2390 2103 2424 2117
rect 2390 2083 2424 2103
rect 2390 2035 2424 2042
rect 2390 2008 2424 2035
rect 2390 1933 2424 1967
rect 2546 2851 2580 2867
rect 2546 2833 2580 2851
rect 2546 2783 2580 2792
rect 2546 2758 2580 2783
rect 2546 2715 2580 2717
rect 2546 2683 2580 2715
rect 2546 2613 2580 2642
rect 2546 2608 2580 2613
rect 2546 2545 2580 2567
rect 2546 2533 2580 2545
rect 2546 2477 2580 2492
rect 2546 2458 2580 2477
rect 2546 2409 2580 2417
rect 2546 2383 2580 2409
rect 2546 2341 2580 2342
rect 2546 2308 2580 2341
rect 2546 2239 2580 2267
rect 2546 2233 2580 2239
rect 2546 2171 2580 2192
rect 2546 2158 2580 2171
rect 2546 2103 2580 2117
rect 2546 2083 2580 2103
rect 2546 2035 2580 2042
rect 2546 2008 2580 2035
rect 2546 1933 2580 1967
rect 2702 2851 2736 2867
rect 2702 2833 2736 2851
rect 2702 2783 2736 2792
rect 2702 2758 2736 2783
rect 2702 2715 2736 2717
rect 2702 2683 2736 2715
rect 2702 2613 2736 2642
rect 2702 2608 2736 2613
rect 2702 2545 2736 2567
rect 2702 2533 2736 2545
rect 2702 2477 2736 2492
rect 2702 2458 2736 2477
rect 2702 2409 2736 2417
rect 2702 2383 2736 2409
rect 2702 2341 2736 2342
rect 2702 2308 2736 2341
rect 2702 2239 2736 2267
rect 2702 2233 2736 2239
rect 2702 2171 2736 2192
rect 2702 2158 2736 2171
rect 2702 2103 2736 2117
rect 2702 2083 2736 2103
rect 2702 2035 2736 2042
rect 2702 2008 2736 2035
rect 2702 1933 2736 1967
rect 2858 2851 2892 2867
rect 2858 2833 2892 2851
rect 2858 2783 2892 2792
rect 2858 2758 2892 2783
rect 2858 2715 2892 2717
rect 2858 2683 2892 2715
rect 2858 2613 2892 2642
rect 2858 2608 2892 2613
rect 2858 2545 2892 2567
rect 2858 2533 2892 2545
rect 2858 2477 2892 2492
rect 2858 2458 2892 2477
rect 2858 2409 2892 2417
rect 2858 2383 2892 2409
rect 2858 2341 2892 2342
rect 2858 2308 2892 2341
rect 2858 2239 2892 2267
rect 2858 2233 2892 2239
rect 2858 2171 2892 2192
rect 2858 2158 2892 2171
rect 2858 2103 2892 2117
rect 2858 2083 2892 2103
rect 2858 2035 2892 2042
rect 2858 2008 2892 2035
rect 2858 1933 2892 1967
rect 3014 2851 3048 2867
rect 3014 2833 3048 2851
rect 3014 2783 3048 2792
rect 3014 2758 3048 2783
rect 3014 2715 3048 2717
rect 3014 2683 3048 2715
rect 3014 2613 3048 2642
rect 3014 2608 3048 2613
rect 3014 2545 3048 2567
rect 3014 2533 3048 2545
rect 3014 2477 3048 2492
rect 3014 2458 3048 2477
rect 3014 2409 3048 2417
rect 3014 2383 3048 2409
rect 3014 2341 3048 2342
rect 3014 2308 3048 2341
rect 3014 2239 3048 2267
rect 3014 2233 3048 2239
rect 3014 2171 3048 2192
rect 3014 2158 3048 2171
rect 3014 2103 3048 2117
rect 3014 2083 3048 2103
rect 3014 2035 3048 2042
rect 3014 2008 3048 2035
rect 3014 1933 3048 1967
rect 3170 2851 3204 2867
rect 3170 2833 3204 2851
rect 3170 2783 3204 2792
rect 3170 2758 3204 2783
rect 3170 2715 3204 2717
rect 3170 2683 3204 2715
rect 3170 2613 3204 2642
rect 3170 2608 3204 2613
rect 3170 2545 3204 2567
rect 3170 2533 3204 2545
rect 3170 2477 3204 2492
rect 3170 2458 3204 2477
rect 3170 2409 3204 2417
rect 3170 2383 3204 2409
rect 3170 2341 3204 2342
rect 3170 2308 3204 2341
rect 3170 2239 3204 2267
rect 3170 2233 3204 2239
rect 3170 2171 3204 2192
rect 3170 2158 3204 2171
rect 3170 2103 3204 2117
rect 3170 2083 3204 2103
rect 3170 2035 3204 2042
rect 3170 2008 3204 2035
rect 3170 1933 3204 1967
rect 3326 2851 3360 2867
rect 3326 2833 3360 2851
rect 3326 2783 3360 2792
rect 3326 2758 3360 2783
rect 3326 2715 3360 2717
rect 3326 2683 3360 2715
rect 3326 2613 3360 2642
rect 3326 2608 3360 2613
rect 3326 2545 3360 2567
rect 3326 2533 3360 2545
rect 3326 2477 3360 2492
rect 3326 2458 3360 2477
rect 3326 2409 3360 2417
rect 3326 2383 3360 2409
rect 3326 2341 3360 2342
rect 3326 2308 3360 2341
rect 3326 2239 3360 2267
rect 3326 2233 3360 2239
rect 3326 2171 3360 2192
rect 3326 2158 3360 2171
rect 3326 2103 3360 2117
rect 3326 2083 3360 2103
rect 3326 2035 3360 2042
rect 3326 2008 3360 2035
rect 3326 1933 3360 1967
rect 3482 2851 3516 2867
rect 3482 2833 3516 2851
rect 3482 2783 3516 2792
rect 3482 2758 3516 2783
rect 3482 2715 3516 2717
rect 3482 2683 3516 2715
rect 3482 2613 3516 2642
rect 3482 2608 3516 2613
rect 3482 2545 3516 2567
rect 3482 2533 3516 2545
rect 3482 2477 3516 2492
rect 3482 2458 3516 2477
rect 3482 2409 3516 2417
rect 3482 2383 3516 2409
rect 3482 2341 3516 2342
rect 3482 2308 3516 2341
rect 3482 2239 3516 2267
rect 3482 2233 3516 2239
rect 3482 2171 3516 2192
rect 3482 2158 3516 2171
rect 3482 2103 3516 2117
rect 3482 2083 3516 2103
rect 3482 2035 3516 2042
rect 3482 2008 3516 2035
rect 3482 1933 3516 1967
rect 3638 2851 3672 2867
rect 3638 2833 3672 2851
rect 3638 2783 3672 2789
rect 3638 2755 3672 2783
rect 3638 2681 3672 2711
rect 3638 2677 3672 2681
rect 3638 2613 3672 2633
rect 3638 2599 3672 2613
rect 3638 2545 3672 2554
rect 3638 2520 3672 2545
rect 3638 2443 3672 2475
rect 3638 2441 3672 2443
rect 3638 2375 3672 2396
rect 3638 2362 3672 2375
rect 3638 2307 3672 2317
rect 3638 2283 3672 2307
rect 3638 2205 3672 2238
rect 3638 2204 3672 2205
rect 3638 2137 3672 2159
rect 3638 2125 3672 2137
rect 3638 2069 3672 2080
rect 3638 2046 3672 2069
rect 3794 2851 3828 2867
rect 3794 2833 3828 2851
rect 3794 2783 3828 2792
rect 3794 2758 3828 2783
rect 3794 2715 3828 2717
rect 3794 2683 3828 2715
rect 3794 2613 3828 2642
rect 3794 2608 3828 2613
rect 3794 2545 3828 2567
rect 3794 2533 3828 2545
rect 3794 2477 3828 2492
rect 3794 2458 3828 2477
rect 3794 2409 3828 2417
rect 3794 2383 3828 2409
rect 3794 2341 3828 2342
rect 3794 2308 3828 2341
rect 3794 2239 3828 2267
rect 3794 2233 3828 2239
rect 3794 2171 3828 2192
rect 3794 2158 3828 2171
rect 3794 2103 3828 2117
rect 3794 2083 3828 2103
rect 3794 2035 3828 2042
rect 3794 2008 3828 2035
rect 3794 1933 3828 1967
rect 3950 2851 3984 2867
rect 3950 2833 3984 2851
rect 3950 2783 3984 2790
rect 3950 2756 3984 2783
rect 3950 2681 3984 2712
rect 3950 2678 3984 2681
rect 3950 2613 3984 2634
rect 3950 2600 3984 2613
rect 3950 2545 3984 2556
rect 3950 2522 3984 2545
rect 3950 2477 3984 2478
rect 3950 2444 3984 2477
rect 3950 2375 3984 2400
rect 3950 2366 3984 2375
rect 3950 2307 3984 2322
rect 3950 2288 3984 2307
rect 3950 2239 3984 2244
rect 3950 2210 3984 2239
rect 3950 2137 3984 2166
rect 3950 2132 3984 2137
rect 3950 2069 3984 2088
rect 3950 2054 3984 2069
rect 4106 2851 4140 2867
rect 4106 2833 4140 2851
rect 4106 2783 4140 2792
rect 4106 2758 4140 2783
rect 4106 2715 4140 2717
rect 4106 2683 4140 2715
rect 4106 2613 4140 2642
rect 4106 2608 4140 2613
rect 4673 2811 4707 2827
rect 4673 2793 4707 2811
rect 4673 2743 4707 2753
rect 4673 2719 4707 2743
rect 4673 2675 4707 2679
rect 4673 2645 4707 2675
rect 4304 2569 4311 2603
rect 4311 2569 4338 2603
rect 4388 2569 4406 2603
rect 4406 2569 4422 2603
rect 4471 2569 4501 2603
rect 4501 2569 4505 2603
rect 4106 2545 4140 2567
rect 4106 2533 4140 2545
rect 4106 2477 4140 2492
rect 4106 2458 4140 2477
rect 4673 2573 4707 2605
rect 4673 2571 4707 2573
rect 4673 2505 4707 2531
rect 4673 2497 4707 2505
rect 4106 2409 4140 2417
rect 4106 2383 4140 2409
rect 4106 2341 4140 2342
rect 4106 2308 4140 2341
rect 4106 2239 4140 2267
rect 4106 2233 4140 2239
rect 4106 2171 4140 2192
rect 4106 2158 4140 2171
rect 4106 2103 4140 2117
rect 4106 2083 4140 2103
rect 4106 2035 4140 2042
rect 4106 2008 4140 2035
rect 4106 1933 4140 1967
rect 4216 2443 4250 2459
rect 4216 2425 4250 2443
rect 4216 2375 4250 2377
rect 4216 2343 4250 2375
rect 4216 2273 4250 2295
rect 4216 2261 4250 2273
rect 4216 2205 4250 2213
rect 4216 2179 4250 2205
rect 4216 2103 4250 2131
rect 4216 2097 4250 2103
rect 4216 2035 4250 2049
rect 4216 2015 4250 2035
rect 4216 1933 4250 1967
rect 4372 2443 4406 2459
rect 4372 2425 4406 2443
rect 4372 2375 4406 2377
rect 4372 2343 4406 2375
rect 4372 2273 4406 2295
rect 4372 2261 4406 2273
rect 4372 2205 4406 2213
rect 4372 2179 4406 2205
rect 4372 2103 4406 2131
rect 4372 2097 4406 2103
rect 4372 2035 4406 2049
rect 4372 2015 4406 2035
rect 4372 1933 4406 1967
rect 4528 2443 4562 2459
rect 4528 2425 4562 2443
rect 4528 2375 4562 2377
rect 4528 2343 4562 2375
rect 4528 2273 4562 2295
rect 4528 2261 4562 2273
rect 4528 2205 4562 2213
rect 4528 2179 4562 2205
rect 4528 2103 4562 2131
rect 4528 2097 4562 2103
rect 4528 2035 4562 2049
rect 4528 2015 4562 2035
rect 4528 1933 4562 1967
rect 4673 2437 4707 2457
rect 4673 2423 4707 2437
rect 4673 2369 4707 2383
rect 4673 2349 4707 2369
rect 4673 2301 4707 2309
rect 4673 2275 4707 2301
rect 4673 2233 4707 2235
rect 4673 2201 4707 2233
rect 4673 2131 4707 2161
rect 4673 2127 4707 2131
rect 4673 2063 4707 2086
rect 4673 2052 4707 2063
rect 4673 1995 4707 2011
rect 4673 1977 4707 1995
rect 4673 1927 4707 1936
rect 4673 1902 4707 1927
rect 433 1850 467 1862
rect 433 1828 467 1850
rect 717 1839 751 1873
rect 817 1839 851 1873
rect 917 1839 951 1873
rect 1245 1839 1277 1873
rect 1277 1839 1279 1873
rect 1318 1839 1351 1873
rect 1351 1839 1352 1873
rect 1391 1839 1425 1873
rect 1464 1839 1498 1873
rect 1537 1839 1571 1873
rect 1610 1839 1644 1873
rect 1682 1839 1716 1873
rect 1754 1839 1755 1873
rect 1755 1839 1788 1873
rect 1826 1839 1829 1873
rect 1829 1839 1860 1873
rect 1898 1839 1903 1873
rect 1903 1839 1932 1873
rect 1970 1839 1977 1873
rect 1977 1839 2004 1873
rect 2166 1839 2173 1873
rect 2173 1839 2200 1873
rect 2239 1839 2244 1873
rect 2244 1839 2273 1873
rect 2312 1839 2315 1873
rect 2315 1839 2346 1873
rect 2385 1839 2387 1873
rect 2387 1839 2419 1873
rect 2457 1839 2459 1873
rect 2459 1839 2491 1873
rect 2529 1839 2531 1873
rect 2531 1839 2563 1873
rect 2762 1839 2763 1873
rect 2763 1839 2796 1873
rect 2845 1839 2869 1873
rect 2869 1839 2879 1873
rect 2928 1839 2941 1873
rect 2941 1839 2962 1873
rect 3011 1839 3013 1873
rect 3013 1839 3045 1873
rect 3094 1839 3123 1873
rect 3123 1839 3128 1873
rect 3176 1839 3194 1873
rect 3194 1839 3210 1873
rect 3258 1839 3265 1873
rect 3265 1839 3292 1873
rect 3661 1839 3680 1873
rect 3680 1839 3695 1873
rect 3734 1839 3753 1873
rect 3753 1839 3768 1873
rect 3807 1839 3826 1873
rect 3826 1839 3841 1873
rect 3880 1839 3899 1873
rect 3899 1839 3914 1873
rect 3953 1839 3972 1873
rect 3972 1839 3987 1873
rect 4025 1839 4045 1873
rect 4045 1839 4059 1873
rect 433 1782 467 1788
rect 433 1754 467 1782
rect 4673 1859 4707 1861
rect 4673 1827 4707 1859
rect 4673 1754 4707 1786
rect 4673 1752 4707 1754
rect 1067 1680 1069 1714
rect 1069 1680 1101 1714
rect 1144 1680 1171 1714
rect 1171 1680 1178 1714
rect 1221 1680 1239 1714
rect 1239 1680 1255 1714
rect 1298 1680 1307 1714
rect 1307 1680 1332 1714
rect 1375 1680 1409 1714
rect 1451 1680 1477 1714
rect 1477 1680 1485 1714
rect 1527 1680 1545 1714
rect 1545 1680 1561 1714
rect 1603 1680 1613 1714
rect 1613 1680 1637 1714
rect 1679 1680 1681 1714
rect 1681 1680 1713 1714
rect 1755 1680 1783 1714
rect 1783 1680 1789 1714
rect 1831 1680 1851 1714
rect 1851 1680 1865 1714
rect 1907 1680 1919 1714
rect 1919 1680 1941 1714
rect 1983 1680 1987 1714
rect 1987 1680 2017 1714
rect 2059 1680 2089 1714
rect 2089 1680 2093 1714
rect 2135 1680 2157 1714
rect 2157 1680 2169 1714
rect 2396 1680 2429 1714
rect 2429 1680 2430 1714
rect 2476 1680 2497 1714
rect 2497 1680 2510 1714
rect 2556 1680 2565 1714
rect 2565 1680 2590 1714
rect 2636 1680 2667 1714
rect 2667 1680 2670 1714
rect 2716 1680 2735 1714
rect 2735 1680 2750 1714
rect 2795 1680 2803 1714
rect 2803 1680 2829 1714
rect 2874 1680 2905 1714
rect 2905 1680 2908 1714
rect 2984 1680 3007 1714
rect 3007 1680 3018 1714
rect 3059 1680 3075 1714
rect 3075 1680 3093 1714
rect 3134 1680 3143 1714
rect 3143 1680 3168 1714
rect 3209 1680 3211 1714
rect 3211 1680 3243 1714
rect 3284 1680 3313 1714
rect 3313 1680 3318 1714
rect 3359 1680 3381 1714
rect 3381 1680 3393 1714
rect 3434 1680 3449 1714
rect 3449 1680 3468 1714
rect 4173 1680 4197 1714
rect 4197 1680 4207 1714
rect 4257 1680 4265 1714
rect 4265 1680 4291 1714
rect 4341 1680 4367 1714
rect 4367 1680 4375 1714
rect 4424 1680 4435 1714
rect 4435 1680 4458 1714
rect 4507 1680 4537 1714
rect 4537 1680 4541 1714
rect 4590 1680 4605 1714
rect 4605 1680 4624 1714
rect 4896 3034 4930 3050
rect 4896 3016 4930 3034
rect 4896 2966 4930 2976
rect 4896 2942 4930 2966
rect 4896 2898 4930 2902
rect 4896 2868 4930 2898
rect 4896 2796 4930 2828
rect 4896 2794 4930 2796
rect 4896 2728 4930 2754
rect 4896 2720 4930 2728
rect 4896 2660 4930 2680
rect 4896 2646 4930 2660
rect 4896 2592 4930 2606
rect 4896 2572 4930 2592
rect 4896 2524 4930 2532
rect 4896 2498 4930 2524
rect 4896 2456 4930 2458
rect 4896 2424 4930 2456
rect 4896 2354 4930 2384
rect 4896 2350 4930 2354
rect 4896 2286 4930 2310
rect 4896 2276 4930 2286
rect 4896 2218 4930 2236
rect 4896 2202 4930 2218
rect 4896 2150 4930 2161
rect 4896 2127 4930 2150
rect 4896 2082 4930 2086
rect 4896 2052 4930 2082
rect 4896 1980 4930 2011
rect 4896 1977 4930 1980
rect 4896 1912 4930 1936
rect 4896 1902 4930 1912
rect 4896 1844 4930 1861
rect 4896 1827 4930 1844
rect 4896 1776 4930 1786
rect 4896 1752 4930 1776
rect 4896 1708 4930 1711
rect 4896 1677 4930 1708
rect 4896 1606 4930 1636
rect 4896 1602 4930 1606
rect 4896 1527 4930 1561
rect 957 1457 986 1490
rect 986 1457 991 1490
rect 1031 1457 1054 1490
rect 1054 1457 1065 1490
rect 1105 1457 1122 1490
rect 1122 1457 1139 1490
rect 1179 1457 1190 1490
rect 1190 1457 1213 1490
rect 1253 1457 1258 1490
rect 1258 1457 1287 1490
rect 1327 1457 1360 1490
rect 1360 1457 1361 1490
rect 1401 1457 1428 1490
rect 1428 1457 1435 1490
rect 1475 1457 1496 1490
rect 1496 1457 1509 1490
rect 1549 1457 1564 1490
rect 1564 1457 1583 1490
rect 1623 1457 1632 1490
rect 1632 1457 1657 1490
rect 1697 1457 1700 1490
rect 1700 1457 1731 1490
rect 1771 1457 1802 1490
rect 1802 1457 1805 1490
rect 1845 1457 1870 1490
rect 1870 1457 1879 1490
rect 1919 1457 1938 1490
rect 1938 1457 1953 1490
rect 1993 1457 2006 1490
rect 2006 1457 2027 1490
rect 2068 1457 2074 1490
rect 2074 1457 2102 1490
rect 2143 1457 2176 1490
rect 2176 1457 2177 1490
rect 2375 1457 2380 1490
rect 2380 1457 2409 1490
rect 2449 1457 2482 1490
rect 2482 1457 2483 1490
rect 2523 1457 2550 1490
rect 2550 1457 2557 1490
rect 2597 1457 2618 1490
rect 2618 1457 2631 1490
rect 2671 1457 2686 1490
rect 2686 1457 2705 1490
rect 2745 1457 2754 1490
rect 2754 1457 2779 1490
rect 2819 1457 2822 1490
rect 2822 1457 2853 1490
rect 2893 1457 2924 1490
rect 2924 1457 2927 1490
rect 2967 1457 2992 1490
rect 2992 1457 3001 1490
rect 3041 1457 3060 1490
rect 3060 1457 3075 1490
rect 3115 1457 3128 1490
rect 3128 1457 3149 1490
rect 3190 1457 3196 1490
rect 3196 1457 3224 1490
rect 3265 1457 3298 1490
rect 3298 1457 3299 1490
rect 3340 1457 3366 1490
rect 3366 1457 3374 1490
rect 3415 1457 3434 1490
rect 3434 1457 3449 1490
rect 3490 1457 3502 1490
rect 3502 1457 3524 1490
rect 3565 1457 3570 1490
rect 3570 1457 3599 1490
rect 3640 1457 3672 1490
rect 3672 1457 3674 1490
rect 3715 1457 3740 1490
rect 3740 1457 3749 1490
rect 3790 1457 3808 1490
rect 3808 1457 3824 1490
rect 3865 1457 3876 1490
rect 3876 1457 3899 1490
rect 4112 1457 4114 1489
rect 4114 1457 4146 1489
rect 4191 1457 4216 1489
rect 4216 1457 4225 1489
rect 4270 1457 4284 1489
rect 4284 1457 4304 1489
rect 4349 1457 4352 1489
rect 4352 1457 4383 1489
rect 4428 1457 4454 1489
rect 4454 1457 4462 1489
rect 4506 1457 4522 1489
rect 4522 1457 4540 1489
rect 4584 1457 4590 1489
rect 4590 1457 4618 1489
rect 4662 1457 4692 1489
rect 4692 1457 4696 1489
rect 4740 1457 4760 1489
rect 4760 1457 4774 1489
rect 4818 1457 4828 1489
rect 4828 1457 4852 1489
rect 957 1456 991 1457
rect 1031 1456 1065 1457
rect 1105 1456 1139 1457
rect 1179 1456 1213 1457
rect 1253 1456 1287 1457
rect 1327 1456 1361 1457
rect 1401 1456 1435 1457
rect 1475 1456 1509 1457
rect 1549 1456 1583 1457
rect 1623 1456 1657 1457
rect 1697 1456 1731 1457
rect 1771 1456 1805 1457
rect 1845 1456 1879 1457
rect 1919 1456 1953 1457
rect 1993 1456 2027 1457
rect 2068 1456 2102 1457
rect 2143 1456 2177 1457
rect 2375 1456 2409 1457
rect 2449 1456 2483 1457
rect 2523 1456 2557 1457
rect 2597 1456 2631 1457
rect 2671 1456 2705 1457
rect 2745 1456 2779 1457
rect 2819 1456 2853 1457
rect 2893 1456 2927 1457
rect 2967 1456 3001 1457
rect 3041 1456 3075 1457
rect 3115 1456 3149 1457
rect 3190 1456 3224 1457
rect 3265 1456 3299 1457
rect 3340 1456 3374 1457
rect 3415 1456 3449 1457
rect 3490 1456 3524 1457
rect 3565 1456 3599 1457
rect 3640 1456 3674 1457
rect 3715 1456 3749 1457
rect 3790 1456 3824 1457
rect 3865 1456 3899 1457
rect 4112 1455 4146 1457
rect 4191 1455 4225 1457
rect 4270 1455 4304 1457
rect 4349 1455 4383 1457
rect 4428 1455 4462 1457
rect 4506 1455 4540 1457
rect 4584 1455 4618 1457
rect 4662 1455 4696 1457
rect 4740 1455 4774 1457
rect 4818 1455 4852 1457
rect 5170 3238 5177 3272
rect 5177 3238 5204 3272
rect 5245 3238 5279 3272
rect 5320 3238 5347 3272
rect 5347 3238 5354 3272
rect 5395 3238 5415 3272
rect 5415 3238 5429 3272
rect 5470 3238 5483 3272
rect 5483 3238 5504 3272
rect 5545 3238 5551 3272
rect 5551 3238 5579 3272
rect 5619 3238 5653 3272
rect 5693 3238 5721 3272
rect 5721 3238 5727 3272
rect 5767 3238 5789 3272
rect 5789 3238 5801 3272
rect 5841 3238 5857 3272
rect 5857 3238 5875 3272
rect 5915 3238 5925 3272
rect 5925 3238 5949 3272
rect 5989 3238 5993 3272
rect 5993 3238 6023 3272
rect 6063 3238 6095 3272
rect 6095 3238 6097 3272
rect 6137 3238 6163 3272
rect 6163 3238 6171 3272
rect 6211 3238 6231 3272
rect 6231 3238 6245 3272
rect 6285 3238 6299 3272
rect 6299 3238 6319 3272
rect 6359 3238 6367 3272
rect 6367 3238 6393 3272
rect 6433 3238 6435 3272
rect 6435 3238 6467 3272
rect 6507 3238 6537 3272
rect 6537 3238 6541 3272
rect 6581 3238 6605 3272
rect 6605 3238 6615 3272
rect 6655 3238 6673 3272
rect 6673 3238 6689 3272
rect 6729 3238 6741 3272
rect 6741 3238 6763 3272
rect 6803 3238 6809 3272
rect 6809 3238 6837 3272
rect 5098 3170 5099 3198
rect 5099 3170 5132 3198
rect 5098 3164 5132 3170
rect 5098 3102 5099 3124
rect 5099 3102 5132 3124
rect 5098 3090 5132 3102
rect 6877 3191 6911 3200
rect 6877 3166 6911 3191
rect 6877 3123 6911 3126
rect 6877 3092 6911 3123
rect 5098 3034 5099 3050
rect 5099 3034 5132 3050
rect 5098 3016 5132 3034
rect 5098 2966 5099 2976
rect 5099 2966 5132 2976
rect 5098 2942 5132 2966
rect 5098 2898 5099 2902
rect 5099 2898 5132 2902
rect 5098 2868 5132 2898
rect 5098 2796 5132 2828
rect 5098 2794 5099 2796
rect 5099 2794 5132 2796
rect 5098 2728 5132 2754
rect 5098 2720 5099 2728
rect 5099 2720 5132 2728
rect 5098 2660 5132 2680
rect 5098 2646 5099 2660
rect 5099 2646 5132 2660
rect 5098 2592 5132 2606
rect 5098 2572 5099 2592
rect 5099 2572 5132 2592
rect 5098 2524 5132 2532
rect 5098 2498 5099 2524
rect 5099 2498 5132 2524
rect 5098 2456 5132 2458
rect 5098 2424 5099 2456
rect 5099 2424 5132 2456
rect 5098 2354 5099 2384
rect 5099 2354 5132 2384
rect 5098 2350 5132 2354
rect 5098 2286 5099 2310
rect 5099 2286 5132 2310
rect 5098 2276 5132 2286
rect 5098 2218 5099 2236
rect 5099 2218 5132 2236
rect 5098 2202 5132 2218
rect 5098 2150 5099 2162
rect 5099 2150 5132 2162
rect 5098 2128 5132 2150
rect 5098 2082 5099 2088
rect 5099 2082 5132 2088
rect 5098 2054 5132 2082
rect 5098 1980 5132 2013
rect 5098 1979 5099 1980
rect 5099 1979 5132 1980
rect 5098 1912 5132 1938
rect 5098 1904 5099 1912
rect 5099 1904 5132 1912
rect 5098 1844 5132 1863
rect 5098 1829 5099 1844
rect 5099 1829 5132 1844
rect 5098 1776 5132 1788
rect 5098 1754 5099 1776
rect 5099 1754 5132 1776
rect 5098 1708 5132 1713
rect 5098 1679 5099 1708
rect 5099 1679 5132 1708
rect 5443 3015 5467 3049
rect 5467 3015 5477 3049
rect 5530 3015 5535 3049
rect 5535 3015 5564 3049
rect 5640 3015 5671 3049
rect 5671 3015 5674 3049
rect 5712 3015 5739 3049
rect 5739 3015 5746 3049
rect 5784 3015 5807 3049
rect 5807 3015 5818 3049
rect 5856 3015 5875 3049
rect 5875 3015 5890 3049
rect 5928 3015 5943 3049
rect 5943 3015 5962 3049
rect 6001 3015 6011 3049
rect 6011 3015 6035 3049
rect 6074 3015 6079 3049
rect 6079 3015 6108 3049
rect 6147 3015 6181 3049
rect 6220 3015 6249 3049
rect 6249 3015 6254 3049
rect 6293 3015 6317 3049
rect 6317 3015 6327 3049
rect 6366 3015 6385 3049
rect 6385 3015 6400 3049
rect 6439 3015 6453 3049
rect 6453 3015 6473 3049
rect 6512 3015 6521 3049
rect 6521 3015 6546 3049
rect 6585 3015 6589 3049
rect 6589 3015 6619 3049
rect 5357 2947 5391 2977
rect 5357 2943 5391 2947
rect 5357 2879 5391 2902
rect 5357 2868 5391 2879
rect 6657 2941 6691 2975
rect 5357 2811 5391 2827
rect 5357 2793 5391 2811
rect 5357 2743 5391 2752
rect 5357 2718 5391 2743
rect 5357 2675 5391 2677
rect 5357 2643 5391 2675
rect 5357 2573 5391 2602
rect 5357 2568 5391 2573
rect 5357 2505 5391 2528
rect 5357 2494 5391 2505
rect 5357 2437 5391 2454
rect 5357 2420 5391 2437
rect 5357 2369 5391 2380
rect 5357 2346 5391 2369
rect 5357 2301 5391 2306
rect 5357 2272 5391 2301
rect 5357 2199 5391 2232
rect 5357 2198 5391 2199
rect 5357 2131 5391 2158
rect 5357 2124 5391 2131
rect 5357 2063 5391 2084
rect 5357 2050 5391 2063
rect 5357 1995 5391 2010
rect 5357 1976 5391 1995
rect 5357 1927 5391 1936
rect 5357 1902 5391 1927
rect 5502 2851 5536 2867
rect 5502 2833 5536 2851
rect 5502 2783 5536 2792
rect 5502 2758 5536 2783
rect 5502 2715 5536 2717
rect 5502 2683 5536 2715
rect 5502 2613 5536 2642
rect 5502 2608 5536 2613
rect 5502 2545 5536 2567
rect 5502 2533 5536 2545
rect 5502 2477 5536 2492
rect 5502 2458 5536 2477
rect 5502 2409 5536 2417
rect 5502 2383 5536 2409
rect 5502 2341 5536 2342
rect 5502 2308 5536 2341
rect 5502 2239 5536 2267
rect 5502 2233 5536 2239
rect 5502 2171 5536 2192
rect 5502 2158 5536 2171
rect 5502 2103 5536 2117
rect 5502 2083 5536 2103
rect 5502 2035 5536 2042
rect 5502 2008 5536 2035
rect 5502 1933 5536 1967
rect 5658 2851 5692 2867
rect 5658 2833 5692 2851
rect 5658 2783 5692 2788
rect 5658 2754 5692 2783
rect 5658 2681 5692 2709
rect 5658 2675 5692 2681
rect 5658 2613 5692 2630
rect 5658 2596 5692 2613
rect 5658 2545 5692 2551
rect 5658 2517 5692 2545
rect 5658 2443 5692 2472
rect 5658 2438 5692 2443
rect 5658 2375 5692 2393
rect 5658 2359 5692 2375
rect 5658 2307 5692 2314
rect 5658 2280 5692 2307
rect 5658 2205 5692 2234
rect 5658 2200 5692 2205
rect 5658 2137 5692 2154
rect 5658 2120 5692 2137
rect 5812 2851 5846 2867
rect 5812 2833 5814 2851
rect 5814 2833 5846 2851
rect 5812 2783 5846 2792
rect 5812 2758 5814 2783
rect 5814 2758 5846 2783
rect 5812 2715 5846 2717
rect 5812 2683 5814 2715
rect 5814 2683 5846 2715
rect 5812 2613 5814 2642
rect 5814 2613 5846 2642
rect 5812 2608 5846 2613
rect 5812 2545 5814 2567
rect 5814 2545 5846 2567
rect 5812 2533 5846 2545
rect 5812 2477 5814 2492
rect 5814 2477 5846 2492
rect 5812 2458 5846 2477
rect 5812 2409 5814 2417
rect 5814 2409 5846 2417
rect 5812 2383 5846 2409
rect 5812 2341 5814 2342
rect 5814 2341 5846 2342
rect 5812 2308 5846 2341
rect 5812 2239 5846 2267
rect 5812 2233 5814 2239
rect 5814 2233 5846 2239
rect 5812 2171 5846 2192
rect 5812 2158 5814 2171
rect 5814 2158 5846 2171
rect 5812 2103 5846 2117
rect 5812 2083 5814 2103
rect 5814 2083 5846 2103
rect 5812 2035 5846 2042
rect 5812 2008 5814 2035
rect 5814 2008 5846 2035
rect 5812 1933 5814 1967
rect 5814 1933 5846 1967
rect 6030 2851 6064 2867
rect 6030 2833 6064 2851
rect 6030 2783 6064 2792
rect 6030 2758 6064 2783
rect 6030 2715 6064 2717
rect 6030 2683 6064 2715
rect 6030 2613 6064 2642
rect 6030 2608 6064 2613
rect 6030 2545 6064 2567
rect 6030 2533 6064 2545
rect 6030 2477 6064 2492
rect 6030 2458 6064 2477
rect 6030 2409 6064 2417
rect 6030 2383 6064 2409
rect 6030 2341 6064 2342
rect 6030 2308 6064 2341
rect 6030 2239 6064 2267
rect 6030 2233 6064 2239
rect 6030 2171 6064 2192
rect 6030 2158 6064 2171
rect 6030 2103 6064 2117
rect 6030 2083 6064 2103
rect 6030 2035 6064 2042
rect 6030 2008 6064 2035
rect 6030 1933 6064 1967
rect 6246 2851 6280 2867
rect 6246 2833 6280 2851
rect 6246 2783 6280 2792
rect 6246 2758 6280 2783
rect 6246 2715 6280 2717
rect 6246 2683 6280 2715
rect 6246 2613 6280 2642
rect 6246 2608 6280 2613
rect 6246 2545 6280 2567
rect 6246 2533 6280 2545
rect 6512 2833 6546 2867
rect 6512 2754 6546 2788
rect 6512 2675 6546 2709
rect 6512 2595 6546 2629
rect 6246 2477 6280 2492
rect 6246 2458 6280 2477
rect 6246 2409 6280 2417
rect 6246 2383 6280 2409
rect 6246 2341 6280 2342
rect 6246 2308 6280 2341
rect 6356 2503 6390 2509
rect 6356 2475 6390 2503
rect 6356 2367 6390 2389
rect 6356 2355 6390 2367
rect 6512 2515 6546 2549
rect 6512 2435 6546 2469
rect 6512 2367 6546 2389
rect 6512 2355 6546 2367
rect 6657 2870 6691 2901
rect 6657 2867 6691 2870
rect 6657 2802 6691 2827
rect 6657 2793 6691 2802
rect 6657 2734 6691 2753
rect 6657 2719 6691 2734
rect 6657 2666 6691 2679
rect 6657 2645 6691 2666
rect 6657 2598 6691 2605
rect 6657 2571 6691 2598
rect 6657 2530 6691 2531
rect 6657 2497 6691 2530
rect 6657 2428 6691 2457
rect 6657 2423 6691 2428
rect 6657 2360 6691 2383
rect 6657 2349 6691 2360
rect 6657 2292 6691 2309
rect 6657 2275 6691 2292
rect 6246 2239 6280 2267
rect 6436 2239 6451 2273
rect 6451 2239 6470 2273
rect 6508 2239 6519 2273
rect 6519 2239 6542 2273
rect 6246 2233 6280 2239
rect 6246 2171 6280 2192
rect 6246 2158 6280 2171
rect 6246 2103 6280 2117
rect 6246 2083 6280 2103
rect 6246 2035 6280 2042
rect 6246 2008 6280 2035
rect 6246 1933 6280 1967
rect 6657 2224 6691 2235
rect 6657 2201 6691 2224
rect 6657 2156 6691 2161
rect 6657 2127 6691 2156
rect 6657 2054 6691 2086
rect 6657 2052 6691 2054
rect 6657 1986 6691 2011
rect 6657 1977 6691 1986
rect 5357 1859 5391 1862
rect 5357 1828 5391 1859
rect 6657 1918 6691 1936
rect 6657 1902 6691 1918
rect 5563 1839 5597 1873
rect 5648 1839 5658 1873
rect 5658 1839 5682 1873
rect 5733 1839 5753 1873
rect 5753 1839 5767 1873
rect 5879 1839 5909 1873
rect 5909 1839 5913 1873
rect 5956 1839 5987 1873
rect 5987 1839 5990 1873
rect 6033 1839 6065 1873
rect 6065 1839 6067 1873
rect 6110 1839 6142 1873
rect 6142 1839 6144 1873
rect 6186 1839 6219 1873
rect 6219 1839 6220 1873
rect 5357 1754 5391 1788
rect 6657 1850 6691 1861
rect 6657 1827 6691 1850
rect 6657 1782 6691 1786
rect 6657 1752 6691 1782
rect 5429 1680 5459 1714
rect 5459 1680 5463 1714
rect 5511 1680 5527 1714
rect 5527 1680 5545 1714
rect 5592 1680 5595 1714
rect 5595 1680 5626 1714
rect 5673 1680 5697 1714
rect 5697 1680 5707 1714
rect 5754 1680 5765 1714
rect 5765 1680 5788 1714
rect 6566 1680 6581 1714
rect 6581 1680 6600 1714
rect 6877 3021 6911 3052
rect 6877 3018 6911 3021
rect 6877 2953 6911 2978
rect 6877 2944 6911 2953
rect 6877 2885 6911 2904
rect 6877 2870 6911 2885
rect 6877 2817 6911 2830
rect 6877 2796 6911 2817
rect 6877 2749 6911 2757
rect 6877 2723 6911 2749
rect 6877 2681 6911 2684
rect 6877 2650 6911 2681
rect 6877 2579 6911 2611
rect 6877 2577 6911 2579
rect 6877 2511 6911 2538
rect 6877 2504 6911 2511
rect 6877 2443 6911 2465
rect 6877 2431 6911 2443
rect 6877 2375 6911 2392
rect 6877 2358 6911 2375
rect 6877 2307 6911 2319
rect 6877 2285 6911 2307
rect 6877 2239 6911 2246
rect 6877 2212 6911 2239
rect 6877 2171 6911 2173
rect 6877 2139 6911 2171
rect 6877 2069 6911 2100
rect 6877 2066 6911 2069
rect 6877 2001 6911 2027
rect 6877 1993 6911 2001
rect 6877 1933 6911 1954
rect 6877 1920 6911 1933
rect 6877 1865 6911 1881
rect 6877 1847 6911 1865
rect 6877 1797 6911 1808
rect 6877 1774 6911 1797
rect 6877 1729 6911 1735
rect 6877 1701 6911 1729
rect 5098 1606 5099 1638
rect 5099 1606 5132 1638
rect 5098 1604 5132 1606
rect 5098 1529 5132 1563
rect 6877 1661 6911 1662
rect 6877 1628 6911 1661
rect 6877 1559 6911 1589
rect 6877 1555 6911 1559
rect 6241 1491 6275 1492
rect 6319 1491 6353 1492
rect 6397 1491 6431 1492
rect 6476 1491 6510 1492
rect 6555 1491 6589 1492
rect 6634 1491 6668 1492
rect 6713 1491 6747 1492
rect 6792 1491 6826 1492
rect 5170 1457 5201 1491
rect 5201 1457 5204 1491
rect 5242 1457 5269 1491
rect 5269 1457 5276 1491
rect 5314 1457 5337 1491
rect 5337 1457 5348 1491
rect 5386 1457 5405 1491
rect 5405 1457 5420 1491
rect 5458 1457 5473 1491
rect 5473 1457 5492 1491
rect 5530 1457 5541 1491
rect 5541 1457 5564 1491
rect 5602 1457 5609 1491
rect 5609 1457 5636 1491
rect 5675 1457 5677 1491
rect 5677 1457 5709 1491
rect 5748 1457 5779 1491
rect 5779 1457 5782 1491
rect 6241 1458 6255 1491
rect 6255 1458 6275 1491
rect 6319 1458 6323 1491
rect 6323 1458 6353 1491
rect 6397 1458 6425 1491
rect 6425 1458 6431 1491
rect 6476 1458 6493 1491
rect 6493 1458 6510 1491
rect 6555 1458 6561 1491
rect 6561 1458 6589 1491
rect 6634 1458 6663 1491
rect 6663 1458 6668 1491
rect 6713 1458 6731 1491
rect 6731 1458 6747 1491
rect 6792 1458 6799 1491
rect 6799 1458 6826 1491
rect 6871 1458 6905 1492
rect 7077 3238 7111 3272
rect 7155 3238 7182 3272
rect 7182 3238 7189 3272
rect 7233 3238 7250 3272
rect 7250 3238 7267 3272
rect 7311 3238 7318 3272
rect 7318 3238 7345 3272
rect 7390 3238 7420 3272
rect 7420 3238 7424 3272
rect 7469 3238 7488 3272
rect 7488 3238 7503 3272
rect 7548 3238 7556 3272
rect 7556 3238 7582 3272
rect 7627 3238 7658 3272
rect 7658 3238 7661 3272
rect 7737 3238 7760 3272
rect 7760 3238 7771 3272
rect 7812 3238 7828 3272
rect 7828 3238 7846 3272
rect 7887 3238 7896 3272
rect 7896 3238 7921 3272
rect 7962 3238 7964 3272
rect 7964 3238 7996 3272
rect 8037 3238 8066 3272
rect 8066 3238 8071 3272
rect 8112 3238 8134 3272
rect 8134 3238 8146 3272
rect 8187 3238 8202 3272
rect 8202 3238 8221 3272
rect 8262 3238 8270 3272
rect 8270 3238 8296 3272
rect 8338 3238 8372 3272
rect 8414 3238 8440 3272
rect 8440 3238 8448 3272
rect 8490 3238 8508 3272
rect 8508 3238 8524 3272
rect 8566 3238 8576 3272
rect 8576 3238 8600 3272
rect 8642 3238 8644 3272
rect 8644 3238 8676 3272
rect 8718 3238 8746 3272
rect 8746 3238 8752 3272
rect 8794 3238 8814 3272
rect 8814 3238 8828 3272
rect 8870 3238 8882 3272
rect 8882 3238 8904 3272
rect 8946 3238 8950 3272
rect 8950 3238 8980 3272
rect 6999 3170 7033 3200
rect 6999 3166 7033 3170
rect 6999 3102 7033 3127
rect 6999 3093 7033 3102
rect 6999 3034 7033 3054
rect 6999 3020 7033 3034
rect 9018 3191 9052 3198
rect 9018 3164 9052 3191
rect 9018 3123 9052 3124
rect 9018 3090 9052 3123
rect 6999 2966 7033 2981
rect 6999 2947 7033 2966
rect 6999 2898 7033 2908
rect 6999 2874 7033 2898
rect 6999 2830 7033 2835
rect 6999 2801 7033 2830
rect 6999 2728 7033 2762
rect 6999 2660 7033 2689
rect 6999 2655 7033 2660
rect 6999 2592 7033 2616
rect 6999 2582 7033 2592
rect 6999 2524 7033 2543
rect 6999 2509 7033 2524
rect 6999 2456 7033 2470
rect 6999 2436 7033 2456
rect 6999 2388 7033 2397
rect 6999 2363 7033 2388
rect 6999 2320 7033 2324
rect 6999 2290 7033 2320
rect 6999 2218 7033 2251
rect 6999 2217 7033 2218
rect 6999 2150 7033 2178
rect 6999 2144 7033 2150
rect 6999 2082 7033 2105
rect 6999 2071 7033 2082
rect 6999 2014 7033 2032
rect 6999 1998 7033 2014
rect 6999 1946 7033 1960
rect 6999 1926 7033 1946
rect 6999 1878 7033 1888
rect 6999 1854 7033 1878
rect 6999 1810 7033 1816
rect 6999 1782 7033 1810
rect 6999 1742 7033 1744
rect 6999 1710 7033 1742
rect 7302 3015 7333 3049
rect 7333 3015 7336 3049
rect 7380 3015 7401 3049
rect 7401 3015 7414 3049
rect 7458 3015 7469 3049
rect 7469 3015 7492 3049
rect 7536 3015 7537 3049
rect 7537 3015 7570 3049
rect 7646 3015 7673 3049
rect 7673 3015 7680 3049
rect 7722 3015 7741 3049
rect 7741 3015 7756 3049
rect 7799 3015 7809 3049
rect 7809 3015 7833 3049
rect 7876 3015 7877 3049
rect 7877 3015 7910 3049
rect 7953 3015 7979 3049
rect 7979 3015 7987 3049
rect 8030 3015 8047 3049
rect 8047 3015 8064 3049
rect 8107 3015 8115 3049
rect 8115 3015 8141 3049
rect 8184 3015 8217 3049
rect 8217 3015 8218 3049
rect 8261 3015 8285 3049
rect 8285 3015 8295 3049
rect 8338 3015 8353 3049
rect 8353 3015 8372 3049
rect 8415 3015 8421 3049
rect 8421 3015 8449 3049
rect 8492 3015 8523 3049
rect 8523 3015 8526 3049
rect 8569 3015 8591 3049
rect 8591 3015 8603 3049
rect 8646 3015 8659 3049
rect 8659 3015 8680 3049
rect 8723 3015 8727 3049
rect 8727 3015 8757 3049
rect 7225 2947 7259 2977
rect 7225 2943 7259 2947
rect 7225 2879 7259 2903
rect 7225 2869 7259 2879
rect 8795 2941 8829 2975
rect 8018 2878 8052 2912
rect 7225 2811 7259 2829
rect 7225 2795 7259 2811
rect 7225 2743 7259 2755
rect 7225 2721 7259 2743
rect 7225 2675 7259 2682
rect 7225 2648 7259 2675
rect 7225 2607 7259 2609
rect 7225 2575 7259 2607
rect 7225 2505 7259 2536
rect 7225 2502 7259 2505
rect 7225 2437 7259 2463
rect 7225 2429 7259 2437
rect 7225 2369 7259 2390
rect 7225 2356 7259 2369
rect 7225 2301 7259 2317
rect 7225 2283 7259 2301
rect 7225 2233 7259 2244
rect 7225 2210 7259 2233
rect 7225 2165 7259 2171
rect 7225 2137 7259 2165
rect 7225 2097 7259 2098
rect 7225 2064 7259 2097
rect 7225 1995 7259 2025
rect 7225 1991 7259 1995
rect 7225 1927 7259 1952
rect 7225 1918 7259 1927
rect 7370 2851 7404 2867
rect 7370 2833 7404 2851
rect 7370 2783 7404 2792
rect 7370 2758 7404 2783
rect 7370 2715 7404 2717
rect 7370 2683 7404 2715
rect 7370 2613 7404 2642
rect 7370 2608 7404 2613
rect 7370 2545 7404 2567
rect 7370 2533 7404 2545
rect 7370 2477 7404 2492
rect 7370 2458 7404 2477
rect 7370 2409 7404 2417
rect 7370 2383 7404 2409
rect 7370 2341 7404 2342
rect 7370 2308 7404 2341
rect 7370 2239 7404 2267
rect 7370 2233 7404 2239
rect 7370 2171 7404 2192
rect 7370 2158 7404 2171
rect 7370 2103 7404 2117
rect 7370 2083 7404 2103
rect 7370 2035 7404 2042
rect 7370 2008 7404 2035
rect 7370 1933 7404 1967
rect 7586 2851 7620 2867
rect 7586 2833 7620 2851
rect 7586 2783 7620 2792
rect 7586 2758 7620 2783
rect 7586 2715 7620 2717
rect 7586 2683 7620 2715
rect 7586 2613 7620 2642
rect 7586 2608 7620 2613
rect 7586 2545 7620 2567
rect 7586 2533 7620 2545
rect 7586 2477 7620 2492
rect 7586 2458 7620 2477
rect 7586 2409 7620 2417
rect 7586 2383 7620 2409
rect 7586 2341 7620 2342
rect 7586 2308 7620 2341
rect 7586 2239 7620 2267
rect 7586 2233 7620 2239
rect 7586 2171 7620 2192
rect 7586 2158 7620 2171
rect 7586 2103 7620 2117
rect 7586 2083 7620 2103
rect 7586 2035 7620 2042
rect 7586 2008 7620 2035
rect 7586 1933 7620 1967
rect 7802 2851 7836 2867
rect 7802 2833 7836 2851
rect 7802 2783 7836 2792
rect 7802 2758 7836 2783
rect 7802 2715 7836 2717
rect 7802 2683 7836 2715
rect 7802 2613 7836 2642
rect 7802 2608 7836 2613
rect 7802 2545 7836 2567
rect 7802 2533 7836 2545
rect 7802 2477 7836 2492
rect 7802 2458 7836 2477
rect 7802 2409 7836 2417
rect 7802 2383 7836 2409
rect 7802 2341 7836 2342
rect 7802 2308 7836 2341
rect 7802 2239 7836 2267
rect 7802 2233 7836 2239
rect 7802 2171 7836 2192
rect 7802 2158 7836 2171
rect 7802 2103 7836 2117
rect 7802 2083 7836 2103
rect 7802 2035 7836 2042
rect 7802 2008 7836 2035
rect 7802 1933 7836 1967
rect 8018 2817 8052 2840
rect 8018 2806 8052 2817
rect 8018 2749 8052 2768
rect 8018 2734 8052 2749
rect 8018 2681 8052 2696
rect 8018 2662 8052 2681
rect 8018 2613 8052 2624
rect 8018 2590 8052 2613
rect 8018 2545 8052 2551
rect 8018 2517 8052 2545
rect 8018 2477 8052 2478
rect 8018 2444 8052 2477
rect 8018 2375 8052 2405
rect 8018 2371 8052 2375
rect 8018 2307 8052 2332
rect 8018 2298 8052 2307
rect 8018 2239 8052 2259
rect 8018 2225 8052 2239
rect 8018 2171 8052 2186
rect 8018 2152 8052 2171
rect 8018 2103 8052 2113
rect 8018 2079 8052 2103
rect 8018 2035 8052 2040
rect 8018 2006 8052 2035
rect 8018 1933 8052 1967
rect 8174 2851 8208 2867
rect 8174 2833 8208 2851
rect 8174 2783 8208 2788
rect 8174 2754 8208 2783
rect 8174 2681 8208 2709
rect 8174 2675 8208 2681
rect 8174 2613 8208 2630
rect 8174 2596 8208 2613
rect 8174 2545 8208 2551
rect 8174 2517 8208 2545
rect 8174 2443 8208 2472
rect 8174 2438 8208 2443
rect 8174 2375 8208 2393
rect 8174 2359 8208 2375
rect 8174 2307 8208 2314
rect 8174 2280 8208 2307
rect 8174 2205 8208 2234
rect 8174 2200 8208 2205
rect 8174 2137 8208 2154
rect 8174 2120 8208 2137
rect 8330 2851 8364 2867
rect 8330 2833 8364 2851
rect 8330 2783 8364 2792
rect 8330 2758 8364 2783
rect 8330 2715 8364 2717
rect 8330 2683 8364 2715
rect 8330 2613 8364 2642
rect 8330 2608 8364 2613
rect 8330 2545 8364 2567
rect 8330 2533 8364 2545
rect 8330 2477 8364 2492
rect 8330 2458 8364 2477
rect 8330 2409 8364 2417
rect 8330 2383 8364 2409
rect 8330 2341 8364 2342
rect 8330 2308 8364 2341
rect 8330 2239 8364 2267
rect 8330 2233 8364 2239
rect 8330 2171 8364 2192
rect 8330 2158 8364 2171
rect 8330 2103 8364 2117
rect 8330 2083 8364 2103
rect 8330 2035 8364 2042
rect 8330 2008 8364 2035
rect 8330 1933 8364 1967
rect 8486 2851 8520 2867
rect 8486 2833 8520 2851
rect 8486 2783 8520 2788
rect 8486 2754 8520 2783
rect 8486 2681 8520 2709
rect 8486 2675 8520 2681
rect 8486 2613 8520 2630
rect 8486 2596 8520 2613
rect 8486 2545 8520 2551
rect 8486 2517 8520 2545
rect 8486 2443 8520 2472
rect 8486 2438 8520 2443
rect 8486 2375 8520 2393
rect 8486 2359 8520 2375
rect 8486 2307 8520 2314
rect 8486 2280 8520 2307
rect 8486 2205 8520 2234
rect 8486 2200 8520 2205
rect 8486 2137 8520 2154
rect 8486 2120 8520 2137
rect 8642 2851 8676 2867
rect 8642 2833 8676 2851
rect 8642 2783 8676 2792
rect 8642 2758 8676 2783
rect 8642 2715 8676 2717
rect 8642 2683 8676 2715
rect 8642 2613 8676 2642
rect 8642 2608 8676 2613
rect 8642 2545 8676 2567
rect 8642 2533 8676 2545
rect 8642 2477 8676 2492
rect 8642 2458 8676 2477
rect 8642 2409 8676 2417
rect 8642 2383 8676 2409
rect 8642 2341 8676 2342
rect 8642 2308 8676 2341
rect 8642 2239 8676 2267
rect 8642 2233 8676 2239
rect 8642 2171 8676 2192
rect 8642 2158 8676 2171
rect 8642 2103 8676 2117
rect 8642 2083 8676 2103
rect 8642 2035 8676 2042
rect 8642 2008 8676 2035
rect 8642 1933 8676 1967
rect 8795 2870 8829 2901
rect 8795 2867 8829 2870
rect 8795 2802 8829 2827
rect 8795 2793 8829 2802
rect 8795 2734 8829 2753
rect 8795 2719 8829 2734
rect 8795 2666 8829 2679
rect 8795 2645 8829 2666
rect 8795 2598 8829 2605
rect 8795 2571 8829 2598
rect 8795 2530 8829 2531
rect 8795 2497 8829 2530
rect 8795 2428 8829 2457
rect 8795 2423 8829 2428
rect 8795 2360 8829 2383
rect 8795 2349 8829 2360
rect 8795 2292 8829 2309
rect 8795 2275 8829 2292
rect 8795 2224 8829 2235
rect 8795 2201 8829 2224
rect 8795 2156 8829 2161
rect 8795 2127 8829 2156
rect 8795 2054 8829 2086
rect 8795 2052 8829 2054
rect 8795 1986 8829 2011
rect 8795 1977 8829 1986
rect 7225 1859 7259 1879
rect 7225 1845 7259 1859
rect 8795 1918 8829 1936
rect 8795 1902 8829 1918
rect 7451 1839 7465 1873
rect 7465 1839 7485 1873
rect 7529 1839 7541 1873
rect 7541 1839 7563 1873
rect 7606 1839 7616 1873
rect 7616 1839 7640 1873
rect 7683 1839 7691 1873
rect 7691 1839 7717 1873
rect 7760 1839 7766 1873
rect 7766 1839 7794 1873
rect 7837 1839 7841 1873
rect 7841 1839 7871 1873
rect 7914 1839 7916 1873
rect 7916 1839 7948 1873
rect 8101 1839 8113 1873
rect 8113 1839 8135 1873
rect 8179 1839 8185 1873
rect 8185 1839 8213 1873
rect 8257 1839 8291 1873
rect 8335 1839 8367 1873
rect 8367 1839 8369 1873
rect 8413 1839 8439 1873
rect 8439 1839 8447 1873
rect 8490 1839 8510 1873
rect 8510 1839 8524 1873
rect 8567 1839 8581 1873
rect 8581 1839 8601 1873
rect 7225 1788 7259 1806
rect 7225 1772 7259 1788
rect 8795 1850 8829 1861
rect 8795 1827 8829 1850
rect 8795 1782 8829 1786
rect 8795 1752 8829 1782
rect 7780 1680 7803 1714
rect 7803 1680 7814 1714
rect 7853 1680 7871 1714
rect 7871 1680 7887 1714
rect 7926 1680 7939 1714
rect 7939 1680 7960 1714
rect 7999 1680 8007 1714
rect 8007 1680 8033 1714
rect 8072 1680 8075 1714
rect 8075 1680 8106 1714
rect 8145 1680 8177 1714
rect 8177 1680 8179 1714
rect 8218 1680 8245 1714
rect 8245 1680 8252 1714
rect 8291 1680 8313 1714
rect 8313 1680 8325 1714
rect 8363 1680 8381 1714
rect 8381 1680 8397 1714
rect 8435 1680 8449 1714
rect 8449 1680 8469 1714
rect 8507 1680 8517 1714
rect 8517 1680 8541 1714
rect 8579 1680 8585 1714
rect 8585 1680 8613 1714
rect 8651 1680 8653 1714
rect 8653 1680 8685 1714
rect 8723 1680 8755 1714
rect 8755 1680 8757 1714
rect 9018 3021 9052 3050
rect 9018 3016 9052 3021
rect 9018 2953 9052 2976
rect 9018 2942 9052 2953
rect 9018 2885 9052 2902
rect 9018 2868 9052 2885
rect 9018 2817 9052 2828
rect 9018 2794 9052 2817
rect 9018 2749 9052 2754
rect 9018 2720 9052 2749
rect 9018 2647 9052 2680
rect 9018 2646 9052 2647
rect 9018 2579 9052 2606
rect 9018 2572 9052 2579
rect 9018 2511 9052 2532
rect 9018 2498 9052 2511
rect 9018 2443 9052 2458
rect 9018 2424 9052 2443
rect 9018 2375 9052 2384
rect 9018 2350 9052 2375
rect 9018 2307 9052 2310
rect 9018 2276 9052 2307
rect 9018 2205 9052 2236
rect 9018 2202 9052 2205
rect 9018 2137 9052 2162
rect 9018 2128 9052 2137
rect 9018 2069 9052 2088
rect 9018 2054 9052 2069
rect 9018 2001 9052 2013
rect 9018 1979 9052 2001
rect 9018 1933 9052 1938
rect 9018 1904 9052 1933
rect 9018 1831 9052 1863
rect 9018 1829 9052 1831
rect 9018 1763 9052 1788
rect 9018 1754 9052 1763
rect 6999 1640 7033 1672
rect 6999 1638 7033 1640
rect 6999 1566 7033 1600
rect 6999 1494 7033 1528
rect 9018 1695 9052 1713
rect 9018 1679 9052 1695
rect 9588 3054 9622 3088
rect 9673 3054 9707 3088
rect 9759 3054 9793 3088
rect 9845 3054 9879 3088
rect 9931 3054 9965 3088
rect 10041 3054 10075 3088
rect 10116 3054 10150 3088
rect 10191 3054 10225 3088
rect 10266 3054 10300 3088
rect 10341 3054 10375 3088
rect 10416 3054 10450 3088
rect 10491 3054 10525 3088
rect 10566 3054 10600 3088
rect 10641 3054 10675 3088
rect 10716 3054 10750 3088
rect 10791 3054 10825 3088
rect 10866 3054 10900 3088
rect 10941 3054 10975 3088
rect 11016 3054 11050 3088
rect 11091 3054 11125 3088
rect 11167 3054 11201 3088
rect 11243 3054 11277 3088
rect 11319 3054 11353 3088
rect 11395 3054 11429 3088
rect 11471 3054 11505 3088
rect 11547 3054 11581 3088
rect 11623 3054 11657 3088
rect 9503 2982 9537 3016
rect 9503 2938 9537 2943
rect 9503 2909 9537 2938
rect 11695 2982 11729 3016
rect 9503 2836 9537 2870
rect 9503 2768 9537 2797
rect 9503 2763 9537 2768
rect 9503 2700 9537 2724
rect 9503 2690 9537 2700
rect 9503 2632 9537 2651
rect 9503 2617 9537 2632
rect 9503 2564 9537 2578
rect 9503 2544 9537 2564
rect 9503 2496 9537 2506
rect 9503 2472 9537 2496
rect 9503 2428 9537 2434
rect 9503 2400 9537 2428
rect 9503 2360 9537 2362
rect 9503 2328 9537 2360
rect 9503 2258 9537 2290
rect 9503 2256 9537 2258
rect 9503 2190 9537 2218
rect 9503 2184 9537 2190
rect 9503 2122 9537 2146
rect 9503 2112 9537 2122
rect 9503 2054 9537 2074
rect 9503 2040 9537 2054
rect 9503 1986 9537 2002
rect 9503 1968 9537 1986
rect 9503 1918 9537 1930
rect 9503 1896 9537 1918
rect 9648 2875 9682 2909
rect 9960 2875 9994 2909
rect 9648 2817 9682 2837
rect 9648 2803 9682 2817
rect 9648 2749 9682 2765
rect 9648 2731 9682 2749
rect 9648 2681 9682 2693
rect 9648 2659 9682 2681
rect 9648 2613 9682 2621
rect 9648 2587 9682 2613
rect 9648 2545 9682 2549
rect 9648 2515 9682 2545
rect 9648 2443 9682 2477
rect 9648 2375 9682 2405
rect 9648 2371 9682 2375
rect 9648 2307 9682 2332
rect 9648 2298 9682 2307
rect 9648 2239 9682 2259
rect 9648 2225 9682 2239
rect 9648 2171 9682 2186
rect 9648 2152 9682 2171
rect 9648 2103 9682 2113
rect 9648 2079 9682 2103
rect 9648 2035 9682 2040
rect 9648 2006 9682 2035
rect 9648 1933 9682 1967
rect 9803 2749 9804 2782
rect 9804 2749 9837 2782
rect 9803 2748 9837 2749
rect 9803 2681 9804 2708
rect 9804 2681 9837 2708
rect 9803 2674 9837 2681
rect 9803 2613 9804 2634
rect 9804 2613 9837 2634
rect 9803 2600 9837 2613
rect 9803 2545 9804 2560
rect 9804 2545 9837 2560
rect 9803 2526 9837 2545
rect 9803 2477 9804 2486
rect 9804 2477 9837 2486
rect 9803 2452 9837 2477
rect 9803 2409 9804 2412
rect 9804 2409 9837 2412
rect 9803 2378 9837 2409
rect 9803 2307 9837 2338
rect 9803 2304 9804 2307
rect 9804 2304 9837 2307
rect 9803 2239 9837 2264
rect 9803 2230 9804 2239
rect 9804 2230 9837 2239
rect 9803 2171 9837 2190
rect 9803 2156 9804 2171
rect 9804 2156 9837 2171
rect 9803 2103 9837 2116
rect 9803 2082 9804 2103
rect 9804 2082 9837 2103
rect 9803 2035 9837 2042
rect 9803 2008 9804 2035
rect 9804 2008 9837 2035
rect 9803 1933 9804 1967
rect 9804 1933 9837 1967
rect 10272 2875 10306 2909
rect 9960 2817 9994 2837
rect 9960 2803 9994 2817
rect 9960 2749 9994 2765
rect 9960 2731 9994 2749
rect 9960 2681 9994 2693
rect 9960 2659 9994 2681
rect 9960 2613 9994 2621
rect 9960 2587 9994 2613
rect 9960 2545 9994 2549
rect 9960 2515 9994 2545
rect 9960 2443 9994 2477
rect 9960 2375 9994 2405
rect 9960 2371 9994 2375
rect 9960 2307 9994 2332
rect 9960 2298 9994 2307
rect 9960 2239 9994 2259
rect 9960 2225 9994 2239
rect 9960 2171 9994 2186
rect 9960 2152 9994 2171
rect 9960 2103 9994 2113
rect 9960 2079 9994 2103
rect 9960 2035 9994 2040
rect 9960 2006 9994 2035
rect 9960 1933 9994 1967
rect 10116 2749 10150 2782
rect 10116 2748 10150 2749
rect 10116 2681 10150 2705
rect 10116 2671 10150 2681
rect 10116 2613 10150 2628
rect 10116 2594 10150 2613
rect 10116 2545 10150 2551
rect 10116 2517 10150 2545
rect 10116 2443 10150 2474
rect 10116 2440 10150 2443
rect 10116 2375 10150 2397
rect 10116 2363 10150 2375
rect 10116 2307 10150 2320
rect 10116 2286 10150 2307
rect 10116 2239 10150 2243
rect 10116 2209 10150 2239
rect 10116 2137 10150 2166
rect 10116 2132 10150 2137
rect 10116 2069 10150 2088
rect 10116 2054 10150 2069
rect 10584 2875 10618 2909
rect 10272 2817 10306 2837
rect 10272 2803 10306 2817
rect 10272 2749 10306 2765
rect 10272 2731 10306 2749
rect 10272 2681 10306 2693
rect 10272 2659 10306 2681
rect 10272 2613 10306 2621
rect 10272 2587 10306 2613
rect 10272 2545 10306 2549
rect 10272 2515 10306 2545
rect 10272 2443 10306 2477
rect 10272 2375 10306 2405
rect 10272 2371 10306 2375
rect 10272 2307 10306 2332
rect 10272 2298 10306 2307
rect 10272 2239 10306 2259
rect 10272 2225 10306 2239
rect 10272 2171 10306 2186
rect 10272 2152 10306 2171
rect 10272 2103 10306 2113
rect 10272 2079 10306 2103
rect 10272 2035 10306 2040
rect 10272 2006 10306 2035
rect 10272 1933 10306 1967
rect 10428 2749 10462 2782
rect 10428 2748 10462 2749
rect 10428 2681 10462 2705
rect 10428 2671 10462 2681
rect 10428 2613 10462 2628
rect 10428 2594 10462 2613
rect 10428 2545 10462 2551
rect 10428 2517 10462 2545
rect 10428 2443 10462 2474
rect 10428 2440 10462 2443
rect 10428 2375 10462 2397
rect 10428 2363 10462 2375
rect 10428 2307 10462 2320
rect 10428 2286 10462 2307
rect 10428 2239 10462 2243
rect 10428 2209 10462 2239
rect 10428 2137 10462 2166
rect 10428 2132 10462 2137
rect 10428 2069 10462 2088
rect 10428 2054 10462 2069
rect 10896 2875 10930 2909
rect 10584 2817 10618 2837
rect 10584 2803 10618 2817
rect 10584 2749 10618 2765
rect 10584 2731 10618 2749
rect 10584 2681 10618 2693
rect 10584 2659 10618 2681
rect 10584 2613 10618 2621
rect 10584 2587 10618 2613
rect 10584 2545 10618 2549
rect 10584 2515 10618 2545
rect 10584 2443 10618 2477
rect 10584 2375 10618 2405
rect 10584 2371 10618 2375
rect 10584 2307 10618 2332
rect 10584 2298 10618 2307
rect 10584 2239 10618 2259
rect 10584 2225 10618 2239
rect 10584 2171 10618 2186
rect 10584 2152 10618 2171
rect 10584 2103 10618 2113
rect 10584 2079 10618 2103
rect 10584 2035 10618 2040
rect 10584 2006 10618 2035
rect 10584 1933 10618 1967
rect 10740 2783 10774 2810
rect 10740 2776 10774 2783
rect 10740 2715 10774 2731
rect 10740 2697 10774 2715
rect 10740 2647 10774 2651
rect 10740 2617 10774 2647
rect 10740 2545 10774 2571
rect 10740 2537 10774 2545
rect 10740 2477 10774 2491
rect 10740 2457 10774 2477
rect 10740 2409 10774 2411
rect 10740 2377 10774 2409
rect 10740 2307 10774 2331
rect 10740 2297 10774 2307
rect 10740 2239 10774 2251
rect 10740 2217 10774 2239
rect 10740 2137 10774 2171
rect 10740 2069 10774 2091
rect 10740 2057 10774 2069
rect 11208 2875 11242 2909
rect 10896 2817 10930 2837
rect 10896 2803 10930 2817
rect 10896 2749 10930 2765
rect 10896 2731 10930 2749
rect 10896 2681 10930 2693
rect 10896 2659 10930 2681
rect 10896 2613 10930 2621
rect 10896 2587 10930 2613
rect 10896 2545 10930 2549
rect 10896 2515 10930 2545
rect 10896 2443 10930 2477
rect 10896 2375 10930 2405
rect 10896 2371 10930 2375
rect 10896 2307 10930 2332
rect 10896 2298 10930 2307
rect 10896 2239 10930 2259
rect 10896 2225 10930 2239
rect 10896 2171 10930 2186
rect 10896 2152 10930 2171
rect 10896 2103 10930 2113
rect 10896 2079 10930 2103
rect 10896 2035 10930 2040
rect 10896 2006 10930 2035
rect 10896 1933 10930 1967
rect 11052 2783 11086 2810
rect 11052 2776 11086 2783
rect 11052 2715 11086 2734
rect 11052 2700 11086 2715
rect 11052 2647 11086 2658
rect 11052 2624 11086 2647
rect 11052 2579 11086 2582
rect 11052 2548 11086 2579
rect 11052 2477 11086 2506
rect 11052 2472 11086 2477
rect 11052 2409 11086 2429
rect 11052 2395 11086 2409
rect 11052 2341 11086 2352
rect 11052 2318 11086 2341
rect 11052 2273 11086 2275
rect 11052 2241 11086 2273
rect 11052 2171 11086 2198
rect 11052 2164 11086 2171
rect 11052 2103 11086 2121
rect 11052 2087 11086 2103
rect 11052 2035 11086 2044
rect 11052 2010 11086 2035
rect 11052 1933 11086 1967
rect 11520 2875 11554 2909
rect 11208 2817 11242 2837
rect 11208 2803 11242 2817
rect 11208 2749 11242 2765
rect 11208 2731 11242 2749
rect 11208 2681 11242 2693
rect 11208 2659 11242 2681
rect 11208 2613 11242 2621
rect 11208 2587 11242 2613
rect 11208 2545 11242 2549
rect 11208 2515 11242 2545
rect 11208 2443 11242 2477
rect 11208 2375 11242 2405
rect 11208 2371 11242 2375
rect 11208 2307 11242 2332
rect 11208 2298 11242 2307
rect 11208 2239 11242 2259
rect 11208 2225 11242 2239
rect 11208 2171 11242 2186
rect 11208 2152 11242 2171
rect 11208 2103 11242 2113
rect 11208 2079 11242 2103
rect 11208 2035 11242 2040
rect 11208 2006 11242 2035
rect 11208 1933 11242 1967
rect 11364 2749 11398 2782
rect 11364 2748 11398 2749
rect 11364 2681 11398 2708
rect 11364 2674 11398 2681
rect 11364 2613 11398 2634
rect 11364 2600 11398 2613
rect 11364 2545 11398 2560
rect 11364 2526 11398 2545
rect 11364 2477 11398 2486
rect 11364 2452 11398 2477
rect 11364 2409 11398 2412
rect 11364 2378 11398 2409
rect 11364 2307 11398 2338
rect 11364 2304 11398 2307
rect 11364 2239 11398 2264
rect 11364 2230 11398 2239
rect 11364 2171 11398 2190
rect 11364 2156 11398 2171
rect 11364 2103 11398 2116
rect 11364 2082 11398 2103
rect 11364 2035 11398 2042
rect 11364 2008 11398 2035
rect 11364 1933 11398 1967
rect 11520 2817 11554 2837
rect 11520 2803 11554 2817
rect 11520 2749 11554 2765
rect 11520 2731 11554 2749
rect 11520 2681 11554 2693
rect 11520 2659 11554 2681
rect 11520 2613 11554 2621
rect 11520 2587 11554 2613
rect 11520 2545 11554 2549
rect 11520 2515 11554 2545
rect 11520 2443 11554 2477
rect 11520 2375 11554 2405
rect 11520 2371 11554 2375
rect 11520 2307 11554 2332
rect 11520 2298 11554 2307
rect 11520 2239 11554 2259
rect 11520 2225 11554 2239
rect 11520 2171 11554 2186
rect 11520 2152 11554 2171
rect 11520 2103 11554 2113
rect 11520 2079 11554 2103
rect 11520 2035 11554 2040
rect 11520 2006 11554 2035
rect 11520 1933 11554 1967
rect 11695 2913 11729 2944
rect 11695 2910 11729 2913
rect 11695 2845 11729 2872
rect 11695 2838 11729 2845
rect 11695 2777 11729 2800
rect 11695 2766 11729 2777
rect 11695 2709 11729 2728
rect 11695 2694 11729 2709
rect 11695 2641 11729 2656
rect 11695 2622 11729 2641
rect 11695 2573 11729 2584
rect 11695 2550 11729 2573
rect 11695 2505 11729 2512
rect 11695 2478 11729 2505
rect 11695 2437 11729 2440
rect 11695 2406 11729 2437
rect 11695 2335 11729 2368
rect 11695 2334 11729 2335
rect 11695 2267 11729 2296
rect 11695 2262 11729 2267
rect 11695 2199 11729 2224
rect 11695 2190 11729 2199
rect 11695 2131 11729 2151
rect 11695 2117 11729 2131
rect 11695 2063 11729 2078
rect 11695 2044 11729 2063
rect 11695 1995 11729 2005
rect 11695 1971 11729 1995
rect 11695 1898 11729 1932
rect 9503 1850 9537 1858
rect 9503 1824 9537 1850
rect 9711 1839 9743 1873
rect 9743 1839 9745 1873
rect 9796 1839 9804 1873
rect 9804 1839 9830 1873
rect 9881 1839 9899 1873
rect 9899 1839 9915 1873
rect 10286 1839 10318 1873
rect 10318 1839 10320 1873
rect 10362 1839 10392 1873
rect 10392 1839 10396 1873
rect 10437 1839 10466 1873
rect 10466 1839 10471 1873
rect 10512 1839 10540 1873
rect 10540 1839 10546 1873
rect 10587 1839 10614 1873
rect 10614 1839 10621 1873
rect 10662 1839 10688 1873
rect 10688 1839 10696 1873
rect 10737 1839 10762 1873
rect 10762 1839 10771 1873
rect 10812 1839 10836 1873
rect 10836 1839 10846 1873
rect 10954 1839 10957 1873
rect 10957 1839 10988 1873
rect 11047 1839 11052 1873
rect 11052 1839 11081 1873
rect 11140 1839 11147 1873
rect 11147 1839 11174 1873
rect 11271 1839 11303 1873
rect 11303 1839 11305 1873
rect 11364 1839 11398 1873
rect 11457 1839 11459 1873
rect 11459 1839 11491 1873
rect 9503 1782 9537 1786
rect 9503 1752 9537 1782
rect 11695 1828 11729 1859
rect 11695 1825 11729 1828
rect 11695 1760 11729 1786
rect 11695 1752 11729 1760
rect 9517 1680 9551 1714
rect 10278 1680 10301 1714
rect 10301 1680 10312 1714
rect 10353 1680 10369 1714
rect 10369 1680 10387 1714
rect 10428 1680 10437 1714
rect 10437 1680 10462 1714
rect 10503 1680 10505 1714
rect 10505 1680 10537 1714
rect 10578 1680 10607 1714
rect 10607 1680 10612 1714
rect 10653 1680 10675 1714
rect 10675 1680 10687 1714
rect 10728 1680 10743 1714
rect 10743 1680 10762 1714
rect 10803 1680 10811 1714
rect 10811 1680 10837 1714
rect 10878 1680 10879 1714
rect 10879 1680 10912 1714
rect 10953 1680 10981 1714
rect 10981 1680 10987 1714
rect 11028 1680 11049 1714
rect 11049 1680 11062 1714
rect 11103 1680 11117 1714
rect 11117 1680 11137 1714
rect 11177 1680 11185 1714
rect 11185 1680 11211 1714
rect 11251 1680 11253 1714
rect 11253 1680 11285 1714
rect 11325 1680 11355 1714
rect 11355 1680 11359 1714
rect 11399 1680 11423 1714
rect 11423 1680 11433 1714
rect 11473 1680 11491 1714
rect 11491 1680 11507 1714
rect 11547 1680 11559 1714
rect 11559 1680 11581 1714
rect 11621 1680 11627 1714
rect 11627 1680 11655 1714
rect 11994 3030 12028 3064
rect 12066 3030 12090 3064
rect 12090 3030 12100 3064
rect 12138 3030 12158 3064
rect 12158 3030 12172 3064
rect 12210 3030 12226 3064
rect 12226 3030 12244 3064
rect 12282 3030 12294 3064
rect 12294 3030 12316 3064
rect 12354 3030 12362 3064
rect 12362 3030 12388 3064
rect 12426 3030 12430 3064
rect 12430 3030 12460 3064
rect 12498 3030 12532 3064
rect 12570 3030 12600 3064
rect 12600 3030 12604 3064
rect 12642 3030 12668 3064
rect 12668 3030 12676 3064
rect 12714 3030 12736 3064
rect 12736 3030 12748 3064
rect 12786 3030 12804 3064
rect 12804 3030 12820 3064
rect 12858 3030 12872 3064
rect 12872 3030 12892 3064
rect 12930 3030 12940 3064
rect 12940 3030 12964 3064
rect 13002 3030 13008 3064
rect 13008 3030 13036 3064
rect 13074 3030 13076 3064
rect 13076 3030 13108 3064
rect 13146 3030 13178 3064
rect 13178 3030 13180 3064
rect 13218 3030 13246 3064
rect 13246 3030 13252 3064
rect 13290 3030 13314 3064
rect 13314 3030 13324 3064
rect 13362 3030 13382 3064
rect 13382 3030 13396 3064
rect 13434 3030 13450 3064
rect 13450 3030 13468 3064
rect 13506 3030 13518 3064
rect 13518 3030 13540 3064
rect 13578 3030 13586 3064
rect 13586 3030 13612 3064
rect 13650 3030 13654 3064
rect 13654 3030 13684 3064
rect 13722 3030 13756 3064
rect 13794 3030 13824 3064
rect 13824 3030 13828 3064
rect 13866 3030 13892 3064
rect 13892 3030 13900 3064
rect 13938 3030 13960 3064
rect 13960 3030 13972 3064
rect 14010 3030 14028 3064
rect 14028 3030 14044 3064
rect 14082 3030 14096 3064
rect 14096 3030 14116 3064
rect 14154 3030 14164 3064
rect 14164 3030 14188 3064
rect 14226 3030 14232 3064
rect 14232 3030 14260 3064
rect 14298 3030 14300 3064
rect 14300 3030 14332 3064
rect 14370 3030 14402 3064
rect 14402 3030 14404 3064
rect 14442 3030 14470 3064
rect 14470 3030 14476 3064
rect 14514 3030 14538 3064
rect 14538 3030 14548 3064
rect 14586 3030 14606 3064
rect 14606 3030 14620 3064
rect 14658 3030 14674 3064
rect 14674 3030 14692 3064
rect 14730 3030 14742 3064
rect 14742 3030 14764 3064
rect 14802 3030 14810 3064
rect 14810 3030 14836 3064
rect 14874 3030 14878 3064
rect 14878 3030 14908 3064
rect 14946 3030 14980 3064
rect 15018 3030 15048 3064
rect 15048 3030 15052 3064
rect 15090 3030 15116 3064
rect 15116 3030 15124 3064
rect 15162 3030 15184 3064
rect 15184 3030 15196 3064
rect 15234 3030 15252 3064
rect 15252 3030 15268 3064
rect 15306 3030 15320 3064
rect 15320 3030 15340 3064
rect 15378 3030 15388 3064
rect 15388 3030 15412 3064
rect 15450 3030 15456 3064
rect 15456 3030 15484 3064
rect 15522 3030 15524 3064
rect 15524 3030 15556 3064
rect 15594 3030 15626 3064
rect 15626 3030 15628 3064
rect 15666 3030 15694 3064
rect 15694 3030 15700 3064
rect 15738 3030 15762 3064
rect 15762 3030 15772 3064
rect 15810 3030 15830 3064
rect 15830 3030 15844 3064
rect 15882 3030 15898 3064
rect 15898 3030 15916 3064
rect 15954 3030 15966 3064
rect 15966 3030 15988 3064
rect 16026 3030 16034 3064
rect 16034 3030 16060 3064
rect 16098 3030 16102 3064
rect 16102 3030 16132 3064
rect 16170 3030 16204 3064
rect 16243 3030 16272 3064
rect 16272 3030 16277 3064
rect 16316 3030 16340 3064
rect 16340 3030 16350 3064
rect 16389 3030 16408 3064
rect 16408 3030 16423 3064
rect 16462 3030 16476 3064
rect 16476 3030 16496 3064
rect 16572 3030 16578 3064
rect 16578 3030 16606 3064
rect 16646 3030 16680 3064
rect 16720 3030 16748 3064
rect 16748 3030 16754 3064
rect 16794 3030 16816 3064
rect 16816 3030 16828 3064
rect 16868 3030 16884 3064
rect 16884 3030 16902 3064
rect 16942 3030 16952 3064
rect 16952 3030 16976 3064
rect 17016 3030 17020 3064
rect 17020 3030 17050 3064
rect 11922 2962 11956 2992
rect 11922 2958 11956 2962
rect 11922 2894 11956 2919
rect 11922 2885 11956 2894
rect 11922 2826 11956 2846
rect 11922 2812 11956 2826
rect 11922 2758 11956 2773
rect 11922 2739 11956 2758
rect 14535 2927 14569 2961
rect 14535 2856 14569 2887
rect 14535 2853 14569 2856
rect 12208 2744 12232 2778
rect 12232 2744 12242 2778
rect 12281 2744 12302 2778
rect 12302 2744 12315 2778
rect 12354 2744 12372 2778
rect 12372 2744 12388 2778
rect 12427 2744 12442 2778
rect 12442 2744 12461 2778
rect 12500 2744 12512 2778
rect 12512 2744 12534 2778
rect 12573 2744 12582 2778
rect 12582 2744 12607 2778
rect 12646 2744 12651 2778
rect 12651 2744 12680 2778
rect 12719 2744 12720 2778
rect 12720 2744 12753 2778
rect 12792 2744 12823 2778
rect 12823 2744 12826 2778
rect 12865 2744 12892 2778
rect 12892 2744 12899 2778
rect 12938 2744 12961 2778
rect 12961 2744 12972 2778
rect 13011 2744 13030 2778
rect 13030 2744 13045 2778
rect 13084 2744 13099 2778
rect 13099 2744 13118 2778
rect 13157 2744 13168 2778
rect 13168 2744 13191 2778
rect 13230 2744 13237 2778
rect 13237 2744 13264 2778
rect 13303 2744 13306 2778
rect 13306 2744 13337 2778
rect 13376 2744 13410 2778
rect 13449 2744 13479 2778
rect 13479 2744 13483 2778
rect 13522 2744 13548 2778
rect 13548 2744 13556 2778
rect 13595 2744 13617 2778
rect 13617 2744 13629 2778
rect 13668 2744 13686 2778
rect 13686 2744 13702 2778
rect 13741 2744 13755 2778
rect 13755 2744 13775 2778
rect 13814 2744 13824 2778
rect 13824 2744 13848 2778
rect 13887 2744 13893 2778
rect 13893 2744 13921 2778
rect 13960 2744 13962 2778
rect 13962 2744 13994 2778
rect 14032 2744 14065 2778
rect 14065 2744 14066 2778
rect 14104 2744 14134 2778
rect 14134 2744 14138 2778
rect 14176 2744 14203 2778
rect 14203 2744 14210 2778
rect 14535 2787 14569 2813
rect 14535 2779 14569 2787
rect 17088 2976 17122 2992
rect 17088 2958 17122 2976
rect 17088 2908 17122 2920
rect 17088 2886 17122 2908
rect 17088 2840 17122 2848
rect 17088 2814 17122 2840
rect 11922 2690 11956 2700
rect 11922 2666 11956 2690
rect 14896 2744 14911 2778
rect 14911 2744 14930 2778
rect 14970 2744 14981 2778
rect 14981 2744 15004 2778
rect 15044 2744 15051 2778
rect 15051 2744 15078 2778
rect 15118 2744 15121 2778
rect 15121 2744 15152 2778
rect 15192 2744 15226 2778
rect 15266 2744 15296 2778
rect 15296 2744 15300 2778
rect 15340 2744 15365 2778
rect 15365 2744 15374 2778
rect 15414 2744 15434 2778
rect 15434 2744 15448 2778
rect 15488 2744 15503 2778
rect 15503 2744 15522 2778
rect 15562 2744 15572 2778
rect 15572 2744 15596 2778
rect 15636 2744 15641 2778
rect 15641 2744 15670 2778
rect 15710 2744 15744 2778
rect 15784 2744 15813 2778
rect 15813 2744 15818 2778
rect 15858 2744 15882 2778
rect 15882 2744 15892 2778
rect 15932 2744 15951 2778
rect 15951 2744 15966 2778
rect 16006 2744 16020 2778
rect 16020 2744 16040 2778
rect 16080 2744 16089 2778
rect 16089 2744 16114 2778
rect 16154 2744 16158 2778
rect 16158 2744 16188 2778
rect 16228 2744 16262 2778
rect 16302 2744 16331 2778
rect 16331 2744 16336 2778
rect 16376 2744 16400 2778
rect 16400 2744 16410 2778
rect 16450 2744 16469 2778
rect 16469 2744 16484 2778
rect 16524 2744 16538 2778
rect 16538 2744 16558 2778
rect 16598 2744 16607 2778
rect 16607 2744 16632 2778
rect 16672 2744 16676 2778
rect 16676 2744 16706 2778
rect 16745 2744 16779 2778
rect 14535 2718 14569 2739
rect 14535 2705 14569 2718
rect 11922 2622 11956 2627
rect 11922 2593 11956 2622
rect 12252 2626 12268 2660
rect 12268 2626 12286 2660
rect 12326 2626 12336 2660
rect 12336 2626 12360 2660
rect 12400 2626 12404 2660
rect 12404 2626 12434 2660
rect 12474 2626 12506 2660
rect 12506 2626 12508 2660
rect 12548 2626 12574 2660
rect 12574 2626 12582 2660
rect 12622 2626 12642 2660
rect 12642 2626 12656 2660
rect 12696 2626 12710 2660
rect 12710 2626 12730 2660
rect 12770 2626 12778 2660
rect 12778 2626 12804 2660
rect 12844 2626 12846 2660
rect 12846 2626 12878 2660
rect 12918 2626 12948 2660
rect 12948 2626 12952 2660
rect 12992 2626 13016 2660
rect 13016 2626 13026 2660
rect 13066 2626 13084 2660
rect 13084 2626 13100 2660
rect 13140 2626 13152 2660
rect 13152 2626 13174 2660
rect 13214 2626 13220 2660
rect 13220 2626 13248 2660
rect 13288 2626 13322 2660
rect 13362 2626 13390 2660
rect 13390 2626 13396 2660
rect 13436 2626 13458 2660
rect 13458 2626 13470 2660
rect 13510 2626 13526 2660
rect 13526 2626 13544 2660
rect 13584 2626 13594 2660
rect 13594 2626 13618 2660
rect 13658 2626 13662 2660
rect 13662 2626 13692 2660
rect 13732 2626 13764 2660
rect 13764 2626 13766 2660
rect 13806 2626 13832 2660
rect 13832 2626 13840 2660
rect 13880 2626 13900 2660
rect 13900 2626 13914 2660
rect 13954 2626 13968 2660
rect 13968 2626 13988 2660
rect 14028 2626 14036 2660
rect 14036 2626 14062 2660
rect 14102 2626 14104 2660
rect 14104 2626 14136 2660
rect 14176 2626 14206 2660
rect 14206 2626 14210 2660
rect 14535 2649 14569 2665
rect 14535 2631 14569 2649
rect 17088 2772 17122 2776
rect 17088 2742 17122 2772
rect 17088 2670 17122 2704
rect 15145 2626 15150 2660
rect 15150 2626 15179 2660
rect 15218 2626 15252 2660
rect 15291 2626 15320 2660
rect 15320 2626 15325 2660
rect 15364 2626 15388 2660
rect 15388 2626 15398 2660
rect 15437 2626 15456 2660
rect 15456 2626 15471 2660
rect 15510 2626 15524 2660
rect 15524 2626 15544 2660
rect 15583 2626 15592 2660
rect 15592 2626 15617 2660
rect 15656 2626 15660 2660
rect 15660 2626 15690 2660
rect 15729 2626 15762 2660
rect 15762 2626 15763 2660
rect 15802 2626 15830 2660
rect 15830 2626 15836 2660
rect 15875 2626 15898 2660
rect 15898 2626 15909 2660
rect 15948 2626 15966 2660
rect 15966 2626 15982 2660
rect 16021 2626 16034 2660
rect 16034 2626 16055 2660
rect 16094 2626 16102 2660
rect 16102 2626 16128 2660
rect 16167 2626 16170 2660
rect 16170 2626 16201 2660
rect 16240 2626 16272 2660
rect 16272 2626 16274 2660
rect 16313 2626 16340 2660
rect 16340 2626 16347 2660
rect 16386 2626 16408 2660
rect 16408 2626 16420 2660
rect 16459 2626 16476 2660
rect 16476 2626 16493 2660
rect 16532 2626 16544 2660
rect 16544 2626 16566 2660
rect 16604 2626 16612 2660
rect 16612 2626 16638 2660
rect 16676 2626 16680 2660
rect 16680 2626 16710 2660
rect 16748 2626 16782 2660
rect 16820 2626 16850 2660
rect 16850 2626 16854 2660
rect 11922 2520 11956 2554
rect 11922 2452 11956 2481
rect 11922 2447 11956 2452
rect 14266 2565 14300 2588
rect 14266 2554 14300 2565
rect 14266 2492 14300 2508
rect 14266 2474 14300 2492
rect 11922 2384 11956 2408
rect 11922 2374 11956 2384
rect 12252 2390 12268 2424
rect 12268 2390 12286 2424
rect 12325 2390 12336 2424
rect 12336 2390 12359 2424
rect 12398 2390 12404 2424
rect 12404 2390 12432 2424
rect 12471 2390 12472 2424
rect 12472 2390 12505 2424
rect 12544 2390 12574 2424
rect 12574 2390 12578 2424
rect 12617 2390 12642 2424
rect 12642 2390 12651 2424
rect 12690 2390 12710 2424
rect 12710 2390 12724 2424
rect 12763 2390 12778 2424
rect 12778 2390 12797 2424
rect 12836 2390 12846 2424
rect 12846 2390 12870 2424
rect 12909 2390 12914 2424
rect 12914 2390 12943 2424
rect 12982 2390 13016 2424
rect 13055 2390 13084 2424
rect 13084 2390 13089 2424
rect 13128 2390 13152 2424
rect 13152 2390 13162 2424
rect 13200 2390 13220 2424
rect 13220 2390 13234 2424
rect 13272 2390 13288 2424
rect 13288 2390 13306 2424
rect 13344 2390 13356 2424
rect 13356 2390 13378 2424
rect 13416 2390 13424 2424
rect 13424 2390 13450 2424
rect 13488 2390 13492 2424
rect 13492 2390 13522 2424
rect 13560 2390 13594 2424
rect 13632 2390 13662 2424
rect 13662 2390 13666 2424
rect 13704 2390 13730 2424
rect 13730 2390 13738 2424
rect 13776 2390 13798 2424
rect 13798 2390 13810 2424
rect 13848 2390 13866 2424
rect 13866 2390 13882 2424
rect 13920 2390 13934 2424
rect 13934 2390 13954 2424
rect 14266 2419 14300 2427
rect 14266 2393 14300 2419
rect 11922 2316 11956 2335
rect 11922 2301 11956 2316
rect 11922 2248 11956 2262
rect 11922 2228 11956 2248
rect 11922 2180 11956 2189
rect 11922 2155 11956 2180
rect 14266 2312 14300 2346
rect 14266 2234 14300 2265
rect 14266 2231 14300 2234
rect 12420 2154 12438 2188
rect 12438 2154 12454 2188
rect 12494 2154 12506 2188
rect 12506 2154 12528 2188
rect 12568 2154 12574 2188
rect 12574 2154 12602 2188
rect 12642 2154 12676 2188
rect 12716 2154 12744 2188
rect 12744 2154 12750 2188
rect 12789 2154 12812 2188
rect 12812 2154 12823 2188
rect 12862 2154 12880 2188
rect 12880 2154 12896 2188
rect 12935 2154 12948 2188
rect 12948 2154 12969 2188
rect 13008 2154 13016 2188
rect 13016 2154 13042 2188
rect 13081 2154 13084 2188
rect 13084 2154 13115 2188
rect 13154 2154 13186 2188
rect 13186 2154 13188 2188
rect 13227 2154 13254 2188
rect 13254 2154 13261 2188
rect 13300 2154 13322 2188
rect 13322 2154 13334 2188
rect 13373 2154 13390 2188
rect 13390 2154 13407 2188
rect 13446 2154 13458 2188
rect 13458 2154 13480 2188
rect 13519 2154 13526 2188
rect 13526 2154 13553 2188
rect 13592 2154 13594 2188
rect 13594 2154 13626 2188
rect 13665 2154 13696 2188
rect 13696 2154 13699 2188
rect 13738 2154 13764 2188
rect 13764 2154 13772 2188
rect 13811 2154 13832 2188
rect 13832 2154 13845 2188
rect 13884 2154 13900 2188
rect 13900 2154 13918 2188
rect 13957 2154 13968 2188
rect 13968 2154 13991 2188
rect 14030 2154 14036 2188
rect 14036 2154 14064 2188
rect 14103 2154 14104 2188
rect 14104 2154 14137 2188
rect 14176 2154 14206 2188
rect 14206 2154 14210 2188
rect 14266 2161 14300 2184
rect 11922 2112 11956 2116
rect 11922 2082 11956 2112
rect 11922 2010 11956 2044
rect 11922 1942 11956 1972
rect 11922 1938 11956 1942
rect 14266 2150 14300 2161
rect 14266 2087 14300 2103
rect 14266 2069 14300 2087
rect 14266 2013 14300 2022
rect 14266 1988 14300 2013
rect 14535 2580 14569 2591
rect 14535 2557 14569 2580
rect 14535 2511 14569 2517
rect 14535 2483 14569 2511
rect 14535 2442 14569 2443
rect 14535 2409 14569 2442
rect 14535 2339 14569 2369
rect 14535 2335 14569 2339
rect 14535 2270 14569 2295
rect 14535 2261 14569 2270
rect 14535 2201 14569 2221
rect 14535 2187 14569 2201
rect 14535 2132 14569 2147
rect 14535 2113 14569 2132
rect 14535 2063 14569 2073
rect 14535 2039 14569 2063
rect 14535 1994 14569 1998
rect 14535 1964 14569 1994
rect 14780 2565 14814 2588
rect 14780 2554 14814 2565
rect 14780 2492 14814 2508
rect 14780 2474 14814 2492
rect 14780 2419 14814 2427
rect 17088 2602 17122 2632
rect 17088 2598 17122 2602
rect 17088 2534 17122 2559
rect 17088 2525 17122 2534
rect 17088 2466 17122 2486
rect 17088 2452 17122 2466
rect 14780 2393 14814 2419
rect 14896 2390 14912 2424
rect 14912 2390 14930 2424
rect 14971 2390 14980 2424
rect 14980 2390 15005 2424
rect 15046 2390 15048 2424
rect 15048 2390 15080 2424
rect 15121 2390 15150 2424
rect 15150 2390 15155 2424
rect 15196 2390 15218 2424
rect 15218 2390 15230 2424
rect 15271 2390 15286 2424
rect 15286 2390 15305 2424
rect 15346 2390 15354 2424
rect 15354 2390 15380 2424
rect 15420 2390 15422 2424
rect 15422 2390 15454 2424
rect 15494 2390 15524 2424
rect 15524 2390 15528 2424
rect 15568 2390 15592 2424
rect 15592 2390 15602 2424
rect 15642 2390 15660 2424
rect 15660 2390 15676 2424
rect 15716 2390 15728 2424
rect 15728 2390 15750 2424
rect 15790 2390 15796 2424
rect 15796 2390 15824 2424
rect 15864 2390 15898 2424
rect 15938 2390 15966 2424
rect 15966 2390 15972 2424
rect 16012 2390 16034 2424
rect 16034 2390 16046 2424
rect 16086 2390 16102 2424
rect 16102 2390 16120 2424
rect 16160 2390 16170 2424
rect 16170 2390 16194 2424
rect 16234 2390 16238 2424
rect 16238 2390 16268 2424
rect 16308 2390 16340 2424
rect 16340 2390 16342 2424
rect 16382 2390 16408 2424
rect 16408 2390 16416 2424
rect 16456 2390 16476 2424
rect 16476 2390 16490 2424
rect 16530 2390 16544 2424
rect 16544 2390 16564 2424
rect 16604 2390 16612 2424
rect 16612 2390 16638 2424
rect 14780 2312 14814 2346
rect 14780 2234 14814 2265
rect 14780 2231 14814 2234
rect 17088 2398 17122 2413
rect 17088 2379 17122 2398
rect 17088 2330 17122 2340
rect 17088 2306 17122 2330
rect 17088 2262 17122 2267
rect 17088 2233 17122 2262
rect 14780 2161 14814 2184
rect 14780 2150 14814 2161
rect 15064 2154 15082 2188
rect 15082 2154 15098 2188
rect 15138 2154 15150 2188
rect 15150 2154 15172 2188
rect 15212 2154 15218 2188
rect 15218 2154 15246 2188
rect 15286 2154 15320 2188
rect 15360 2154 15388 2188
rect 15388 2154 15394 2188
rect 15433 2154 15456 2188
rect 15456 2154 15467 2188
rect 15506 2154 15524 2188
rect 15524 2154 15540 2188
rect 15579 2154 15592 2188
rect 15592 2154 15613 2188
rect 15652 2154 15660 2188
rect 15660 2154 15686 2188
rect 15725 2154 15728 2188
rect 15728 2154 15759 2188
rect 15798 2154 15830 2188
rect 15830 2154 15832 2188
rect 15871 2154 15898 2188
rect 15898 2154 15905 2188
rect 15944 2154 15966 2188
rect 15966 2154 15978 2188
rect 16017 2154 16034 2188
rect 16034 2154 16051 2188
rect 16090 2154 16102 2188
rect 16102 2154 16124 2188
rect 16163 2154 16170 2188
rect 16170 2154 16197 2188
rect 16236 2154 16238 2188
rect 16238 2154 16270 2188
rect 16309 2154 16340 2188
rect 16340 2154 16343 2188
rect 16382 2154 16408 2188
rect 16408 2154 16416 2188
rect 16455 2154 16476 2188
rect 16476 2154 16489 2188
rect 16528 2154 16544 2188
rect 16544 2154 16562 2188
rect 16601 2154 16612 2188
rect 16612 2154 16635 2188
rect 16674 2154 16680 2188
rect 16680 2154 16708 2188
rect 16747 2154 16748 2188
rect 16748 2154 16781 2188
rect 16820 2154 16850 2188
rect 16850 2154 16854 2188
rect 14780 2087 14814 2103
rect 14780 2069 14814 2087
rect 14780 2013 14814 2022
rect 14780 1988 14814 2013
rect 17088 2160 17122 2194
rect 17088 2092 17122 2121
rect 17088 2087 17122 2092
rect 17088 2024 17122 2048
rect 17088 2014 17122 2024
rect 12252 1918 12268 1952
rect 12268 1918 12286 1952
rect 12325 1918 12336 1952
rect 12336 1918 12359 1952
rect 12398 1918 12404 1952
rect 12404 1918 12432 1952
rect 12471 1918 12472 1952
rect 12472 1918 12505 1952
rect 12544 1918 12574 1952
rect 12574 1918 12578 1952
rect 12617 1918 12642 1952
rect 12642 1918 12651 1952
rect 12690 1918 12710 1952
rect 12710 1918 12724 1952
rect 12763 1918 12778 1952
rect 12778 1918 12797 1952
rect 12836 1918 12846 1952
rect 12846 1918 12870 1952
rect 12909 1918 12914 1952
rect 12914 1918 12943 1952
rect 12982 1918 13016 1952
rect 13055 1918 13084 1952
rect 13084 1918 13089 1952
rect 13128 1918 13152 1952
rect 13152 1918 13162 1952
rect 13200 1918 13220 1952
rect 13220 1918 13234 1952
rect 13272 1918 13288 1952
rect 13288 1918 13306 1952
rect 13344 1918 13356 1952
rect 13356 1918 13378 1952
rect 13416 1918 13424 1952
rect 13424 1918 13450 1952
rect 13488 1918 13492 1952
rect 13492 1918 13522 1952
rect 13560 1918 13594 1952
rect 13632 1918 13662 1952
rect 13662 1918 13666 1952
rect 13704 1918 13730 1952
rect 13730 1918 13738 1952
rect 13776 1918 13798 1952
rect 13798 1918 13810 1952
rect 13848 1918 13866 1952
rect 13866 1918 13882 1952
rect 13920 1918 13934 1952
rect 13934 1918 13954 1952
rect 11922 1874 11956 1900
rect 11922 1866 11956 1874
rect 11922 1794 11956 1828
rect 11922 1742 11956 1756
rect 11922 1722 11956 1742
rect 14535 1890 14569 1923
rect 14535 1889 14569 1890
rect 14896 1918 14912 1952
rect 14912 1918 14930 1952
rect 14971 1918 14980 1952
rect 14980 1918 15005 1952
rect 15046 1918 15048 1952
rect 15048 1918 15080 1952
rect 15121 1918 15150 1952
rect 15150 1918 15155 1952
rect 15196 1918 15218 1952
rect 15218 1918 15230 1952
rect 15271 1918 15286 1952
rect 15286 1918 15305 1952
rect 15346 1918 15354 1952
rect 15354 1918 15380 1952
rect 15420 1918 15422 1952
rect 15422 1918 15454 1952
rect 15494 1918 15524 1952
rect 15524 1918 15528 1952
rect 15568 1918 15592 1952
rect 15592 1918 15602 1952
rect 15642 1918 15660 1952
rect 15660 1918 15676 1952
rect 15716 1918 15728 1952
rect 15728 1918 15750 1952
rect 15790 1918 15796 1952
rect 15796 1918 15824 1952
rect 15864 1918 15898 1952
rect 15938 1918 15966 1952
rect 15966 1918 15972 1952
rect 16012 1918 16034 1952
rect 16034 1918 16046 1952
rect 16086 1918 16102 1952
rect 16102 1918 16120 1952
rect 16160 1918 16170 1952
rect 16170 1918 16194 1952
rect 16234 1918 16238 1952
rect 16238 1918 16268 1952
rect 16308 1918 16340 1952
rect 16340 1918 16342 1952
rect 16382 1918 16408 1952
rect 16408 1918 16416 1952
rect 16456 1918 16476 1952
rect 16476 1918 16490 1952
rect 16530 1918 16544 1952
rect 16544 1918 16564 1952
rect 16604 1918 16612 1952
rect 16612 1918 16638 1952
rect 17088 1956 17122 1975
rect 17088 1941 17122 1956
rect 14535 1821 14569 1848
rect 14535 1814 14569 1821
rect 14535 1752 14569 1773
rect 14535 1739 14569 1752
rect 17088 1888 17122 1902
rect 17088 1868 17122 1888
rect 17088 1820 17122 1829
rect 17088 1795 17122 1820
rect 17088 1752 17122 1756
rect 17088 1722 17122 1752
rect 11994 1650 12024 1684
rect 12024 1650 12028 1684
rect 12068 1650 12092 1684
rect 12092 1650 12102 1684
rect 12142 1650 12160 1684
rect 12160 1650 12176 1684
rect 12216 1650 12228 1684
rect 12228 1650 12250 1684
rect 12290 1650 12296 1684
rect 12296 1650 12324 1684
rect 12364 1650 12398 1684
rect 12438 1650 12466 1684
rect 12466 1650 12472 1684
rect 12512 1650 12534 1684
rect 12534 1650 12546 1684
rect 12586 1650 12602 1684
rect 12602 1650 12620 1684
rect 12660 1650 12670 1684
rect 12670 1650 12694 1684
rect 12734 1650 12738 1684
rect 12738 1650 12768 1684
rect 12808 1650 12840 1684
rect 12840 1650 12842 1684
rect 12882 1650 12908 1684
rect 12908 1650 12916 1684
rect 12956 1650 12976 1684
rect 12976 1650 12990 1684
rect 13030 1650 13044 1684
rect 13044 1650 13064 1684
rect 13104 1650 13112 1684
rect 13112 1650 13138 1684
rect 13178 1650 13180 1684
rect 13180 1650 13212 1684
rect 13252 1650 13282 1684
rect 13282 1650 13286 1684
rect 13326 1650 13350 1684
rect 13350 1650 13360 1684
rect 13399 1650 13418 1684
rect 13418 1650 13433 1684
rect 13472 1650 13486 1684
rect 13486 1650 13506 1684
rect 13545 1650 13554 1684
rect 13554 1650 13579 1684
rect 13618 1650 13622 1684
rect 13622 1650 13652 1684
rect 13691 1650 13724 1684
rect 13724 1650 13725 1684
rect 13764 1650 13792 1684
rect 13792 1650 13798 1684
rect 13837 1650 13860 1684
rect 13860 1650 13871 1684
rect 13910 1650 13928 1684
rect 13928 1650 13944 1684
rect 13983 1650 13996 1684
rect 13996 1650 14017 1684
rect 14056 1650 14064 1684
rect 14064 1650 14090 1684
rect 14129 1650 14132 1684
rect 14132 1650 14163 1684
rect 14202 1650 14234 1684
rect 14234 1650 14236 1684
rect 14275 1650 14302 1684
rect 14302 1650 14309 1684
rect 14348 1650 14370 1684
rect 14370 1650 14382 1684
rect 14421 1650 14438 1684
rect 14438 1650 14455 1684
rect 14494 1650 14506 1684
rect 14506 1650 14528 1684
rect 14567 1650 14574 1684
rect 14574 1650 14601 1684
rect 14640 1650 14642 1684
rect 14642 1650 14674 1684
rect 14713 1650 14744 1684
rect 14744 1650 14747 1684
rect 14786 1650 14812 1684
rect 14812 1650 14820 1684
rect 14859 1650 14880 1684
rect 14880 1650 14893 1684
rect 14932 1650 14948 1684
rect 14948 1650 14966 1684
rect 15005 1650 15016 1684
rect 15016 1650 15039 1684
rect 15078 1650 15084 1684
rect 15084 1650 15112 1684
rect 15151 1650 15152 1684
rect 15152 1650 15185 1684
rect 15224 1650 15254 1684
rect 15254 1650 15258 1684
rect 15297 1650 15322 1684
rect 15322 1650 15331 1684
rect 15370 1650 15390 1684
rect 15390 1650 15404 1684
rect 15443 1650 15458 1684
rect 15458 1650 15477 1684
rect 15516 1650 15526 1684
rect 15526 1650 15550 1684
rect 15589 1650 15594 1684
rect 15594 1650 15623 1684
rect 15855 1650 15866 1684
rect 15866 1650 15889 1684
rect 15929 1650 15934 1684
rect 15934 1650 15963 1684
rect 16003 1650 16036 1684
rect 16036 1650 16037 1684
rect 16077 1650 16104 1684
rect 16104 1650 16111 1684
rect 16151 1650 16172 1684
rect 16172 1650 16185 1684
rect 16225 1650 16240 1684
rect 16240 1650 16259 1684
rect 16299 1650 16308 1684
rect 16308 1650 16333 1684
rect 16373 1650 16376 1684
rect 16376 1650 16407 1684
rect 16447 1650 16478 1684
rect 16478 1650 16481 1684
rect 16521 1650 16546 1684
rect 16546 1650 16555 1684
rect 16595 1650 16614 1684
rect 16614 1650 16629 1684
rect 16668 1650 16682 1684
rect 16682 1650 16702 1684
rect 16741 1650 16750 1684
rect 16750 1650 16775 1684
rect 16814 1650 16818 1684
rect 16818 1650 16848 1684
rect 16887 1650 16920 1684
rect 16920 1650 16921 1684
rect 16960 1650 16988 1684
rect 16988 1650 16994 1684
rect 9018 1627 9052 1638
rect 9018 1604 9052 1627
rect 9018 1559 9052 1563
rect 9018 1529 9052 1559
rect 7799 1457 7815 1491
rect 7815 1457 7833 1491
rect 7876 1457 7883 1491
rect 7883 1457 7910 1491
rect 7953 1457 7985 1491
rect 7985 1457 7987 1491
rect 8030 1457 8053 1491
rect 8053 1457 8064 1491
rect 8106 1457 8121 1491
rect 8121 1457 8140 1491
rect 8182 1457 8189 1491
rect 8189 1457 8216 1491
rect 8258 1457 8291 1491
rect 8291 1457 8292 1491
rect 8334 1457 8359 1491
rect 8359 1457 8368 1491
rect 8410 1457 8427 1491
rect 8427 1457 8444 1491
rect 8486 1457 8495 1491
rect 8495 1457 8520 1491
rect 8562 1457 8563 1491
rect 8563 1457 8596 1491
rect 8638 1457 8665 1491
rect 8665 1457 8672 1491
rect 8714 1457 8733 1491
rect 8733 1457 8748 1491
rect 8790 1457 8801 1491
rect 8801 1457 8824 1491
rect 8866 1457 8869 1491
rect 8869 1457 8900 1491
rect 8942 1457 8976 1491
rect 5910 1387 5944 1421
rect 6000 1387 6034 1421
rect 6091 1387 6125 1421
rect 6738 1196 6753 1230
rect 6753 1196 6772 1230
rect 6810 1196 6814 1230
rect 6814 1196 6844 1230
rect 7029 1196 7031 1230
rect 7031 1196 7063 1230
rect 7101 1196 7133 1230
rect 7133 1196 7135 1230
rect 7221 1196 7255 1230
rect 7293 1196 7297 1230
rect 7297 1196 7327 1230
rect 7592 1196 7597 1230
rect 7597 1196 7626 1230
rect 7668 1196 7699 1230
rect 7699 1196 7702 1230
rect 7744 1196 7767 1230
rect 7767 1196 7778 1230
rect 7820 1196 7835 1230
rect 7835 1196 7854 1230
rect 7896 1196 7903 1230
rect 7903 1196 7930 1230
rect 7972 1196 8005 1230
rect 8005 1196 8006 1230
rect 8048 1196 8073 1230
rect 8073 1196 8082 1230
rect 8124 1196 8141 1230
rect 8141 1196 8158 1230
rect 8200 1196 8210 1230
rect 8210 1196 8234 1230
rect 8276 1196 8279 1230
rect 8279 1196 8310 1230
rect 8383 1196 8417 1230
rect 8521 1196 8555 1230
rect 9705 1196 9733 1230
rect 9733 1196 9739 1230
rect 9780 1196 9802 1230
rect 9802 1196 9814 1230
rect 9855 1196 9871 1230
rect 9871 1196 9889 1230
rect 9930 1196 9940 1230
rect 9940 1196 9964 1230
rect 10005 1196 10009 1230
rect 10009 1196 10039 1230
rect 10080 1196 10112 1230
rect 10112 1196 10114 1230
rect 10155 1196 10181 1230
rect 10181 1196 10189 1230
rect 10230 1196 10250 1230
rect 10250 1196 10264 1230
rect 10305 1196 10319 1230
rect 10319 1196 10339 1230
rect 10380 1196 10388 1230
rect 10388 1196 10414 1230
rect 10455 1196 10457 1230
rect 10457 1196 10489 1230
rect 10530 1196 10561 1230
rect 10561 1196 10564 1230
rect 10605 1196 10630 1230
rect 10630 1196 10639 1230
rect 10680 1196 10699 1230
rect 10699 1196 10714 1230
rect 10755 1196 10768 1230
rect 10768 1196 10789 1230
rect 10830 1196 10837 1230
rect 10837 1196 10864 1230
rect 10905 1196 10906 1230
rect 10906 1196 10939 1230
rect 10980 1196 11009 1230
rect 11009 1196 11014 1230
rect 11055 1196 11078 1230
rect 11078 1196 11089 1230
rect 11257 1196 11269 1230
rect 11269 1196 11291 1230
rect 11330 1196 11337 1230
rect 11337 1196 11364 1230
rect 11403 1196 11405 1230
rect 11405 1196 11437 1230
rect 11476 1196 11507 1230
rect 11507 1196 11510 1230
rect 11549 1196 11575 1230
rect 11575 1196 11583 1230
rect 11622 1196 11643 1230
rect 11643 1196 11656 1230
rect 11695 1196 11711 1230
rect 11711 1196 11729 1230
rect 11768 1196 11779 1230
rect 11779 1196 11802 1230
rect 11841 1196 11847 1230
rect 11847 1196 11875 1230
rect 11914 1196 11915 1230
rect 11915 1196 11948 1230
rect 11987 1196 12017 1230
rect 12017 1196 12021 1230
rect 12060 1196 12085 1230
rect 12085 1196 12094 1230
rect 12133 1196 12153 1230
rect 12153 1196 12167 1230
rect 12206 1196 12221 1230
rect 12221 1196 12240 1230
rect 12279 1196 12289 1230
rect 12289 1196 12313 1230
rect 12352 1196 12357 1230
rect 12357 1196 12386 1230
rect 12425 1196 12459 1230
rect 12498 1196 12527 1230
rect 12527 1196 12532 1230
rect 12571 1196 12595 1230
rect 12595 1196 12605 1230
rect 12644 1196 12663 1230
rect 12663 1196 12678 1230
rect 12717 1196 12731 1230
rect 12731 1196 12751 1230
rect 12790 1196 12799 1230
rect 12799 1196 12824 1230
rect 12863 1196 12867 1230
rect 12867 1196 12897 1230
rect 12936 1196 12969 1230
rect 12969 1196 12970 1230
rect 13009 1196 13037 1230
rect 13037 1196 13043 1230
rect 13082 1196 13105 1230
rect 13105 1196 13116 1230
rect 13155 1196 13173 1230
rect 13173 1196 13189 1230
rect 13228 1196 13241 1230
rect 13241 1196 13262 1230
rect 13301 1196 13310 1230
rect 13310 1196 13335 1230
rect 13374 1196 13379 1230
rect 13379 1196 13408 1230
rect 13447 1196 13448 1230
rect 13448 1196 13481 1230
rect 13520 1196 13552 1230
rect 13552 1196 13554 1230
rect 13593 1196 13621 1230
rect 13621 1196 13627 1230
rect 13666 1196 13690 1230
rect 13690 1196 13700 1230
rect 13739 1196 13759 1230
rect 13759 1196 13773 1230
rect 13812 1196 13828 1230
rect 13828 1196 13846 1230
rect 13885 1196 13897 1230
rect 13897 1196 13919 1230
rect 13958 1196 13966 1230
rect 13966 1196 13992 1230
rect 14031 1196 14035 1230
rect 14035 1196 14065 1230
rect 14104 1196 14138 1230
rect 14177 1196 14207 1230
rect 14207 1196 14211 1230
rect 14250 1196 14276 1230
rect 14276 1196 14284 1230
rect 14323 1196 14345 1230
rect 14345 1196 14357 1230
rect 14396 1196 14414 1230
rect 14414 1196 14430 1230
rect 14469 1196 14483 1230
rect 14483 1196 14503 1230
rect 14542 1196 14552 1230
rect 14552 1196 14576 1230
rect 14615 1196 14621 1230
rect 14621 1196 14649 1230
rect 14688 1196 14690 1230
rect 14690 1196 14722 1230
rect 14761 1196 14794 1230
rect 14794 1196 14795 1230
rect 14833 1196 14863 1230
rect 14863 1196 14867 1230
rect 14905 1196 14932 1230
rect 14932 1196 14939 1230
rect 14977 1196 15001 1230
rect 15001 1196 15011 1230
rect 15252 1196 15267 1230
rect 15267 1196 15286 1230
rect 15369 1196 15401 1230
rect 15401 1196 15403 1230
rect 15829 1196 15832 1230
rect 15832 1196 15863 1230
rect 15913 1196 15943 1230
rect 15943 1196 15947 1230
rect 1613 1032 1622 1066
rect 1622 1032 1647 1066
rect 1689 1032 1690 1066
rect 1690 1032 1723 1066
rect 1765 1032 1792 1066
rect 1792 1032 1799 1066
rect 1841 1032 1860 1066
rect 1860 1032 1875 1066
rect 1917 1032 1928 1066
rect 1928 1032 1951 1066
rect 1993 1032 1996 1066
rect 1996 1032 2027 1066
rect 2069 1032 2098 1066
rect 2098 1032 2103 1066
rect 2145 1032 2166 1066
rect 2166 1032 2179 1066
rect 2221 1032 2234 1066
rect 2234 1032 2255 1066
rect 2296 1032 2302 1066
rect 2302 1032 2330 1066
rect 2966 1034 3000 1068
rect 3049 1066 3083 1068
rect 3132 1066 3166 1068
rect 3215 1066 3249 1068
rect 3299 1066 3333 1068
rect 3383 1066 3417 1068
rect 3049 1034 3057 1066
rect 3057 1034 3083 1066
rect 3132 1034 3159 1066
rect 3159 1034 3166 1066
rect 3215 1034 3227 1066
rect 3227 1034 3249 1066
rect 3299 1034 3329 1066
rect 3329 1034 3333 1066
rect 3383 1034 3397 1066
rect 3397 1034 3417 1066
rect 3942 1010 3976 1019
rect 3942 985 3976 1010
rect 3942 942 3976 946
rect 3942 912 3976 942
rect 3942 840 3976 873
rect 3942 839 3976 840
rect 2260 792 2294 826
rect 2260 720 2294 754
rect 3172 797 3206 831
rect 3172 725 3206 759
rect 3942 772 3976 800
rect 3942 766 3976 772
rect 3942 704 3976 727
rect 3942 693 3976 704
rect 3942 636 3976 654
rect 3942 620 3976 636
rect 3942 568 3976 581
rect 3942 547 3976 568
rect 3942 500 3976 507
rect 3942 473 3976 500
rect 1685 414 1719 448
rect 1895 422 1929 456
rect 1685 342 1719 376
rect 1789 365 1823 399
rect 1895 349 1929 383
rect 2151 415 2185 449
rect 2151 343 2185 377
rect 3085 421 3119 455
rect 3085 349 3119 383
rect 3257 424 3291 458
rect 3257 352 3291 386
rect 3942 432 3976 433
rect 3942 399 3976 432
rect 1789 293 1823 327
rect 3942 330 3976 359
rect 3942 325 3976 330
rect 3942 262 3976 285
rect 3942 251 3976 262
rect 4048 1078 4082 1082
rect 4048 1048 4082 1078
rect 4048 976 4082 1010
rect 4048 908 4082 938
rect 4048 904 4082 908
rect 4048 840 4082 866
rect 4048 832 4082 840
rect 4048 772 4082 794
rect 4048 760 4082 772
rect 4048 704 4082 722
rect 4048 688 4082 704
rect 4048 636 4082 650
rect 4048 616 4082 636
rect 4048 568 4082 577
rect 4048 543 4082 568
rect 4048 500 4082 504
rect 4048 470 4082 500
rect 4048 398 4082 431
rect 4048 397 4082 398
rect 4048 330 4082 358
rect 4048 324 4082 330
rect 4048 262 4082 285
rect 4048 251 4082 262
rect 4154 1078 4188 1082
rect 4154 1048 4188 1078
rect 4154 976 4188 1010
rect 4154 908 4188 938
rect 4154 904 4188 908
rect 4154 840 4188 866
rect 4154 832 4188 840
rect 4154 772 4188 794
rect 4154 760 4188 772
rect 4154 704 4188 722
rect 4154 688 4188 704
rect 4154 636 4188 650
rect 4154 616 4188 636
rect 4154 568 4188 577
rect 4154 543 4188 568
rect 4154 500 4188 504
rect 4154 470 4188 500
rect 4154 398 4188 431
rect 4154 397 4188 398
rect 4154 330 4188 358
rect 4154 324 4188 330
rect 4154 262 4188 285
rect 4154 251 4188 262
rect 4260 1078 4294 1082
rect 4260 1048 4294 1078
rect 4260 976 4294 1010
rect 4260 908 4294 938
rect 4260 904 4294 908
rect 4260 840 4294 866
rect 4260 832 4294 840
rect 4260 772 4294 794
rect 4260 760 4294 772
rect 4260 704 4294 722
rect 4260 688 4294 704
rect 4260 636 4294 650
rect 4260 616 4294 636
rect 4260 568 4294 577
rect 4260 543 4294 568
rect 4260 500 4294 504
rect 4260 470 4294 500
rect 4260 398 4294 431
rect 4260 397 4294 398
rect 4260 330 4294 358
rect 4260 324 4294 330
rect 4260 262 4294 285
rect 4260 251 4294 262
rect 4366 1078 4400 1082
rect 4366 1048 4400 1078
rect 4366 976 4400 1010
rect 4366 908 4400 938
rect 4366 904 4400 908
rect 4366 840 4400 866
rect 4366 832 4400 840
rect 4366 772 4400 794
rect 4366 760 4400 772
rect 4366 704 4400 722
rect 4366 688 4400 704
rect 4366 636 4400 650
rect 4366 616 4400 636
rect 4366 568 4400 577
rect 4366 543 4400 568
rect 4366 500 4400 504
rect 4366 470 4400 500
rect 4366 398 4400 431
rect 4366 397 4400 398
rect 4366 330 4400 358
rect 4366 324 4400 330
rect 4366 262 4400 285
rect 4366 251 4400 262
rect 4472 1078 4506 1082
rect 4472 1048 4506 1078
rect 4472 976 4506 1010
rect 4472 908 4506 938
rect 4472 904 4506 908
rect 4472 840 4506 866
rect 4472 832 4506 840
rect 4472 772 4506 794
rect 4472 760 4506 772
rect 4472 704 4506 722
rect 4472 688 4506 704
rect 4472 636 4506 650
rect 4472 616 4506 636
rect 4472 568 4506 577
rect 4472 543 4506 568
rect 4472 500 4506 504
rect 4472 470 4506 500
rect 4472 398 4506 431
rect 4472 397 4506 398
rect 4472 330 4506 358
rect 4472 324 4506 330
rect 4472 262 4506 285
rect 4472 251 4506 262
rect 4578 1078 4612 1082
rect 4578 1048 4612 1078
rect 4578 976 4612 1010
rect 4578 908 4612 938
rect 4578 904 4612 908
rect 4578 840 4612 866
rect 4578 832 4612 840
rect 4578 772 4612 794
rect 4578 760 4612 772
rect 4578 704 4612 722
rect 4578 688 4612 704
rect 4578 636 4612 650
rect 4578 616 4612 636
rect 4578 568 4612 577
rect 4578 543 4612 568
rect 4578 500 4612 504
rect 4578 470 4612 500
rect 4578 398 4612 431
rect 4578 397 4612 398
rect 4578 330 4612 358
rect 4578 324 4612 330
rect 4578 262 4612 285
rect 4578 251 4612 262
rect 4684 1078 4718 1082
rect 4684 1048 4718 1078
rect 4684 976 4718 1010
rect 4684 908 4718 938
rect 4684 904 4718 908
rect 4684 840 4718 866
rect 4684 832 4718 840
rect 4684 772 4718 794
rect 4684 760 4718 772
rect 4684 704 4718 722
rect 4684 688 4718 704
rect 4684 636 4718 650
rect 4684 616 4718 636
rect 4684 568 4718 577
rect 4684 543 4718 568
rect 4684 500 4718 504
rect 4684 470 4718 500
rect 4684 398 4718 431
rect 4684 397 4718 398
rect 4684 330 4718 358
rect 4684 324 4718 330
rect 4684 262 4718 285
rect 4684 251 4718 262
rect 4790 1078 4824 1082
rect 4790 1048 4824 1078
rect 4790 976 4824 1010
rect 4790 908 4824 938
rect 4790 904 4824 908
rect 4790 840 4824 866
rect 4790 832 4824 840
rect 4790 772 4824 794
rect 4790 760 4824 772
rect 4790 704 4824 722
rect 4790 688 4824 704
rect 4790 636 4824 650
rect 4790 616 4824 636
rect 4790 568 4824 577
rect 4790 543 4824 568
rect 4790 500 4824 504
rect 4790 470 4824 500
rect 4790 398 4824 431
rect 4790 397 4824 398
rect 4790 330 4824 358
rect 4790 324 4824 330
rect 4790 262 4824 285
rect 4790 251 4824 262
rect 4896 1078 4930 1082
rect 4896 1048 4930 1078
rect 4896 976 4930 1010
rect 4896 908 4930 938
rect 4896 904 4930 908
rect 4896 840 4930 866
rect 4896 832 4930 840
rect 4896 772 4930 794
rect 4896 760 4930 772
rect 4896 704 4930 722
rect 4896 688 4930 704
rect 4896 636 4930 650
rect 4896 616 4930 636
rect 4896 568 4930 577
rect 4896 543 4930 568
rect 4896 500 4930 504
rect 4896 470 4930 500
rect 4896 398 4930 431
rect 4896 397 4930 398
rect 4896 330 4930 358
rect 4896 324 4930 330
rect 4896 262 4930 285
rect 4896 251 4930 262
rect 5002 1078 5036 1082
rect 5002 1048 5036 1078
rect 5002 976 5036 1010
rect 5002 908 5036 938
rect 5002 904 5036 908
rect 5002 840 5036 866
rect 5002 832 5036 840
rect 5002 772 5036 794
rect 5002 760 5036 772
rect 5002 704 5036 722
rect 5002 688 5036 704
rect 5002 636 5036 650
rect 5002 616 5036 636
rect 5002 568 5036 577
rect 5002 543 5036 568
rect 5002 500 5036 504
rect 5002 470 5036 500
rect 5002 398 5036 431
rect 5002 397 5036 398
rect 5002 330 5036 358
rect 5002 324 5036 330
rect 5002 262 5036 285
rect 5002 251 5036 262
rect 5108 1078 5142 1082
rect 5108 1048 5142 1078
rect 5108 976 5142 1010
rect 5108 908 5142 938
rect 5108 904 5142 908
rect 5108 840 5142 866
rect 5108 832 5142 840
rect 5108 772 5142 794
rect 5108 760 5142 772
rect 5108 704 5142 722
rect 5108 688 5142 704
rect 5108 636 5142 650
rect 5108 616 5142 636
rect 5108 568 5142 577
rect 5108 543 5142 568
rect 5108 500 5142 504
rect 5108 470 5142 500
rect 5108 398 5142 431
rect 5108 397 5142 398
rect 5108 330 5142 358
rect 5108 324 5142 330
rect 5108 262 5142 285
rect 5108 251 5142 262
rect 5214 1078 5248 1082
rect 5214 1048 5248 1078
rect 5214 976 5248 1010
rect 5214 908 5248 938
rect 5214 904 5248 908
rect 5214 840 5248 866
rect 5214 832 5248 840
rect 5214 772 5248 794
rect 5214 760 5248 772
rect 5214 704 5248 722
rect 5214 688 5248 704
rect 5214 636 5248 650
rect 5214 616 5248 636
rect 5214 568 5248 577
rect 5214 543 5248 568
rect 5214 500 5248 504
rect 5214 470 5248 500
rect 5214 398 5248 431
rect 5214 397 5248 398
rect 5214 330 5248 358
rect 5214 324 5248 330
rect 5214 262 5248 285
rect 5214 251 5248 262
rect 5320 1078 5354 1082
rect 5320 1048 5354 1078
rect 5320 976 5354 1010
rect 5320 908 5354 938
rect 5320 904 5354 908
rect 5320 840 5354 866
rect 5320 832 5354 840
rect 5320 772 5354 794
rect 5320 760 5354 772
rect 5320 704 5354 722
rect 5320 688 5354 704
rect 5320 636 5354 650
rect 5320 616 5354 636
rect 5320 568 5354 577
rect 5320 543 5354 568
rect 5320 500 5354 504
rect 5320 470 5354 500
rect 5320 398 5354 431
rect 5320 397 5354 398
rect 5320 330 5354 358
rect 5320 324 5354 330
rect 5320 262 5354 285
rect 5320 251 5354 262
rect 5426 1078 5460 1082
rect 5426 1048 5460 1078
rect 5426 976 5460 1010
rect 5426 908 5460 938
rect 5426 904 5460 908
rect 5426 840 5460 866
rect 5426 832 5460 840
rect 5426 772 5460 794
rect 5426 760 5460 772
rect 5426 704 5460 722
rect 5426 688 5460 704
rect 5426 636 5460 650
rect 5426 616 5460 636
rect 5426 568 5460 577
rect 5426 543 5460 568
rect 5426 500 5460 504
rect 5426 470 5460 500
rect 5426 398 5460 431
rect 5426 397 5460 398
rect 5426 330 5460 358
rect 5426 324 5460 330
rect 5426 262 5460 285
rect 5426 251 5460 262
rect 5532 1078 5566 1082
rect 5532 1048 5566 1078
rect 5532 976 5566 1010
rect 5532 908 5566 938
rect 5532 904 5566 908
rect 5532 840 5566 866
rect 5532 832 5566 840
rect 5532 772 5566 794
rect 5532 760 5566 772
rect 5532 704 5566 722
rect 5532 688 5566 704
rect 5532 636 5566 650
rect 5532 616 5566 636
rect 5532 568 5566 577
rect 5532 543 5566 568
rect 5532 500 5566 504
rect 5532 470 5566 500
rect 5532 398 5566 431
rect 5532 397 5566 398
rect 5532 330 5566 358
rect 5532 324 5566 330
rect 5532 262 5566 285
rect 5532 251 5566 262
rect 5638 1078 5672 1082
rect 5638 1048 5672 1078
rect 5638 976 5672 1010
rect 5900 1028 5934 1054
rect 5900 1020 5934 1028
rect 5900 960 5934 982
rect 5900 948 5934 960
rect 6116 1130 6150 1146
rect 6116 1112 6150 1130
rect 6116 1062 6150 1074
rect 6116 1040 6150 1062
rect 6548 1130 6582 1146
rect 6548 1112 6582 1130
rect 6548 1062 6582 1074
rect 6333 1028 6366 1054
rect 6366 1028 6367 1054
rect 6333 1020 6367 1028
rect 6333 960 6366 982
rect 6366 960 6367 982
rect 6333 948 6367 960
rect 6548 1040 6582 1062
rect 6658 1070 6692 1100
rect 6658 1066 6692 1070
rect 6658 1002 6692 1027
rect 6658 993 6692 1002
rect 5638 908 5672 938
rect 5638 904 5672 908
rect 6658 934 6692 954
rect 6658 920 6692 934
rect 5957 866 5961 900
rect 5961 866 5991 900
rect 6040 866 6071 900
rect 6071 866 6074 900
rect 6123 866 6146 900
rect 6146 866 6157 900
rect 6206 866 6221 900
rect 6221 866 6240 900
rect 6289 866 6296 900
rect 6296 866 6323 900
rect 6372 866 6406 900
rect 6455 866 6487 900
rect 6487 866 6489 900
rect 6658 866 6692 880
rect 5638 840 5672 866
rect 5638 832 5672 840
rect 6658 846 6692 866
rect 5638 772 5672 794
rect 5638 760 5672 772
rect 5638 704 5672 722
rect 5638 688 5672 704
rect 5638 636 5672 650
rect 5638 616 5672 636
rect 5900 800 5934 804
rect 5900 770 5934 800
rect 5900 698 5934 732
rect 6116 698 6150 712
rect 6116 678 6150 698
rect 6116 630 6150 640
rect 6116 606 6150 630
rect 6333 800 6367 804
rect 6333 770 6366 800
rect 6366 770 6367 800
rect 6333 698 6366 732
rect 6366 698 6367 732
rect 6548 698 6582 712
rect 6548 678 6582 698
rect 6548 630 6582 640
rect 6548 606 6582 630
rect 6658 798 6692 806
rect 6658 772 6692 798
rect 6658 730 6692 732
rect 6658 698 6692 730
rect 6658 628 6692 658
rect 6658 624 6692 628
rect 5638 568 5672 577
rect 5638 543 5672 568
rect 6658 560 6692 584
rect 6658 550 6692 560
rect 5638 500 5672 504
rect 5638 470 5672 500
rect 5957 494 5961 528
rect 5961 494 5991 528
rect 6040 494 6071 528
rect 6071 494 6074 528
rect 6123 494 6146 528
rect 6146 494 6157 528
rect 6206 494 6221 528
rect 6221 494 6240 528
rect 6289 494 6296 528
rect 6296 494 6323 528
rect 6372 494 6406 528
rect 6455 494 6487 528
rect 6487 494 6489 528
rect 6814 1070 6848 1100
rect 6814 1066 6848 1070
rect 6814 1002 6848 1020
rect 6814 986 6848 1002
rect 6814 934 6848 940
rect 6814 906 6848 934
rect 6814 832 6848 859
rect 6814 825 6848 832
rect 6814 764 6848 778
rect 6814 744 6848 764
rect 6814 696 6848 697
rect 6814 663 6848 696
rect 6814 594 6848 616
rect 6814 582 6848 594
rect 6970 968 7004 986
rect 6970 952 7004 968
rect 6970 900 7004 908
rect 6970 874 7004 900
rect 6970 798 7004 830
rect 6970 796 7004 798
rect 6970 730 7004 752
rect 6970 718 7004 730
rect 6970 662 7004 674
rect 6970 640 7004 662
rect 6970 594 7004 595
rect 6970 561 7004 594
rect 6658 476 6692 510
rect 5638 398 5672 431
rect 5638 397 5672 398
rect 5638 330 5672 358
rect 5638 324 5672 330
rect 5638 262 5672 285
rect 5638 251 5672 262
rect 5900 434 5934 450
rect 5900 416 5934 434
rect 5900 366 5934 378
rect 5900 344 5934 366
rect 6116 332 6150 358
rect 6116 324 6150 332
rect 6116 264 6150 286
rect 6116 252 6150 264
rect 6332 434 6366 450
rect 6332 416 6366 434
rect 6332 366 6366 378
rect 6332 344 6366 366
rect 6658 402 6692 436
rect 7126 1070 7160 1100
rect 7126 1066 7160 1070
rect 7126 1002 7160 1020
rect 7126 986 7160 1002
rect 7126 934 7160 940
rect 7126 906 7160 934
rect 7126 832 7160 859
rect 7126 825 7160 832
rect 7126 764 7160 778
rect 7126 744 7160 764
rect 7126 696 7160 697
rect 7126 663 7160 696
rect 7126 594 7160 616
rect 7126 582 7160 594
rect 7236 976 7270 986
rect 7236 952 7270 976
rect 7236 908 7270 912
rect 7236 878 7270 908
rect 7236 806 7270 838
rect 7236 804 7270 806
rect 7236 738 7270 764
rect 7236 730 7270 738
rect 7236 670 7270 690
rect 7236 656 7270 670
rect 7236 602 7270 616
rect 7236 582 7270 602
rect 6970 482 7004 516
rect 6970 403 7004 437
rect 7236 534 7270 541
rect 7236 507 7270 534
rect 7236 432 7270 466
rect 6548 332 6582 358
rect 6548 324 6582 332
rect 6548 264 6582 286
rect 6548 252 6582 264
rect 7236 364 7270 391
rect 7236 357 7270 364
rect 7236 296 7270 316
rect 7236 282 7270 296
rect 7236 228 7270 241
rect 7236 207 7270 228
rect 7236 160 7270 166
rect 7236 132 7270 160
rect 7392 1078 7426 1082
rect 7392 1048 7426 1078
rect 7392 976 7426 1004
rect 7392 970 7426 976
rect 7392 908 7426 926
rect 7392 892 7426 908
rect 7392 840 7426 848
rect 7392 814 7426 840
rect 7392 738 7426 770
rect 7392 736 7426 738
rect 7392 670 7426 692
rect 7392 658 7426 670
rect 7392 602 7426 614
rect 7392 580 7426 602
rect 7392 534 7426 536
rect 7392 502 7426 534
rect 7392 432 7426 458
rect 7392 424 7426 432
rect 7392 364 7426 380
rect 7392 346 7426 364
rect 7392 296 7426 301
rect 7392 267 7426 296
rect 7392 194 7426 222
rect 7392 188 7426 194
rect 7502 1078 7536 1094
rect 7502 1060 7536 1078
rect 7502 1010 7536 1019
rect 7502 985 7536 1010
rect 7502 942 7536 944
rect 7502 910 7536 942
rect 7502 840 7536 869
rect 7502 835 7536 840
rect 7502 772 7536 794
rect 7502 760 7536 772
rect 7502 704 7536 719
rect 7502 685 7536 704
rect 7502 636 7536 644
rect 7502 610 7536 636
rect 7502 568 7536 569
rect 7502 535 7536 568
rect 7502 466 7536 494
rect 7502 460 7536 466
rect 7502 398 7536 419
rect 7502 385 7536 398
rect 7502 330 7536 344
rect 7502 310 7536 330
rect 7502 262 7536 269
rect 7502 235 7536 262
rect 7502 160 7536 194
rect 7718 976 7752 1008
rect 7718 974 7752 976
rect 7718 908 7752 934
rect 7718 900 7752 908
rect 7718 840 7752 860
rect 7718 826 7752 840
rect 7718 772 7752 786
rect 7718 752 7752 772
rect 7718 704 7752 712
rect 7718 678 7752 704
rect 7718 636 7752 638
rect 7718 604 7752 636
rect 7718 534 7752 564
rect 7718 530 7752 534
rect 7718 466 7752 490
rect 7718 456 7752 466
rect 7718 398 7752 416
rect 7718 382 7752 398
rect 7718 330 7752 342
rect 7718 308 7752 330
rect 7718 262 7752 268
rect 7718 234 7752 262
rect 7718 160 7752 194
rect 7934 1078 7968 1094
rect 7934 1060 7968 1078
rect 7934 1010 7968 1019
rect 7934 985 7968 1010
rect 7934 942 7968 944
rect 7934 910 7968 942
rect 7934 840 7968 869
rect 7934 835 7968 840
rect 7934 772 7968 794
rect 7934 760 7968 772
rect 7934 704 7968 719
rect 7934 685 7968 704
rect 7934 636 7968 644
rect 7934 610 7968 636
rect 7934 568 7968 569
rect 7934 535 7968 568
rect 7934 466 7968 494
rect 7934 460 7968 466
rect 7934 398 7968 419
rect 7934 385 7968 398
rect 7934 330 7968 344
rect 7934 310 7968 330
rect 7934 262 7968 269
rect 7934 235 7968 262
rect 7934 160 7968 194
rect 8150 874 8184 886
rect 8150 852 8184 874
rect 8150 806 8184 810
rect 8150 776 8184 806
rect 8150 704 8184 733
rect 8150 699 8184 704
rect 8150 636 8184 656
rect 8150 622 8184 636
rect 8150 568 8184 579
rect 8150 545 8184 568
rect 8150 500 8184 502
rect 8150 468 8184 500
rect 8150 398 8184 425
rect 8150 391 8184 398
rect 8150 330 8184 348
rect 8150 314 8184 330
rect 8150 262 8184 271
rect 8150 237 8184 262
rect 8150 160 8184 194
rect 8366 1078 8400 1094
rect 8366 1060 8400 1078
rect 8366 1010 8400 1019
rect 8366 985 8400 1010
rect 8366 942 8400 944
rect 8366 910 8400 942
rect 8366 840 8400 869
rect 8366 835 8400 840
rect 8366 772 8400 794
rect 8366 760 8400 772
rect 8366 704 8400 719
rect 8366 685 8400 704
rect 8366 636 8400 644
rect 8366 610 8400 636
rect 8366 568 8400 569
rect 8366 535 8400 568
rect 8366 466 8400 494
rect 8366 460 8400 466
rect 8366 398 8400 419
rect 8366 385 8400 398
rect 8366 330 8400 344
rect 8366 310 8400 330
rect 8366 262 8400 269
rect 8366 235 8400 262
rect 8366 160 8400 194
rect 8582 976 8616 1008
rect 8582 974 8616 976
rect 8582 908 8616 934
rect 8582 900 8616 908
rect 8582 840 8616 860
rect 8582 826 8616 840
rect 8582 772 8616 786
rect 8582 752 8616 772
rect 8582 704 8616 712
rect 8582 678 8616 704
rect 8582 636 8616 638
rect 8582 604 8616 636
rect 8582 534 8616 564
rect 8582 530 8616 534
rect 8582 466 8616 490
rect 8582 456 8616 466
rect 8582 398 8616 416
rect 8582 382 8616 398
rect 8582 330 8616 342
rect 8582 308 8616 330
rect 8582 262 8616 268
rect 8582 234 8616 262
rect 8582 160 8616 194
rect 8798 976 8832 1008
rect 8798 974 8832 976
rect 8798 908 8832 934
rect 8798 900 8832 908
rect 8798 840 8832 860
rect 8798 826 8832 840
rect 8798 772 8832 786
rect 8798 752 8832 772
rect 8798 704 8832 712
rect 8798 678 8832 704
rect 8798 636 8832 638
rect 8798 604 8832 636
rect 8798 534 8832 564
rect 8798 530 8832 534
rect 8798 466 8832 490
rect 8798 456 8832 466
rect 8798 398 8832 416
rect 8798 382 8832 398
rect 8798 330 8832 342
rect 8798 308 8832 330
rect 8798 262 8832 268
rect 8798 234 8832 262
rect 8798 160 8832 194
rect 9014 976 9048 1008
rect 9014 974 9048 976
rect 9014 908 9048 934
rect 9014 900 9048 908
rect 9014 840 9048 860
rect 9014 826 9048 840
rect 9014 772 9048 786
rect 9014 752 9048 772
rect 9014 704 9048 712
rect 9014 678 9048 704
rect 9014 636 9048 638
rect 9014 604 9048 636
rect 9014 534 9048 564
rect 9014 530 9048 534
rect 9014 466 9048 490
rect 9014 456 9048 466
rect 9014 398 9048 416
rect 9014 382 9048 398
rect 9014 330 9048 342
rect 9014 308 9048 330
rect 9014 262 9048 268
rect 9014 234 9048 262
rect 9014 160 9048 194
rect 9230 976 9264 1008
rect 9230 974 9264 976
rect 9230 908 9264 934
rect 9230 900 9264 908
rect 9230 840 9264 860
rect 9230 826 9264 840
rect 9230 772 9264 786
rect 9230 752 9264 772
rect 9230 704 9264 712
rect 9230 678 9264 704
rect 9230 636 9264 638
rect 9230 604 9264 636
rect 9230 534 9264 564
rect 9230 530 9264 534
rect 9230 466 9264 490
rect 9230 456 9264 466
rect 9230 398 9264 416
rect 9230 382 9264 398
rect 9230 330 9264 342
rect 9230 308 9264 330
rect 9230 262 9264 268
rect 9230 234 9264 262
rect 9230 160 9264 194
rect 9446 976 9480 1008
rect 9446 974 9480 976
rect 9446 908 9480 934
rect 9446 900 9480 908
rect 9446 840 9480 860
rect 9446 826 9480 840
rect 9446 772 9480 786
rect 9446 752 9480 772
rect 9446 704 9480 712
rect 9446 678 9480 704
rect 9446 636 9480 638
rect 9446 604 9480 636
rect 9446 534 9480 564
rect 9446 530 9480 534
rect 9446 466 9480 490
rect 9446 456 9480 466
rect 9446 398 9480 416
rect 9446 382 9480 398
rect 9446 330 9480 342
rect 9446 308 9480 330
rect 9446 262 9480 268
rect 9446 234 9480 262
rect 9446 160 9480 194
rect 9662 976 9696 1008
rect 9662 974 9696 976
rect 9662 908 9696 934
rect 9662 900 9696 908
rect 9662 840 9696 860
rect 9662 826 9696 840
rect 9662 772 9696 786
rect 9662 752 9696 772
rect 9662 704 9696 712
rect 9662 678 9696 704
rect 9662 636 9696 638
rect 9662 604 9696 636
rect 9662 534 9696 564
rect 9662 530 9696 534
rect 9662 466 9696 490
rect 9662 456 9696 466
rect 9662 398 9696 416
rect 9662 382 9696 398
rect 9662 330 9696 342
rect 9662 308 9696 330
rect 9662 262 9696 268
rect 9662 234 9696 262
rect 9662 160 9696 194
rect 9878 1078 9912 1094
rect 9878 1060 9912 1078
rect 9878 1010 9912 1019
rect 9878 985 9912 1010
rect 9878 942 9912 944
rect 9878 910 9912 942
rect 9878 840 9912 869
rect 9878 835 9912 840
rect 9878 772 9912 794
rect 9878 760 9912 772
rect 9878 704 9912 719
rect 9878 685 9912 704
rect 9878 636 9912 644
rect 9878 610 9912 636
rect 9878 568 9912 569
rect 9878 535 9912 568
rect 9878 466 9912 494
rect 9878 460 9912 466
rect 9878 398 9912 419
rect 9878 385 9912 398
rect 9878 330 9912 344
rect 9878 310 9912 330
rect 9878 262 9912 269
rect 9878 235 9912 262
rect 9878 160 9912 194
rect 10094 1078 10128 1094
rect 10094 1060 10128 1078
rect 10094 1010 10128 1019
rect 10094 985 10128 1010
rect 10094 942 10128 944
rect 10094 910 10128 942
rect 10094 840 10128 869
rect 10094 835 10128 840
rect 10094 772 10128 794
rect 10094 760 10128 772
rect 10094 704 10128 719
rect 10094 685 10128 704
rect 10094 636 10128 644
rect 10094 610 10128 636
rect 10094 568 10128 569
rect 10094 535 10128 568
rect 10094 466 10128 494
rect 10094 460 10128 466
rect 10094 398 10128 419
rect 10094 385 10128 398
rect 10094 330 10128 344
rect 10094 310 10128 330
rect 10094 262 10128 269
rect 10094 235 10128 262
rect 10094 160 10128 194
rect 10310 976 10344 1008
rect 10310 974 10344 976
rect 10310 908 10344 934
rect 10310 900 10344 908
rect 10310 840 10344 860
rect 10310 826 10344 840
rect 10310 772 10344 786
rect 10310 752 10344 772
rect 10310 704 10344 712
rect 10310 678 10344 704
rect 10310 636 10344 638
rect 10310 604 10344 636
rect 10310 534 10344 564
rect 10310 530 10344 534
rect 10310 466 10344 490
rect 10310 456 10344 466
rect 10310 398 10344 416
rect 10310 382 10344 398
rect 10310 330 10344 342
rect 10310 308 10344 330
rect 10310 262 10344 268
rect 10310 234 10344 262
rect 10310 160 10344 194
rect 10526 1078 10560 1094
rect 10526 1060 10560 1078
rect 10526 1010 10560 1019
rect 10526 985 10560 1010
rect 10526 942 10560 944
rect 10526 910 10560 942
rect 10526 840 10560 869
rect 10526 835 10560 840
rect 10526 772 10560 794
rect 10526 760 10560 772
rect 10526 704 10560 719
rect 10526 685 10560 704
rect 10526 636 10560 644
rect 10526 610 10560 636
rect 10526 568 10560 569
rect 10526 535 10560 568
rect 10526 466 10560 494
rect 10526 460 10560 466
rect 10526 398 10560 419
rect 10526 385 10560 398
rect 10526 330 10560 344
rect 10526 310 10560 330
rect 10526 262 10560 269
rect 10526 235 10560 262
rect 10526 160 10560 194
rect 10742 976 10776 1008
rect 10742 974 10776 976
rect 10742 908 10776 934
rect 10742 900 10776 908
rect 10742 840 10776 860
rect 10742 826 10776 840
rect 10742 772 10776 786
rect 10742 752 10776 772
rect 10742 704 10776 712
rect 10742 678 10776 704
rect 10742 636 10776 638
rect 10742 604 10776 636
rect 10742 534 10776 564
rect 10742 530 10776 534
rect 10742 466 10776 490
rect 10742 456 10776 466
rect 10742 398 10776 416
rect 10742 382 10776 398
rect 10742 330 10776 342
rect 10742 308 10776 330
rect 10742 262 10776 268
rect 10742 234 10776 262
rect 10742 160 10776 194
rect 10958 1078 10992 1094
rect 10958 1060 10992 1078
rect 10958 1010 10992 1019
rect 10958 985 10992 1010
rect 10958 942 10992 944
rect 10958 910 10992 942
rect 10958 840 10992 869
rect 10958 835 10992 840
rect 10958 772 10992 794
rect 10958 760 10992 772
rect 10958 704 10992 719
rect 10958 685 10992 704
rect 10958 636 10992 644
rect 10958 610 10992 636
rect 10958 568 10992 569
rect 10958 535 10992 568
rect 10958 466 10992 494
rect 10958 460 10992 466
rect 10958 398 10992 419
rect 10958 385 10992 398
rect 10958 330 10992 344
rect 10958 310 10992 330
rect 10958 262 10992 269
rect 10958 235 10992 262
rect 10958 160 10992 194
rect 11174 976 11208 1008
rect 11174 974 11208 976
rect 11174 908 11208 934
rect 11174 900 11208 908
rect 11174 840 11208 860
rect 11174 826 11208 840
rect 11174 772 11208 786
rect 11174 752 11208 772
rect 11174 704 11208 712
rect 11174 678 11208 704
rect 11174 636 11208 638
rect 11174 604 11208 636
rect 11174 534 11208 564
rect 11174 530 11208 534
rect 11174 466 11208 490
rect 11174 456 11208 466
rect 11174 398 11208 416
rect 11174 382 11208 398
rect 11174 330 11208 342
rect 11174 308 11208 330
rect 11174 262 11208 268
rect 11174 234 11208 262
rect 11174 160 11208 194
rect 11390 1078 11424 1094
rect 11390 1060 11424 1078
rect 11390 1010 11424 1019
rect 11390 985 11424 1010
rect 11390 942 11424 944
rect 11390 910 11424 942
rect 11390 840 11424 869
rect 11390 835 11424 840
rect 11390 772 11424 794
rect 11390 760 11424 772
rect 11390 704 11424 719
rect 11390 685 11424 704
rect 11390 636 11424 644
rect 11390 610 11424 636
rect 11390 568 11424 569
rect 11390 535 11424 568
rect 11390 466 11424 494
rect 11390 460 11424 466
rect 11390 398 11424 419
rect 11390 385 11424 398
rect 11390 330 11424 344
rect 11390 310 11424 330
rect 11390 262 11424 269
rect 11390 235 11424 262
rect 11390 160 11424 194
rect 11606 976 11640 1008
rect 11606 974 11640 976
rect 11606 908 11640 934
rect 11606 900 11640 908
rect 11606 840 11640 860
rect 11606 826 11640 840
rect 11606 772 11640 786
rect 11606 752 11640 772
rect 11606 704 11640 712
rect 11606 678 11640 704
rect 11606 636 11640 638
rect 11606 604 11640 636
rect 11606 534 11640 564
rect 11606 530 11640 534
rect 11606 466 11640 490
rect 11606 456 11640 466
rect 11606 398 11640 416
rect 11606 382 11640 398
rect 11606 330 11640 342
rect 11606 308 11640 330
rect 11606 262 11640 268
rect 11606 234 11640 262
rect 11606 160 11640 194
rect 11823 1078 11857 1094
rect 11823 1060 11856 1078
rect 11856 1060 11857 1078
rect 11823 1010 11857 1019
rect 11823 985 11856 1010
rect 11856 985 11857 1010
rect 11823 942 11857 944
rect 11823 910 11856 942
rect 11856 910 11857 942
rect 11823 840 11856 869
rect 11856 840 11857 869
rect 11823 835 11857 840
rect 11823 772 11856 794
rect 11856 772 11857 794
rect 11823 760 11857 772
rect 11823 704 11856 719
rect 11856 704 11857 719
rect 11823 685 11857 704
rect 11823 636 11856 644
rect 11856 636 11857 644
rect 11823 610 11857 636
rect 11823 568 11856 569
rect 11856 568 11857 569
rect 11823 535 11857 568
rect 11823 466 11857 494
rect 11823 460 11856 466
rect 11856 460 11857 466
rect 11823 398 11857 419
rect 11823 385 11856 398
rect 11856 385 11857 398
rect 11823 330 11857 344
rect 11823 310 11856 330
rect 11856 310 11857 330
rect 11823 262 11857 269
rect 11823 235 11856 262
rect 11856 235 11857 262
rect 11823 160 11856 194
rect 11856 160 11857 194
rect 12038 976 12072 1008
rect 12038 974 12072 976
rect 12038 908 12072 934
rect 12038 900 12072 908
rect 12038 840 12072 860
rect 12038 826 12072 840
rect 12038 772 12072 786
rect 12038 752 12072 772
rect 12038 704 12072 712
rect 12038 678 12072 704
rect 12038 636 12072 638
rect 12038 604 12072 636
rect 12038 534 12072 564
rect 12038 530 12072 534
rect 12038 466 12072 490
rect 12038 456 12072 466
rect 12038 398 12072 416
rect 12038 382 12072 398
rect 12038 330 12072 342
rect 12038 308 12072 330
rect 12038 262 12072 268
rect 12038 234 12072 262
rect 12038 160 12072 194
rect 12254 1078 12288 1094
rect 12254 1060 12288 1078
rect 12254 1010 12288 1019
rect 12254 985 12288 1010
rect 12254 942 12288 944
rect 12254 910 12288 942
rect 12254 840 12288 869
rect 12254 835 12288 840
rect 12254 772 12288 794
rect 12254 760 12288 772
rect 12254 704 12288 719
rect 12254 685 12288 704
rect 12254 636 12288 644
rect 12254 610 12288 636
rect 12254 568 12288 569
rect 12254 535 12288 568
rect 12254 466 12288 494
rect 12254 460 12288 466
rect 12254 398 12288 419
rect 12254 385 12288 398
rect 12254 330 12288 344
rect 12254 310 12288 330
rect 12254 262 12288 269
rect 12254 235 12288 262
rect 12254 160 12288 194
rect 12470 976 12504 1008
rect 12470 974 12504 976
rect 12470 908 12504 934
rect 12470 900 12504 908
rect 12470 840 12504 860
rect 12470 826 12504 840
rect 12470 772 12504 786
rect 12470 752 12504 772
rect 12470 704 12504 712
rect 12470 678 12504 704
rect 12470 636 12504 638
rect 12470 604 12504 636
rect 12470 534 12504 564
rect 12470 530 12504 534
rect 12470 466 12504 490
rect 12470 456 12504 466
rect 12470 398 12504 416
rect 12470 382 12504 398
rect 12470 330 12504 342
rect 12470 308 12504 330
rect 12470 262 12504 268
rect 12470 234 12504 262
rect 12470 160 12504 194
rect 12686 976 12720 1008
rect 12686 974 12720 976
rect 12686 908 12720 934
rect 12686 900 12720 908
rect 12686 840 12720 860
rect 12686 826 12720 840
rect 12686 772 12720 786
rect 12686 752 12720 772
rect 12686 704 12720 712
rect 12686 678 12720 704
rect 12686 636 12720 638
rect 12686 604 12720 636
rect 12686 534 12720 564
rect 12686 530 12720 534
rect 12686 466 12720 490
rect 12686 456 12720 466
rect 12686 398 12720 416
rect 12686 382 12720 398
rect 12686 330 12720 342
rect 12686 308 12720 330
rect 12686 262 12720 268
rect 12686 234 12720 262
rect 12686 160 12720 194
rect 12902 976 12936 1008
rect 12902 974 12936 976
rect 12902 908 12936 934
rect 12902 900 12936 908
rect 12902 840 12936 860
rect 12902 826 12936 840
rect 12902 772 12936 786
rect 12902 752 12936 772
rect 12902 704 12936 712
rect 12902 678 12936 704
rect 12902 636 12936 638
rect 12902 604 12936 636
rect 12902 534 12936 564
rect 12902 530 12936 534
rect 12902 466 12936 490
rect 12902 456 12936 466
rect 12902 398 12936 416
rect 12902 382 12936 398
rect 12902 330 12936 342
rect 12902 308 12936 330
rect 12902 262 12936 268
rect 12902 234 12936 262
rect 12902 160 12936 194
rect 13118 976 13152 1008
rect 13118 974 13152 976
rect 13118 908 13152 934
rect 13118 900 13152 908
rect 13118 840 13152 860
rect 13118 826 13152 840
rect 13118 772 13152 786
rect 13118 752 13152 772
rect 13118 704 13152 712
rect 13118 678 13152 704
rect 13118 636 13152 638
rect 13118 604 13152 636
rect 13118 534 13152 564
rect 13118 530 13152 534
rect 13118 466 13152 490
rect 13118 456 13152 466
rect 13118 398 13152 416
rect 13118 382 13152 398
rect 13118 330 13152 342
rect 13118 308 13152 330
rect 13118 262 13152 268
rect 13118 234 13152 262
rect 13118 160 13152 194
rect 13334 976 13368 1008
rect 13334 974 13368 976
rect 13334 908 13368 934
rect 13334 900 13368 908
rect 13334 840 13368 860
rect 13334 826 13368 840
rect 13334 772 13368 786
rect 13334 752 13368 772
rect 13334 704 13368 712
rect 13334 678 13368 704
rect 13334 636 13368 638
rect 13334 604 13368 636
rect 13334 534 13368 564
rect 13334 530 13368 534
rect 13334 466 13368 490
rect 13334 456 13368 466
rect 13334 398 13368 416
rect 13334 382 13368 398
rect 13334 330 13368 342
rect 13334 308 13368 330
rect 13334 262 13368 268
rect 13334 234 13368 262
rect 13334 160 13368 194
rect 13550 976 13584 1008
rect 13550 974 13584 976
rect 13550 908 13584 934
rect 13550 900 13584 908
rect 13550 840 13584 860
rect 13550 826 13584 840
rect 13550 772 13584 786
rect 13550 752 13584 772
rect 13550 704 13584 712
rect 13550 678 13584 704
rect 13550 636 13584 638
rect 13550 604 13584 636
rect 13550 534 13584 564
rect 13550 530 13584 534
rect 13550 466 13584 490
rect 13550 456 13584 466
rect 13550 398 13584 416
rect 13550 382 13584 398
rect 13550 330 13584 342
rect 13550 308 13584 330
rect 13550 262 13584 268
rect 13550 234 13584 262
rect 13550 160 13584 194
rect 13766 976 13800 1008
rect 13766 974 13800 976
rect 13766 908 13800 934
rect 13766 900 13800 908
rect 13766 840 13800 860
rect 13766 826 13800 840
rect 13766 772 13800 786
rect 13766 752 13800 772
rect 13766 704 13800 712
rect 13766 678 13800 704
rect 13766 636 13800 638
rect 13766 604 13800 636
rect 13766 534 13800 564
rect 13766 530 13800 534
rect 13766 466 13800 490
rect 13766 456 13800 466
rect 13766 398 13800 416
rect 13766 382 13800 398
rect 13766 330 13800 342
rect 13766 308 13800 330
rect 13766 262 13800 268
rect 13766 234 13800 262
rect 13766 160 13800 194
rect 13982 976 14016 1008
rect 13982 974 14016 976
rect 13982 908 14016 934
rect 13982 900 14016 908
rect 13982 840 14016 860
rect 13982 826 14016 840
rect 13982 772 14016 786
rect 13982 752 14016 772
rect 13982 704 14016 712
rect 13982 678 14016 704
rect 13982 636 14016 638
rect 13982 604 14016 636
rect 13982 534 14016 564
rect 13982 530 14016 534
rect 13982 466 14016 490
rect 13982 456 14016 466
rect 13982 398 14016 416
rect 13982 382 14016 398
rect 13982 330 14016 342
rect 13982 308 14016 330
rect 13982 262 14016 268
rect 13982 234 14016 262
rect 13982 160 14016 194
rect 14198 976 14232 1008
rect 14198 974 14232 976
rect 14198 908 14232 934
rect 14198 900 14232 908
rect 14198 840 14232 860
rect 14198 826 14232 840
rect 14198 772 14232 786
rect 14198 752 14232 772
rect 14198 704 14232 712
rect 14198 678 14232 704
rect 14198 636 14232 638
rect 14198 604 14232 636
rect 14198 534 14232 564
rect 14198 530 14232 534
rect 14198 466 14232 490
rect 14198 456 14232 466
rect 14198 398 14232 416
rect 14198 382 14232 398
rect 14198 330 14232 342
rect 14198 308 14232 330
rect 14198 262 14232 268
rect 14198 234 14232 262
rect 14198 160 14232 194
rect 14414 976 14448 1008
rect 14414 974 14448 976
rect 14414 908 14448 934
rect 14414 900 14448 908
rect 14414 840 14448 860
rect 14414 826 14448 840
rect 14414 772 14448 786
rect 14414 752 14448 772
rect 14414 704 14448 712
rect 14414 678 14448 704
rect 14414 636 14448 638
rect 14414 604 14448 636
rect 14414 534 14448 564
rect 14414 530 14448 534
rect 14414 466 14448 490
rect 14414 456 14448 466
rect 14414 398 14448 416
rect 14414 382 14448 398
rect 14414 330 14448 342
rect 14414 308 14448 330
rect 14414 262 14448 268
rect 14414 234 14448 262
rect 14414 160 14448 194
rect 14630 976 14664 1008
rect 14630 974 14664 976
rect 14630 908 14664 934
rect 14630 900 14664 908
rect 14630 840 14664 860
rect 14630 826 14664 840
rect 14630 772 14664 786
rect 14630 752 14664 772
rect 14630 704 14664 712
rect 14630 678 14664 704
rect 14630 636 14664 638
rect 14630 604 14664 636
rect 14630 534 14664 564
rect 14630 530 14664 534
rect 14630 466 14664 490
rect 14630 456 14664 466
rect 14630 398 14664 416
rect 14630 382 14664 398
rect 14630 330 14664 342
rect 14630 308 14664 330
rect 14630 262 14664 268
rect 14630 234 14664 262
rect 14630 160 14664 194
rect 14846 976 14880 1008
rect 14846 974 14880 976
rect 14846 908 14880 934
rect 14846 900 14880 908
rect 14846 840 14880 860
rect 14846 826 14880 840
rect 14846 772 14880 786
rect 14846 752 14880 772
rect 14846 704 14880 712
rect 14846 678 14880 704
rect 14846 636 14880 638
rect 14846 604 14880 636
rect 14846 534 14880 564
rect 14846 530 14880 534
rect 14846 466 14880 490
rect 14846 456 14880 466
rect 14846 398 14880 416
rect 14846 382 14880 398
rect 14846 330 14880 342
rect 14846 308 14880 330
rect 14846 262 14880 268
rect 14846 234 14880 262
rect 14846 160 14880 194
rect 15062 976 15096 1008
rect 15062 974 15096 976
rect 15062 908 15096 934
rect 15062 900 15096 908
rect 15062 840 15096 860
rect 15062 826 15096 840
rect 15062 772 15096 786
rect 15062 752 15096 772
rect 15062 704 15096 712
rect 15062 678 15096 704
rect 15062 636 15096 638
rect 15062 604 15096 636
rect 15062 534 15096 564
rect 15172 1070 15206 1093
rect 15172 1059 15206 1070
rect 15172 1002 15206 1012
rect 15172 978 15206 1002
rect 15172 900 15206 931
rect 15172 897 15206 900
rect 15172 832 15206 850
rect 15172 816 15206 832
rect 15172 764 15206 768
rect 15172 734 15206 764
rect 15172 662 15206 686
rect 15172 652 15206 662
rect 15172 594 15206 604
rect 15172 570 15206 594
rect 15428 1070 15462 1093
rect 15428 1059 15462 1070
rect 15428 1002 15462 1012
rect 15428 978 15462 1002
rect 15428 900 15462 931
rect 15428 897 15462 900
rect 15428 832 15462 850
rect 15428 816 15462 832
rect 15428 764 15462 768
rect 15428 734 15462 764
rect 15428 662 15462 686
rect 15428 652 15462 662
rect 15428 594 15462 604
rect 15428 570 15462 594
rect 15538 1078 15572 1094
rect 15538 1060 15572 1078
rect 15538 1010 15572 1019
rect 15538 985 15572 1010
rect 15538 942 15572 944
rect 15538 910 15572 942
rect 15538 840 15572 869
rect 15538 835 15572 840
rect 15538 772 15572 794
rect 15538 760 15572 772
rect 15538 704 15572 719
rect 15538 685 15572 704
rect 15538 636 15572 644
rect 15538 610 15572 636
rect 15538 568 15572 569
rect 15062 530 15096 534
rect 15062 466 15096 490
rect 15062 456 15096 466
rect 15062 398 15096 416
rect 15062 382 15096 398
rect 15062 330 15096 342
rect 15062 308 15096 330
rect 15062 262 15096 268
rect 15062 234 15096 262
rect 15062 160 15096 194
rect 15538 535 15572 568
rect 15538 466 15572 494
rect 15538 460 15572 466
rect 15538 398 15572 419
rect 15538 385 15572 398
rect 15538 330 15572 344
rect 15538 310 15572 330
rect 15538 262 15572 269
rect 15538 235 15572 262
rect 15538 160 15572 194
rect 15754 1078 15788 1094
rect 15754 1060 15788 1078
rect 15754 1010 15788 1019
rect 15754 985 15788 1010
rect 15754 942 15788 944
rect 15754 910 15788 942
rect 15754 840 15788 869
rect 15754 835 15788 840
rect 15754 772 15788 794
rect 15754 760 15788 772
rect 15754 704 15788 719
rect 15754 685 15788 704
rect 15754 636 15788 644
rect 15754 610 15788 636
rect 15754 568 15788 569
rect 15754 535 15788 568
rect 15754 466 15788 494
rect 15754 460 15788 466
rect 15754 398 15788 419
rect 15754 385 15788 398
rect 15754 330 15788 344
rect 15754 310 15788 330
rect 15754 262 15788 269
rect 15754 235 15788 262
rect 15754 160 15788 194
rect 15970 1078 16004 1094
rect 15970 1060 16004 1078
rect 15970 1010 16004 1019
rect 15970 985 16004 1010
rect 15970 942 16004 944
rect 15970 910 16004 942
rect 15970 840 16004 869
rect 15970 835 16004 840
rect 15970 772 16004 794
rect 15970 760 16004 772
rect 15970 704 16004 719
rect 15970 685 16004 704
rect 15970 636 16004 644
rect 15970 610 16004 636
rect 15970 568 16004 569
rect 15970 535 16004 568
rect 15970 466 16004 494
rect 15970 460 16004 466
rect 15970 398 16004 419
rect 15970 385 16004 398
rect 15970 330 16004 344
rect 15970 310 16004 330
rect 15970 262 16004 269
rect 15970 235 16004 262
rect 15970 160 16004 194
rect 1622 48 1631 82
rect 1631 48 1656 82
rect 1696 48 1705 82
rect 1705 48 1730 82
rect 1770 48 1779 82
rect 1779 48 1804 82
rect 1844 48 1853 82
rect 1853 48 1878 82
rect 1918 48 1927 82
rect 1927 48 1952 82
rect 1992 48 2001 82
rect 2001 48 2026 82
rect 2066 48 2074 82
rect 2074 48 2100 82
rect 2140 48 2147 82
rect 2147 48 2174 82
rect 2214 48 2220 82
rect 2220 48 2248 82
rect 2287 48 2293 82
rect 2293 48 2321 82
rect 2991 48 3003 82
rect 3003 48 3025 82
rect 3065 48 3072 82
rect 3072 48 3099 82
rect 3139 48 3141 82
rect 3141 48 3173 82
rect 3213 48 3244 82
rect 3244 48 3247 82
rect 3288 48 3313 82
rect 3313 48 3322 82
rect 3363 48 3382 82
rect 3382 48 3397 82
rect 3946 40 3958 74
rect 3958 40 3980 74
rect 4020 40 4028 74
rect 4028 40 4054 74
rect 4094 40 4098 74
rect 4098 40 4128 74
rect 4168 40 4202 74
rect 4242 40 4272 74
rect 4272 40 4276 74
rect 4316 40 4342 74
rect 4342 40 4350 74
rect 4390 40 4412 74
rect 4412 40 4424 74
rect 4464 40 4482 74
rect 4482 40 4498 74
rect 4538 40 4552 74
rect 4552 40 4572 74
rect 4612 40 4621 74
rect 4621 40 4646 74
rect 4685 40 4690 74
rect 4690 40 4719 74
rect 4758 40 4759 74
rect 4759 40 4792 74
rect 4831 40 4863 74
rect 4863 40 4865 74
rect 4904 40 4932 74
rect 4932 40 4938 74
rect 4977 40 5001 74
rect 5001 40 5011 74
rect 5050 40 5070 74
rect 5070 40 5084 74
rect 5123 40 5139 74
rect 5139 40 5157 74
rect 5196 40 5208 74
rect 5208 40 5230 74
rect 5269 40 5277 74
rect 5277 40 5303 74
rect 5342 40 5346 74
rect 5346 40 5376 74
rect 5415 40 5449 74
rect 5488 40 5518 74
rect 5518 40 5522 74
rect 5561 40 5587 74
rect 5587 40 5595 74
rect 5634 40 5656 74
rect 5656 40 5668 74
rect 5889 44 5923 78
rect 5962 74 5996 78
rect 6035 74 6069 78
rect 6108 74 6142 78
rect 5962 44 5974 74
rect 5974 44 5996 74
rect 6035 44 6043 74
rect 6043 44 6069 74
rect 6108 44 6112 74
rect 6112 44 6142 74
rect 6181 44 6215 78
rect 6254 74 6288 78
rect 6327 74 6361 78
rect 6400 74 6434 78
rect 6473 74 6507 78
rect 6546 74 6580 78
rect 6619 74 6653 78
rect 6692 74 6726 78
rect 6765 74 6799 78
rect 6838 74 6872 78
rect 6911 74 6945 78
rect 6984 74 7018 78
rect 7057 74 7091 78
rect 7130 74 7164 78
rect 7203 74 7237 78
rect 7276 74 7310 78
rect 7349 74 7383 78
rect 7422 74 7456 78
rect 7495 74 7529 78
rect 7568 74 7602 78
rect 7641 74 7675 78
rect 7714 74 7748 78
rect 7787 74 7821 78
rect 7860 74 7894 78
rect 7933 74 7967 78
rect 8006 74 8040 78
rect 8079 74 8113 78
rect 8152 74 8186 78
rect 8225 74 8259 78
rect 8298 74 8332 78
rect 8371 74 8405 78
rect 8444 74 8478 78
rect 8517 74 8551 78
rect 8590 74 8624 78
rect 8663 74 8697 78
rect 8736 74 8770 78
rect 8809 74 8843 78
rect 8882 74 8916 78
rect 8955 74 8989 78
rect 9028 74 9062 78
rect 9101 74 9135 78
rect 6254 44 6284 74
rect 6284 44 6288 74
rect 6327 44 6352 74
rect 6352 44 6361 74
rect 6400 44 6420 74
rect 6420 44 6434 74
rect 6473 44 6488 74
rect 6488 44 6507 74
rect 6546 44 6556 74
rect 6556 44 6580 74
rect 6619 44 6624 74
rect 6624 44 6653 74
rect 6692 44 6726 74
rect 6765 44 6794 74
rect 6794 44 6799 74
rect 6838 44 6862 74
rect 6862 44 6872 74
rect 6911 44 6930 74
rect 6930 44 6945 74
rect 6984 44 6998 74
rect 6998 44 7018 74
rect 7057 44 7066 74
rect 7066 44 7091 74
rect 7130 44 7134 74
rect 7134 44 7164 74
rect 7203 44 7236 74
rect 7236 44 7237 74
rect 7276 44 7304 74
rect 7304 44 7310 74
rect 7349 44 7372 74
rect 7372 44 7383 74
rect 7422 44 7440 74
rect 7440 44 7456 74
rect 7495 44 7508 74
rect 7508 44 7529 74
rect 7568 44 7576 74
rect 7576 44 7602 74
rect 7641 44 7644 74
rect 7644 44 7675 74
rect 7714 44 7746 74
rect 7746 44 7748 74
rect 7787 44 7814 74
rect 7814 44 7821 74
rect 7860 44 7882 74
rect 7882 44 7894 74
rect 7933 44 7950 74
rect 7950 44 7967 74
rect 8006 44 8018 74
rect 8018 44 8040 74
rect 8079 44 8086 74
rect 8086 44 8113 74
rect 8152 44 8154 74
rect 8154 44 8186 74
rect 8225 44 8256 74
rect 8256 44 8259 74
rect 8298 44 8324 74
rect 8324 44 8332 74
rect 8371 44 8392 74
rect 8392 44 8405 74
rect 8444 44 8460 74
rect 8460 44 8478 74
rect 8517 44 8528 74
rect 8528 44 8551 74
rect 8590 44 8596 74
rect 8596 44 8624 74
rect 8663 44 8664 74
rect 8664 44 8697 74
rect 8736 44 8766 74
rect 8766 44 8770 74
rect 8809 44 8834 74
rect 8834 44 8843 74
rect 8882 44 8902 74
rect 8902 44 8916 74
rect 8955 44 8970 74
rect 8970 44 8989 74
rect 9028 44 9038 74
rect 9038 44 9062 74
rect 9101 44 9106 74
rect 9106 44 9135 74
rect 9174 44 9208 78
rect 9247 74 9281 78
rect 9320 74 9354 78
rect 9393 74 9427 78
rect 9466 74 9500 78
rect 9539 74 9573 78
rect 9612 74 9646 78
rect 9685 74 9719 78
rect 9758 74 9792 78
rect 9831 74 9865 78
rect 9903 74 9937 78
rect 9975 74 10009 78
rect 10047 74 10081 78
rect 10119 74 10153 78
rect 10191 74 10225 78
rect 10263 74 10297 78
rect 10335 74 10369 78
rect 10407 74 10441 78
rect 10479 74 10513 78
rect 10551 74 10585 78
rect 10623 74 10657 78
rect 10695 74 10729 78
rect 10767 74 10801 78
rect 10839 74 10873 78
rect 10911 74 10945 78
rect 10983 74 11017 78
rect 11055 74 11089 78
rect 11127 74 11161 78
rect 11199 74 11233 78
rect 11271 74 11305 78
rect 11343 74 11377 78
rect 11415 74 11449 78
rect 11487 74 11521 78
rect 11559 74 11593 78
rect 11631 74 11665 78
rect 11703 74 11737 78
rect 11775 74 11809 78
rect 11847 74 11881 78
rect 11919 74 11953 78
rect 11991 74 12025 78
rect 12063 74 12097 78
rect 12135 74 12169 78
rect 12207 74 12241 78
rect 12279 74 12313 78
rect 12351 74 12385 78
rect 12423 74 12457 78
rect 12495 74 12529 78
rect 12567 74 12601 78
rect 12639 74 12673 78
rect 12711 74 12745 78
rect 12783 74 12817 78
rect 12855 74 12889 78
rect 12927 74 12961 78
rect 12999 74 13033 78
rect 13071 74 13105 78
rect 13143 74 13177 78
rect 13215 74 13249 78
rect 13287 74 13321 78
rect 13359 74 13393 78
rect 13431 74 13465 78
rect 13503 74 13537 78
rect 13575 74 13609 78
rect 13647 74 13681 78
rect 13719 74 13753 78
rect 13791 74 13825 78
rect 13863 74 13897 78
rect 13935 74 13969 78
rect 14007 74 14041 78
rect 14079 74 14113 78
rect 14151 74 14185 78
rect 14223 74 14257 78
rect 14295 74 14329 78
rect 14367 74 14401 78
rect 14439 74 14473 78
rect 14511 74 14545 78
rect 14583 74 14617 78
rect 14655 74 14689 78
rect 14727 74 14761 78
rect 14799 74 14833 78
rect 14871 74 14905 78
rect 14943 74 14977 78
rect 15015 74 15049 78
rect 15087 74 15121 78
rect 15159 74 15193 78
rect 15231 74 15265 78
rect 15303 74 15337 78
rect 15375 74 15409 78
rect 15447 74 15481 78
rect 15519 74 15553 78
rect 15591 74 15625 78
rect 15663 74 15697 78
rect 15735 74 15769 78
rect 15807 74 15841 78
rect 15879 74 15913 78
rect 15951 74 15985 78
rect 9247 44 9276 74
rect 9276 44 9281 74
rect 9320 44 9344 74
rect 9344 44 9354 74
rect 9393 44 9412 74
rect 9412 44 9427 74
rect 9466 44 9480 74
rect 9480 44 9500 74
rect 9539 44 9548 74
rect 9548 44 9573 74
rect 9612 44 9616 74
rect 9616 44 9646 74
rect 9685 44 9718 74
rect 9718 44 9719 74
rect 9758 44 9786 74
rect 9786 44 9792 74
rect 9831 44 9854 74
rect 9854 44 9865 74
rect 9903 44 9922 74
rect 9922 44 9937 74
rect 9975 44 9990 74
rect 9990 44 10009 74
rect 10047 44 10058 74
rect 10058 44 10081 74
rect 10119 44 10126 74
rect 10126 44 10153 74
rect 10191 44 10194 74
rect 10194 44 10225 74
rect 10263 44 10296 74
rect 10296 44 10297 74
rect 10335 44 10364 74
rect 10364 44 10369 74
rect 10407 44 10432 74
rect 10432 44 10441 74
rect 10479 44 10500 74
rect 10500 44 10513 74
rect 10551 44 10568 74
rect 10568 44 10585 74
rect 10623 44 10636 74
rect 10636 44 10657 74
rect 10695 44 10704 74
rect 10704 44 10729 74
rect 10767 44 10772 74
rect 10772 44 10801 74
rect 10839 44 10840 74
rect 10840 44 10873 74
rect 10911 44 10942 74
rect 10942 44 10945 74
rect 10983 44 11010 74
rect 11010 44 11017 74
rect 11055 44 11078 74
rect 11078 44 11089 74
rect 11127 44 11146 74
rect 11146 44 11161 74
rect 11199 44 11214 74
rect 11214 44 11233 74
rect 11271 44 11282 74
rect 11282 44 11305 74
rect 11343 44 11350 74
rect 11350 44 11377 74
rect 11415 44 11418 74
rect 11418 44 11449 74
rect 11487 44 11520 74
rect 11520 44 11521 74
rect 11559 44 11588 74
rect 11588 44 11593 74
rect 11631 44 11656 74
rect 11656 44 11665 74
rect 11703 44 11724 74
rect 11724 44 11737 74
rect 11775 44 11792 74
rect 11792 44 11809 74
rect 11847 44 11860 74
rect 11860 44 11881 74
rect 11919 44 11928 74
rect 11928 44 11953 74
rect 11991 44 11996 74
rect 11996 44 12025 74
rect 12063 44 12064 74
rect 12064 44 12097 74
rect 12135 44 12166 74
rect 12166 44 12169 74
rect 12207 44 12234 74
rect 12234 44 12241 74
rect 12279 44 12302 74
rect 12302 44 12313 74
rect 12351 44 12370 74
rect 12370 44 12385 74
rect 12423 44 12438 74
rect 12438 44 12457 74
rect 12495 44 12506 74
rect 12506 44 12529 74
rect 12567 44 12574 74
rect 12574 44 12601 74
rect 12639 44 12642 74
rect 12642 44 12673 74
rect 12711 44 12744 74
rect 12744 44 12745 74
rect 12783 44 12812 74
rect 12812 44 12817 74
rect 12855 44 12880 74
rect 12880 44 12889 74
rect 12927 44 12948 74
rect 12948 44 12961 74
rect 12999 44 13016 74
rect 13016 44 13033 74
rect 13071 44 13084 74
rect 13084 44 13105 74
rect 13143 44 13152 74
rect 13152 44 13177 74
rect 13215 44 13220 74
rect 13220 44 13249 74
rect 13287 44 13288 74
rect 13288 44 13321 74
rect 13359 44 13390 74
rect 13390 44 13393 74
rect 13431 44 13458 74
rect 13458 44 13465 74
rect 13503 44 13526 74
rect 13526 44 13537 74
rect 13575 44 13594 74
rect 13594 44 13609 74
rect 13647 44 13662 74
rect 13662 44 13681 74
rect 13719 44 13730 74
rect 13730 44 13753 74
rect 13791 44 13798 74
rect 13798 44 13825 74
rect 13863 44 13866 74
rect 13866 44 13897 74
rect 13935 44 13968 74
rect 13968 44 13969 74
rect 14007 44 14036 74
rect 14036 44 14041 74
rect 14079 44 14104 74
rect 14104 44 14113 74
rect 14151 44 14172 74
rect 14172 44 14185 74
rect 14223 44 14240 74
rect 14240 44 14257 74
rect 14295 44 14308 74
rect 14308 44 14329 74
rect 14367 44 14376 74
rect 14376 44 14401 74
rect 14439 44 14444 74
rect 14444 44 14473 74
rect 14511 44 14512 74
rect 14512 44 14545 74
rect 14583 44 14614 74
rect 14614 44 14617 74
rect 14655 44 14682 74
rect 14682 44 14689 74
rect 14727 44 14750 74
rect 14750 44 14761 74
rect 14799 44 14818 74
rect 14818 44 14833 74
rect 14871 44 14886 74
rect 14886 44 14905 74
rect 14943 44 14954 74
rect 14954 44 14977 74
rect 15015 44 15022 74
rect 15022 44 15049 74
rect 15087 44 15090 74
rect 15090 44 15121 74
rect 15159 44 15192 74
rect 15192 44 15193 74
rect 15231 44 15260 74
rect 15260 44 15265 74
rect 15303 44 15328 74
rect 15328 44 15337 74
rect 15375 44 15396 74
rect 15396 44 15409 74
rect 15447 44 15464 74
rect 15464 44 15481 74
rect 15519 44 15532 74
rect 15532 44 15553 74
rect 15591 44 15600 74
rect 15600 44 15625 74
rect 15663 44 15668 74
rect 15668 44 15697 74
rect 15735 44 15736 74
rect 15736 44 15769 74
rect 15807 44 15838 74
rect 15838 44 15841 74
rect 15879 44 15906 74
rect 15906 44 15913 74
rect 15951 44 15974 74
rect 15974 44 15985 74
<< metal1 >>
rect 9497 3297 11735 3298
rect 204 3272 9058 3278
rect 204 3238 292 3272
rect 326 3238 374 3272
rect 408 3238 456 3272
rect 490 3238 538 3272
rect 572 3238 648 3272
rect 682 3238 720 3272
rect 754 3238 792 3272
rect 826 3238 864 3272
rect 898 3238 936 3272
rect 970 3238 1008 3272
rect 1042 3238 1080 3272
rect 1114 3238 1152 3272
rect 1186 3238 1224 3272
rect 1258 3238 1296 3272
rect 1330 3238 1368 3272
rect 1402 3238 1440 3272
rect 1474 3238 1512 3272
rect 1546 3238 1584 3272
rect 1618 3238 1656 3272
rect 1690 3238 1728 3272
rect 1762 3238 1800 3272
rect 1834 3238 1872 3272
rect 1906 3238 1944 3272
rect 1978 3238 2016 3272
rect 2050 3238 2088 3272
rect 2122 3238 2160 3272
rect 2194 3238 2232 3272
rect 2266 3238 2304 3272
rect 2338 3238 2376 3272
rect 2410 3238 2448 3272
rect 2482 3238 2520 3272
rect 2554 3238 2592 3272
rect 2626 3238 2664 3272
rect 2698 3238 2736 3272
rect 2770 3238 2808 3272
rect 2842 3238 2880 3272
rect 2914 3238 2952 3272
rect 2986 3238 3024 3272
rect 3058 3238 3096 3272
rect 3130 3238 3168 3272
rect 3202 3238 3240 3272
rect 3274 3238 3312 3272
rect 3346 3238 3384 3272
rect 3418 3238 3456 3272
rect 3490 3238 3528 3272
rect 3562 3238 3600 3272
rect 3634 3238 3672 3272
rect 3706 3238 3744 3272
rect 3778 3238 3816 3272
rect 3850 3238 3888 3272
rect 3922 3238 3960 3272
rect 3994 3238 4032 3272
rect 4066 3238 4104 3272
rect 4138 3238 4176 3272
rect 4210 3238 4248 3272
rect 4282 3238 4320 3272
rect 4354 3238 4392 3272
rect 4426 3238 4464 3272
rect 4498 3238 4536 3272
rect 4570 3238 4608 3272
rect 4642 3238 4680 3272
rect 4714 3238 4752 3272
rect 4786 3238 4824 3272
rect 4858 3238 5170 3272
rect 5204 3238 5245 3272
rect 5279 3238 5320 3272
rect 5354 3238 5395 3272
rect 5429 3238 5470 3272
rect 5504 3238 5545 3272
rect 5579 3238 5619 3272
rect 5653 3238 5693 3272
rect 5727 3238 5767 3272
rect 5801 3238 5841 3272
rect 5875 3238 5915 3272
rect 5949 3238 5989 3272
rect 6023 3238 6063 3272
rect 6097 3238 6137 3272
rect 6171 3238 6211 3272
rect 6245 3238 6285 3272
rect 6319 3238 6359 3272
rect 6393 3238 6433 3272
rect 6467 3238 6507 3272
rect 6541 3238 6581 3272
rect 6615 3238 6655 3272
rect 6689 3238 6729 3272
rect 6763 3238 6803 3272
rect 6837 3238 7077 3272
rect 7111 3238 7155 3272
rect 7189 3238 7233 3272
rect 7267 3238 7311 3272
rect 7345 3238 7390 3272
rect 7424 3238 7469 3272
rect 7503 3238 7548 3272
rect 7582 3238 7627 3272
rect 7661 3238 7737 3272
rect 7771 3238 7812 3272
rect 7846 3238 7887 3272
rect 7921 3238 7962 3272
rect 7996 3238 8037 3272
rect 8071 3238 8112 3272
rect 8146 3238 8187 3272
rect 8221 3238 8262 3272
rect 8296 3238 8338 3272
rect 8372 3238 8414 3272
rect 8448 3238 8490 3272
rect 8524 3238 8566 3272
rect 8600 3238 8642 3272
rect 8676 3238 8718 3272
rect 8752 3238 8794 3272
rect 8828 3238 8870 3272
rect 8904 3238 8946 3272
rect 8980 3238 9058 3272
rect 204 3232 9058 3238
rect 204 3200 7039 3232
rect 204 3166 210 3200
rect 244 3198 6877 3200
rect 244 3166 4896 3198
rect 204 3164 4896 3166
rect 4930 3164 5098 3198
rect 5132 3166 6877 3198
rect 6911 3166 6999 3200
rect 7033 3166 7039 3200
tri 7039 3198 7073 3232 nw
tri 8978 3198 9012 3232 ne
rect 9012 3198 9058 3232
rect 5132 3164 7039 3166
rect 204 3127 7039 3164
rect 204 3126 6999 3127
rect 204 3124 6877 3126
rect 204 3113 4896 3124
rect -189 3030 -183 3082
rect -131 3030 -119 3082
rect -67 3030 -61 3082
tri -150 3026 -146 3030 ne
rect -146 3026 -61 3030
tri -146 2992 -112 3026 ne
rect -112 2992 -61 3026
tri -112 2987 -107 2992 ne
rect -107 2764 -61 2992
rect 204 3079 210 3113
rect 244 3090 4896 3113
rect 4930 3090 5098 3124
rect 5132 3092 6877 3124
rect 6911 3093 6999 3126
rect 7033 3093 7039 3127
rect 6911 3092 7039 3093
rect 5132 3090 7039 3092
rect 244 3088 7039 3090
rect 244 3079 251 3088
rect 204 3055 251 3079
tri 251 3055 284 3088 nw
tri 4844 3055 4877 3088 ne
rect 4877 3055 5139 3088
tri 5139 3055 5172 3088 nw
tri 6825 3055 6858 3088 ne
rect 6858 3055 7039 3088
rect 9012 3164 9018 3198
rect 9052 3164 9058 3198
rect 9012 3124 9058 3164
rect 9012 3090 9018 3124
rect 9052 3090 9058 3124
rect 204 3026 250 3055
tri 250 3054 251 3055 nw
rect 204 2992 210 3026
rect 244 2992 250 3026
rect 204 2939 250 2992
rect 204 2905 210 2939
rect 244 2905 250 2939
rect 204 2858 250 2905
rect 193 2812 250 2858
rect 424 3049 4716 3055
tri 4877 3054 4878 3055 ne
rect 4878 3054 5138 3055
tri 5138 3054 5139 3055 nw
tri 4878 3052 4880 3054 ne
rect 4880 3052 5138 3054
tri 4880 3050 4882 3052 ne
rect 4882 3050 5138 3052
rect 424 3015 505 3049
rect 539 3015 577 3049
rect 611 3015 649 3049
rect 683 3015 721 3049
rect 755 3015 794 3049
rect 828 3015 867 3049
rect 901 3015 940 3049
rect 974 3015 1013 3049
rect 1047 3015 1086 3049
rect 1120 3015 1159 3049
rect 1193 3015 1232 3049
rect 1266 3015 1305 3049
rect 1339 3015 1378 3049
rect 1412 3015 1451 3049
rect 1485 3015 1524 3049
rect 1558 3015 1597 3049
rect 1631 3015 1670 3049
rect 1704 3015 1743 3049
rect 1777 3015 1816 3049
rect 1850 3015 1889 3049
rect 1923 3015 1962 3049
rect 1996 3015 2035 3049
rect 2069 3015 2108 3049
rect 2142 3015 2181 3049
rect 2215 3015 2254 3049
rect 2288 3015 2327 3049
rect 2361 3015 2400 3049
rect 2434 3015 2473 3049
rect 2507 3015 2546 3049
rect 2580 3015 2619 3049
rect 2653 3015 2692 3049
rect 2726 3015 2765 3049
rect 2799 3015 2838 3049
rect 2872 3015 2911 3049
rect 2945 3015 2984 3049
rect 3018 3015 3057 3049
rect 3091 3015 3130 3049
rect 3164 3015 3203 3049
rect 3237 3015 3276 3049
rect 3310 3015 3349 3049
rect 3383 3015 3422 3049
rect 3456 3015 3495 3049
rect 3529 3015 3568 3049
rect 3602 3015 3678 3049
rect 3712 3015 3754 3049
rect 3788 3015 3831 3049
rect 3865 3015 3908 3049
rect 3942 3015 3985 3049
rect 4019 3015 4062 3049
rect 4096 3015 4139 3049
rect 4173 3015 4216 3049
rect 4250 3015 4293 3049
rect 4327 3015 4370 3049
rect 4404 3015 4447 3049
rect 4481 3015 4524 3049
rect 4558 3015 4601 3049
rect 4635 3015 4716 3049
tri 4882 3042 4890 3050 ne
rect 424 3009 4716 3015
rect 424 2982 483 3009
tri 483 2982 510 3009 nw
tri 4630 2982 4657 3009 ne
rect 4657 2982 4716 3009
rect 424 2981 482 2982
tri 482 2981 483 2982 nw
tri 4657 2981 4658 2982 ne
rect 4658 2981 4716 2982
rect 424 2978 479 2981
tri 479 2978 482 2981 nw
tri 4658 2978 4661 2981 ne
rect 4661 2978 4716 2981
rect 424 2977 478 2978
tri 478 2977 479 2978 nw
tri 4661 2977 4662 2978 ne
rect 4662 2977 4716 2978
rect 424 2943 433 2977
rect 467 2976 477 2977
tri 477 2976 478 2977 nw
tri 4662 2976 4663 2977 ne
rect 4663 2976 4716 2977
rect 467 2943 476 2976
tri 476 2975 477 2976 nw
tri 4663 2975 4664 2976 ne
rect 4664 2975 4716 2976
rect 424 2902 476 2943
rect 424 2868 433 2902
rect 467 2868 476 2902
rect 827 2891 833 2943
rect 885 2891 897 2943
rect 949 2891 955 2943
rect 4664 2941 4673 2975
rect 4707 2941 4716 2975
tri 836 2879 848 2891 ne
rect 848 2879 938 2891
tri 938 2879 950 2891 nw
rect 424 2827 476 2868
rect 193 2780 239 2812
rect -107 2730 -101 2764
rect -67 2730 -61 2764
rect -107 2684 -61 2730
rect -107 2650 -101 2684
rect -67 2650 -61 2684
rect -107 2604 -61 2650
rect -107 2570 -101 2604
rect -67 2570 -61 2604
rect -107 2523 -61 2570
rect -107 2489 -101 2523
rect -67 2489 -61 2523
rect -107 2442 -61 2489
rect -107 2408 -101 2442
rect -67 2408 -61 2442
rect -107 2361 -61 2408
rect -107 2327 -101 2361
rect -67 2327 -61 2361
rect -107 2280 -61 2327
rect -107 2246 -101 2280
rect -67 2246 -61 2280
rect -107 2234 -61 2246
rect 49 2764 158 2776
rect 49 2730 55 2764
rect 89 2730 158 2764
rect 49 2684 158 2730
rect 49 2650 55 2684
rect 89 2650 158 2684
rect 49 2604 158 2650
rect 49 2570 55 2604
rect 89 2570 158 2604
rect 49 2523 158 2570
rect 49 2489 55 2523
rect 89 2489 158 2523
rect 49 2442 158 2489
rect 49 2408 55 2442
rect 89 2408 158 2442
rect 49 2361 158 2408
rect 49 2327 55 2361
rect 89 2327 158 2361
rect 49 2280 158 2327
rect 49 2246 55 2280
rect 89 2246 158 2280
rect 49 2234 158 2246
tri 95 2221 108 2234 ne
rect 108 2221 158 2234
tri 108 2214 115 2221 ne
rect -71 2190 65 2196
rect -71 2156 -59 2190
rect -25 2156 13 2190
rect 47 2156 65 2190
rect -71 2144 65 2156
tri 97 1638 115 1656 se
rect 115 1638 158 2221
rect 193 2746 199 2780
rect 233 2746 239 2780
rect 193 2705 239 2746
rect 193 2671 199 2705
rect 233 2671 239 2705
rect 193 2630 239 2671
rect 193 2596 199 2630
rect 233 2596 239 2630
rect 193 2555 239 2596
rect 193 2521 199 2555
rect 233 2521 239 2555
rect 193 2480 239 2521
rect 193 2446 199 2480
rect 233 2446 239 2480
rect 193 2405 239 2446
rect 193 2371 199 2405
rect 233 2371 239 2405
rect 193 2330 239 2371
rect 193 2296 199 2330
rect 233 2296 239 2330
rect 193 2255 239 2296
rect 193 2221 199 2255
rect 233 2221 239 2255
rect 193 2180 239 2221
rect 193 2146 199 2180
rect 233 2146 239 2180
rect 193 2106 239 2146
rect 193 2072 199 2106
rect 233 2072 239 2106
rect 193 2032 239 2072
rect 193 1998 199 2032
rect 233 1998 239 2032
rect 193 1958 239 1998
rect 193 1924 199 1958
rect 233 1924 239 1958
rect 193 1890 239 1924
rect 424 2793 433 2827
rect 467 2793 476 2827
rect 424 2752 476 2793
rect 424 2718 433 2752
rect 467 2718 476 2752
rect 424 2677 476 2718
rect 424 2643 433 2677
rect 467 2643 476 2677
rect 424 2602 476 2643
rect 424 2568 433 2602
rect 467 2568 476 2602
rect 424 2528 476 2568
rect 424 2494 433 2528
rect 467 2494 476 2528
rect 424 2454 476 2494
rect 424 2420 433 2454
rect 467 2420 476 2454
rect 424 2380 476 2420
rect 424 2346 433 2380
rect 467 2346 476 2380
rect 424 2306 476 2346
rect 424 2272 433 2306
rect 467 2272 476 2306
rect 424 2232 476 2272
rect 424 2231 433 2232
rect 467 2231 476 2232
rect 424 2166 476 2179
rect 424 2084 476 2114
rect 711 2867 763 2879
tri 848 2867 860 2879 ne
rect 860 2867 926 2879
tri 926 2867 938 2879 nw
rect 1023 2867 1075 2879
rect 711 2833 720 2867
rect 754 2833 763 2867
tri 860 2857 870 2867 ne
rect 711 2788 763 2833
rect 711 2754 720 2788
rect 754 2754 763 2788
rect 711 2709 763 2754
rect 711 2675 720 2709
rect 754 2675 763 2709
rect 711 2630 763 2675
rect 711 2596 720 2630
rect 754 2596 763 2630
rect 711 2551 763 2596
rect 711 2544 720 2551
rect 754 2544 763 2551
rect 711 2480 763 2492
rect 711 2393 763 2428
rect 711 2359 720 2393
rect 754 2359 763 2393
rect 711 2314 763 2359
rect 711 2280 720 2314
rect 754 2280 763 2314
rect 711 2234 763 2280
rect 711 2200 720 2234
rect 754 2200 763 2234
rect 711 2154 763 2200
rect 711 2120 720 2154
rect 754 2120 763 2154
rect 711 2108 763 2120
rect 870 2833 876 2867
rect 910 2833 916 2867
tri 916 2857 926 2867 nw
rect 870 2792 916 2833
rect 870 2758 876 2792
rect 910 2758 916 2792
rect 870 2717 916 2758
rect 870 2683 876 2717
rect 910 2683 916 2717
rect 870 2642 916 2683
rect 870 2608 876 2642
rect 910 2608 916 2642
rect 870 2567 916 2608
rect 870 2533 876 2567
rect 910 2533 916 2567
rect 870 2492 916 2533
rect 870 2458 876 2492
rect 910 2458 916 2492
rect 870 2417 916 2458
rect 870 2383 876 2417
rect 910 2383 916 2417
rect 870 2342 916 2383
rect 870 2308 876 2342
rect 910 2308 916 2342
rect 870 2267 916 2308
rect 870 2233 876 2267
rect 910 2233 916 2267
rect 870 2192 916 2233
rect 870 2158 876 2192
rect 910 2158 916 2192
rect 870 2117 916 2158
rect 424 2050 433 2084
rect 467 2050 476 2084
rect 870 2083 876 2117
rect 910 2083 916 2117
rect 424 2010 476 2050
rect 670 2028 676 2080
rect 728 2028 740 2080
rect 792 2028 798 2080
rect 870 2042 916 2083
rect 424 1976 433 2010
rect 467 1976 476 2010
tri 671 2008 691 2028 ne
rect 691 2008 773 2028
tri 773 2008 793 2028 nw
rect 870 2008 876 2042
rect 910 2008 916 2042
tri 691 1994 705 2008 ne
rect 424 1936 476 1976
rect 424 1902 433 1936
rect 467 1902 476 1936
rect 193 1844 250 1890
rect 204 1812 250 1844
rect 204 1778 210 1812
rect 244 1778 250 1812
rect 204 1735 250 1778
rect 204 1701 210 1735
rect 244 1701 250 1735
rect 204 1663 250 1701
rect 424 1862 476 1902
rect 424 1828 433 1862
rect 467 1828 476 1862
rect 705 1902 759 2008
tri 759 1994 773 2008 nw
rect 870 1967 916 2008
rect 870 1933 876 1967
rect 910 1933 916 1967
rect 870 1921 916 1933
rect 1023 2833 1032 2867
rect 1066 2833 1075 2867
rect 1023 2792 1075 2833
rect 1023 2758 1032 2792
rect 1066 2758 1075 2792
rect 1023 2717 1075 2758
rect 1023 2683 1032 2717
rect 1066 2683 1075 2717
rect 1023 2642 1075 2683
rect 1023 2608 1032 2642
rect 1066 2608 1075 2642
rect 1023 2567 1075 2608
rect 1023 2544 1032 2567
rect 1066 2544 1075 2567
rect 1023 2480 1032 2492
rect 1066 2480 1075 2492
rect 1023 2417 1075 2428
rect 1023 2383 1032 2417
rect 1066 2383 1075 2417
rect 1023 2342 1075 2383
rect 1023 2308 1032 2342
rect 1066 2308 1075 2342
rect 1023 2267 1075 2308
rect 1023 2233 1032 2267
rect 1066 2233 1075 2267
rect 1023 2192 1075 2233
rect 1023 2158 1032 2192
rect 1066 2158 1075 2192
rect 1023 2117 1075 2158
rect 1023 2083 1032 2117
rect 1066 2083 1075 2117
rect 1023 2042 1075 2083
rect 1023 2008 1032 2042
rect 1066 2008 1075 2042
rect 1023 1967 1075 2008
rect 1023 1933 1032 1967
rect 1066 1933 1075 1967
rect 1023 1921 1075 1933
rect 1133 2867 1185 2879
rect 1133 2833 1142 2867
rect 1176 2833 1185 2867
rect 1133 2792 1185 2833
rect 1133 2758 1142 2792
rect 1176 2758 1185 2792
rect 1133 2717 1185 2758
rect 1133 2683 1142 2717
rect 1176 2683 1185 2717
rect 1133 2642 1185 2683
rect 1133 2608 1142 2642
rect 1176 2608 1185 2642
rect 1133 2567 1185 2608
rect 1133 2533 1142 2567
rect 1176 2533 1185 2567
rect 1133 2492 1185 2533
rect 1133 2458 1142 2492
rect 1176 2458 1185 2492
rect 1133 2417 1185 2458
rect 1133 2383 1142 2417
rect 1176 2383 1185 2417
rect 1133 2342 1185 2383
rect 1133 2308 1142 2342
rect 1176 2308 1185 2342
rect 1133 2267 1185 2308
rect 1133 2233 1142 2267
rect 1176 2233 1185 2267
rect 1133 2231 1185 2233
rect 1133 2166 1142 2179
rect 1176 2166 1185 2179
rect 1133 2083 1142 2114
rect 1176 2083 1185 2114
rect 1133 2042 1185 2083
rect 1133 2008 1142 2042
rect 1176 2008 1185 2042
rect 1133 1967 1185 2008
rect 1133 1933 1142 1967
rect 1176 1933 1185 1967
rect 1133 1921 1185 1933
rect 1289 2867 1341 2933
rect 1289 2843 1298 2867
rect 1332 2843 1341 2867
rect 1289 2778 1298 2791
rect 1332 2778 1341 2791
rect 1289 2717 1341 2726
rect 1289 2713 1298 2717
rect 1332 2713 1341 2717
rect 1289 2648 1341 2661
rect 1289 2567 1341 2596
rect 1289 2533 1298 2567
rect 1332 2533 1341 2567
rect 1289 2492 1341 2533
rect 1289 2458 1298 2492
rect 1332 2458 1341 2492
rect 1289 2417 1341 2458
rect 1289 2383 1298 2417
rect 1332 2383 1341 2417
rect 1289 2342 1341 2383
rect 1289 2308 1298 2342
rect 1332 2308 1341 2342
rect 1289 2267 1341 2308
rect 1289 2233 1298 2267
rect 1332 2233 1341 2267
rect 1289 2192 1341 2233
rect 1289 2158 1298 2192
rect 1332 2158 1341 2192
rect 1289 2117 1341 2158
rect 1289 2083 1298 2117
rect 1332 2083 1341 2117
rect 1445 2867 1497 2879
rect 1445 2833 1454 2867
rect 1488 2833 1497 2867
rect 1445 2788 1497 2833
rect 1445 2754 1454 2788
rect 1488 2754 1497 2788
rect 1445 2709 1497 2754
rect 1445 2675 1454 2709
rect 1488 2675 1497 2709
rect 1445 2630 1497 2675
rect 1445 2596 1454 2630
rect 1488 2596 1497 2630
rect 1445 2551 1497 2596
rect 1445 2517 1454 2551
rect 1488 2517 1497 2551
rect 1445 2472 1497 2517
rect 1445 2438 1454 2472
rect 1488 2438 1497 2472
rect 1445 2393 1497 2438
rect 1445 2359 1454 2393
rect 1488 2359 1497 2393
rect 1445 2314 1497 2359
rect 1445 2280 1454 2314
rect 1488 2280 1497 2314
rect 1445 2234 1497 2280
rect 1445 2231 1454 2234
rect 1488 2231 1497 2234
rect 1445 2166 1497 2179
rect 1445 2108 1497 2114
rect 1601 2867 1653 2933
rect 1601 2843 1610 2867
rect 1644 2843 1653 2867
rect 1601 2778 1610 2791
rect 1644 2778 1653 2791
rect 1601 2717 1653 2726
rect 1601 2713 1610 2717
rect 1644 2713 1653 2717
rect 1601 2648 1653 2661
rect 1601 2567 1653 2596
rect 1601 2533 1610 2567
rect 1644 2533 1653 2567
rect 1601 2492 1653 2533
rect 1601 2458 1610 2492
rect 1644 2458 1653 2492
rect 1601 2417 1653 2458
rect 1601 2383 1610 2417
rect 1644 2383 1653 2417
rect 1601 2342 1653 2383
rect 1601 2308 1610 2342
rect 1644 2308 1653 2342
rect 1601 2267 1653 2308
rect 1601 2233 1610 2267
rect 1644 2233 1653 2267
rect 1601 2192 1653 2233
rect 1601 2158 1610 2192
rect 1644 2158 1653 2192
rect 1601 2117 1653 2158
rect 1289 2042 1341 2083
rect 1601 2083 1610 2117
rect 1644 2083 1653 2117
rect 1757 2867 1809 2879
rect 1757 2833 1766 2867
rect 1800 2833 1809 2867
rect 1757 2788 1809 2833
rect 1757 2754 1766 2788
rect 1800 2754 1809 2788
rect 1757 2709 1809 2754
rect 1757 2675 1766 2709
rect 1800 2675 1809 2709
rect 1757 2630 1809 2675
rect 1757 2596 1766 2630
rect 1800 2596 1809 2630
rect 1757 2551 1809 2596
rect 1757 2517 1766 2551
rect 1800 2517 1809 2551
rect 1757 2472 1809 2517
rect 1757 2438 1766 2472
rect 1800 2438 1809 2472
rect 1757 2393 1809 2438
rect 1757 2359 1766 2393
rect 1800 2359 1809 2393
rect 1757 2314 1809 2359
rect 1757 2280 1766 2314
rect 1800 2280 1809 2314
rect 1757 2234 1809 2280
rect 1757 2231 1766 2234
rect 1800 2231 1809 2234
rect 1757 2166 1809 2179
rect 1757 2108 1809 2114
rect 1913 2867 1965 2933
rect 4664 2901 4716 2941
rect 1913 2843 1922 2867
rect 1956 2843 1965 2867
rect 1913 2778 1922 2791
rect 1956 2778 1965 2791
rect 1913 2717 1965 2726
rect 1913 2713 1922 2717
rect 1956 2713 1965 2717
rect 1913 2648 1965 2661
rect 1913 2567 1965 2596
rect 1913 2533 1922 2567
rect 1956 2533 1965 2567
rect 1913 2492 1965 2533
rect 1913 2458 1922 2492
rect 1956 2458 1965 2492
rect 1913 2417 1965 2458
rect 1913 2383 1922 2417
rect 1956 2383 1965 2417
rect 1913 2342 1965 2383
rect 1913 2308 1922 2342
rect 1956 2308 1965 2342
rect 1913 2267 1965 2308
rect 1913 2233 1922 2267
rect 1956 2233 1965 2267
rect 1913 2192 1965 2233
rect 1913 2158 1922 2192
rect 1956 2158 1965 2192
rect 1913 2117 1965 2158
rect 1289 2008 1298 2042
rect 1332 2008 1341 2042
rect 1411 2028 1417 2080
rect 1469 2028 1481 2080
rect 1533 2028 1539 2080
rect 1601 2042 1653 2083
tri 1412 2008 1432 2028 ne
rect 1432 2008 1514 2028
tri 1514 2008 1534 2028 nw
rect 1601 2008 1610 2042
rect 1644 2008 1653 2042
rect 1289 1967 1341 2008
tri 1432 1994 1446 2008 ne
rect 1289 1933 1298 1967
rect 1332 1933 1341 1967
rect 1289 1921 1341 1933
tri 759 1902 770 1913 sw
tri 1435 1902 1446 1913 se
rect 1446 1902 1500 2008
tri 1500 1994 1514 2008 nw
rect 1601 1967 1653 2008
rect 1601 1933 1610 1967
rect 1644 1933 1653 1967
rect 1601 1921 1653 1933
rect 1913 2083 1922 2117
rect 1956 2083 1965 2117
rect 1913 2042 1965 2083
rect 1913 2008 1922 2042
rect 1956 2008 1965 2042
rect 1913 1967 1965 2008
rect 1913 1933 1922 1967
rect 1956 1933 1965 1967
rect 1913 1921 1965 1933
rect 2069 2867 2121 2879
rect 2069 2833 2078 2867
rect 2112 2833 2121 2867
rect 2069 2792 2121 2833
rect 2069 2758 2078 2792
rect 2112 2758 2121 2792
rect 2069 2717 2121 2758
rect 2069 2683 2078 2717
rect 2112 2683 2121 2717
rect 2069 2642 2121 2683
rect 2069 2608 2078 2642
rect 2112 2608 2121 2642
rect 2069 2567 2121 2608
rect 2069 2533 2078 2567
rect 2112 2533 2121 2567
rect 2069 2492 2121 2533
rect 2069 2458 2078 2492
rect 2112 2458 2121 2492
rect 2069 2417 2121 2458
rect 2069 2383 2078 2417
rect 2112 2383 2121 2417
rect 2069 2342 2121 2383
rect 2069 2308 2078 2342
rect 2112 2308 2121 2342
rect 2069 2267 2121 2308
rect 2069 2233 2078 2267
rect 2112 2233 2121 2267
rect 2069 2231 2121 2233
rect 2069 2166 2078 2179
rect 2112 2166 2121 2179
rect 2069 2083 2078 2114
rect 2112 2083 2121 2114
rect 2069 2042 2121 2083
rect 2069 2008 2078 2042
rect 2112 2008 2121 2042
rect 2069 1967 2121 2008
rect 2069 1933 2078 1967
rect 2112 1933 2121 1967
rect 2069 1921 2121 1933
rect 2225 2867 2277 2879
rect 2225 2833 2234 2867
rect 2268 2833 2277 2867
rect 2225 2792 2277 2833
rect 2225 2758 2234 2792
rect 2268 2758 2277 2792
rect 2225 2717 2277 2758
rect 2225 2683 2234 2717
rect 2268 2683 2277 2717
rect 2225 2642 2277 2683
rect 2225 2608 2234 2642
rect 2268 2608 2277 2642
rect 2225 2567 2277 2608
rect 2225 2533 2234 2567
rect 2268 2533 2277 2567
rect 2225 2492 2277 2533
rect 2225 2458 2234 2492
rect 2268 2458 2277 2492
rect 2225 2417 2277 2458
rect 2225 2388 2234 2417
rect 2268 2388 2277 2417
rect 2225 2324 2234 2336
rect 2268 2324 2277 2336
rect 2225 2267 2277 2272
rect 2225 2233 2234 2267
rect 2268 2233 2277 2267
rect 2225 2192 2277 2233
rect 2225 2158 2234 2192
rect 2268 2158 2277 2192
rect 2225 2117 2277 2158
rect 2225 2083 2234 2117
rect 2268 2083 2277 2117
rect 2225 2042 2277 2083
rect 2225 2008 2234 2042
rect 2268 2008 2277 2042
rect 2225 1967 2277 2008
rect 2225 1933 2234 1967
rect 2268 1933 2277 1967
rect 2225 1921 2277 1933
rect 2381 2867 2433 2879
rect 2381 2833 2390 2867
rect 2424 2833 2433 2867
rect 2381 2792 2433 2833
rect 2381 2758 2390 2792
rect 2424 2758 2433 2792
rect 2381 2717 2433 2758
rect 2381 2683 2390 2717
rect 2424 2683 2433 2717
rect 2381 2642 2433 2683
rect 2381 2608 2390 2642
rect 2424 2608 2433 2642
rect 2381 2567 2433 2608
rect 2381 2533 2390 2567
rect 2424 2533 2433 2567
rect 2381 2492 2433 2533
rect 2381 2458 2390 2492
rect 2424 2458 2433 2492
rect 2381 2417 2433 2458
rect 2381 2383 2390 2417
rect 2424 2383 2433 2417
rect 2381 2342 2433 2383
rect 2381 2308 2390 2342
rect 2424 2308 2433 2342
rect 2381 2267 2433 2308
rect 2381 2233 2390 2267
rect 2424 2233 2433 2267
rect 2381 2231 2433 2233
rect 2381 2166 2390 2179
rect 2424 2166 2433 2179
rect 2381 2083 2390 2114
rect 2424 2083 2433 2114
rect 2381 2042 2433 2083
rect 2381 2008 2390 2042
rect 2424 2008 2433 2042
rect 2381 1967 2433 2008
rect 2381 1933 2390 1967
rect 2424 1933 2433 1967
rect 2381 1921 2433 1933
rect 2537 2867 2589 2879
rect 2537 2833 2546 2867
rect 2580 2833 2589 2867
rect 2537 2792 2589 2833
rect 2537 2758 2546 2792
rect 2580 2758 2589 2792
rect 2537 2717 2589 2758
rect 2537 2683 2546 2717
rect 2580 2683 2589 2717
rect 2537 2642 2589 2683
rect 2537 2608 2546 2642
rect 2580 2608 2589 2642
rect 2537 2567 2589 2608
rect 2537 2533 2546 2567
rect 2580 2533 2589 2567
rect 2537 2492 2589 2533
rect 2537 2458 2546 2492
rect 2580 2458 2589 2492
rect 2537 2417 2589 2458
rect 2537 2388 2546 2417
rect 2580 2388 2589 2417
rect 2537 2324 2546 2336
rect 2580 2324 2589 2336
rect 2537 2267 2589 2272
rect 2537 2233 2546 2267
rect 2580 2233 2589 2267
rect 2537 2192 2589 2233
rect 2537 2158 2546 2192
rect 2580 2158 2589 2192
rect 2537 2117 2589 2158
rect 2537 2083 2546 2117
rect 2580 2083 2589 2117
rect 2537 2042 2589 2083
rect 2537 2008 2546 2042
rect 2580 2008 2589 2042
rect 2537 1967 2589 2008
rect 2537 1933 2546 1967
rect 2580 1933 2589 1967
rect 2537 1921 2589 1933
rect 2693 2867 2745 2879
rect 2693 2833 2702 2867
rect 2736 2833 2745 2867
rect 2693 2792 2745 2833
rect 2693 2758 2702 2792
rect 2736 2758 2745 2792
rect 2693 2717 2745 2758
rect 2693 2683 2702 2717
rect 2736 2683 2745 2717
rect 2693 2642 2745 2683
rect 2693 2608 2702 2642
rect 2736 2608 2745 2642
rect 2693 2567 2745 2608
rect 2693 2533 2702 2567
rect 2736 2533 2745 2567
rect 2693 2492 2745 2533
rect 2693 2458 2702 2492
rect 2736 2458 2745 2492
rect 2693 2417 2745 2458
rect 2693 2383 2702 2417
rect 2736 2383 2745 2417
rect 2693 2342 2745 2383
rect 2693 2308 2702 2342
rect 2736 2308 2745 2342
rect 2693 2267 2745 2308
rect 2693 2233 2702 2267
rect 2736 2233 2745 2267
rect 2693 2231 2745 2233
rect 2693 2166 2702 2179
rect 2736 2166 2745 2179
rect 2693 2083 2702 2114
rect 2736 2083 2745 2114
rect 2693 2042 2745 2083
rect 2693 2008 2702 2042
rect 2736 2008 2745 2042
rect 2693 1967 2745 2008
rect 2693 1933 2702 1967
rect 2736 1933 2745 1967
rect 2693 1921 2745 1933
rect 2849 2867 2901 2879
rect 2849 2833 2858 2867
rect 2892 2833 2901 2867
rect 2849 2792 2901 2833
rect 2849 2758 2858 2792
rect 2892 2758 2901 2792
rect 2849 2717 2901 2758
rect 2849 2683 2858 2717
rect 2892 2683 2901 2717
rect 2849 2642 2901 2683
rect 2849 2608 2858 2642
rect 2892 2608 2901 2642
rect 2849 2567 2901 2608
rect 2849 2544 2858 2567
rect 2892 2544 2901 2567
rect 2849 2480 2858 2492
rect 2892 2480 2901 2492
rect 2849 2417 2901 2428
rect 2849 2383 2858 2417
rect 2892 2383 2901 2417
rect 2849 2342 2901 2383
rect 2849 2308 2858 2342
rect 2892 2308 2901 2342
rect 2849 2267 2901 2308
rect 2849 2233 2858 2267
rect 2892 2233 2901 2267
rect 2849 2192 2901 2233
rect 2849 2158 2858 2192
rect 2892 2158 2901 2192
rect 2849 2117 2901 2158
rect 2849 2083 2858 2117
rect 2892 2083 2901 2117
rect 2849 2042 2901 2083
rect 2849 2008 2858 2042
rect 2892 2008 2901 2042
rect 2849 1967 2901 2008
rect 2849 1933 2858 1967
rect 2892 1933 2901 1967
rect 2849 1921 2901 1933
rect 3005 2867 3057 2879
rect 3005 2833 3014 2867
rect 3048 2833 3057 2867
rect 3005 2792 3057 2833
rect 3005 2758 3014 2792
rect 3048 2758 3057 2792
rect 3005 2717 3057 2758
rect 3005 2683 3014 2717
rect 3048 2683 3057 2717
rect 3005 2642 3057 2683
rect 3005 2608 3014 2642
rect 3048 2608 3057 2642
rect 3005 2567 3057 2608
rect 3005 2533 3014 2567
rect 3048 2533 3057 2567
rect 3005 2492 3057 2533
rect 3005 2458 3014 2492
rect 3048 2458 3057 2492
rect 3005 2417 3057 2458
rect 3005 2383 3014 2417
rect 3048 2383 3057 2417
rect 3005 2342 3057 2383
rect 3005 2308 3014 2342
rect 3048 2308 3057 2342
rect 3005 2267 3057 2308
rect 3005 2233 3014 2267
rect 3048 2233 3057 2267
rect 3005 2231 3057 2233
rect 3005 2166 3014 2179
rect 3048 2166 3057 2179
rect 3005 2083 3014 2114
rect 3048 2083 3057 2114
rect 3005 2042 3057 2083
rect 3005 2008 3014 2042
rect 3048 2008 3057 2042
rect 3005 1967 3057 2008
rect 3005 1933 3014 1967
rect 3048 1933 3057 1967
rect 3005 1921 3057 1933
rect 3161 2867 3213 2879
rect 3161 2833 3170 2867
rect 3204 2833 3213 2867
rect 3161 2792 3213 2833
rect 3161 2758 3170 2792
rect 3204 2758 3213 2792
rect 3161 2717 3213 2758
rect 3161 2683 3170 2717
rect 3204 2683 3213 2717
rect 3161 2642 3213 2683
rect 3161 2608 3170 2642
rect 3204 2608 3213 2642
rect 3161 2567 3213 2608
rect 3161 2544 3170 2567
rect 3204 2544 3213 2567
rect 3161 2480 3170 2492
rect 3204 2480 3213 2492
rect 3161 2417 3213 2428
rect 3161 2383 3170 2417
rect 3204 2383 3213 2417
rect 3161 2342 3213 2383
rect 3161 2308 3170 2342
rect 3204 2308 3213 2342
rect 3161 2267 3213 2308
rect 3161 2233 3170 2267
rect 3204 2233 3213 2267
rect 3161 2192 3213 2233
rect 3161 2158 3170 2192
rect 3204 2158 3213 2192
rect 3161 2117 3213 2158
rect 3161 2083 3170 2117
rect 3204 2083 3213 2117
rect 3161 2042 3213 2083
rect 3161 2008 3170 2042
rect 3204 2008 3213 2042
rect 3161 1967 3213 2008
rect 3161 1933 3170 1967
rect 3204 1933 3213 1967
rect 3161 1921 3213 1933
rect 3317 2867 3369 2879
rect 3317 2833 3326 2867
rect 3360 2833 3369 2867
rect 3317 2792 3369 2833
rect 3317 2758 3326 2792
rect 3360 2758 3369 2792
rect 3317 2717 3369 2758
rect 3317 2683 3326 2717
rect 3360 2683 3369 2717
rect 3317 2642 3369 2683
rect 3317 2608 3326 2642
rect 3360 2608 3369 2642
rect 3317 2567 3369 2608
rect 3317 2533 3326 2567
rect 3360 2533 3369 2567
rect 3317 2492 3369 2533
rect 3317 2458 3326 2492
rect 3360 2458 3369 2492
rect 3317 2417 3369 2458
rect 3317 2383 3326 2417
rect 3360 2383 3369 2417
rect 3317 2342 3369 2383
rect 3317 2308 3326 2342
rect 3360 2308 3369 2342
rect 3317 2267 3369 2308
rect 3317 2233 3326 2267
rect 3360 2233 3369 2267
rect 3317 2231 3369 2233
rect 3317 2166 3326 2179
rect 3360 2166 3369 2179
rect 3317 2083 3326 2114
rect 3360 2083 3369 2114
rect 3317 2042 3369 2083
rect 3317 2008 3326 2042
rect 3360 2008 3369 2042
rect 3317 1967 3369 2008
rect 3317 1933 3326 1967
rect 3360 1933 3369 1967
rect 3317 1921 3369 1933
rect 3476 2867 3522 2879
rect 3476 2833 3482 2867
rect 3516 2833 3522 2867
rect 3476 2792 3522 2833
rect 3476 2758 3482 2792
rect 3516 2758 3522 2792
rect 3476 2717 3522 2758
rect 3476 2683 3482 2717
rect 3516 2683 3522 2717
rect 3476 2642 3522 2683
rect 3476 2608 3482 2642
rect 3516 2608 3522 2642
rect 3476 2567 3522 2608
rect 3476 2533 3482 2567
rect 3516 2533 3522 2567
rect 3476 2492 3522 2533
rect 3476 2458 3482 2492
rect 3516 2458 3522 2492
rect 3476 2417 3522 2458
rect 3476 2383 3482 2417
rect 3516 2383 3522 2417
rect 3476 2342 3522 2383
rect 3476 2308 3482 2342
rect 3516 2308 3522 2342
rect 3476 2267 3522 2308
rect 3476 2233 3482 2267
rect 3516 2233 3522 2267
rect 3476 2192 3522 2233
rect 3476 2158 3482 2192
rect 3516 2158 3522 2192
rect 3476 2117 3522 2158
rect 3476 2083 3482 2117
rect 3516 2083 3522 2117
rect 3476 2042 3522 2083
rect 3476 2008 3482 2042
rect 3516 2008 3522 2042
rect 3629 2867 3681 2879
rect 3629 2833 3638 2867
rect 3672 2833 3681 2867
rect 3629 2789 3681 2833
rect 3629 2755 3638 2789
rect 3672 2755 3681 2789
rect 3629 2711 3681 2755
rect 3629 2677 3638 2711
rect 3672 2677 3681 2711
rect 3629 2633 3681 2677
rect 3629 2599 3638 2633
rect 3672 2599 3681 2633
rect 3629 2554 3681 2599
rect 3629 2520 3638 2554
rect 3672 2520 3681 2554
rect 3629 2475 3681 2520
rect 3629 2441 3638 2475
rect 3672 2441 3681 2475
rect 3629 2396 3681 2441
rect 3629 2362 3638 2396
rect 3672 2362 3681 2396
rect 3629 2317 3681 2362
rect 3629 2283 3638 2317
rect 3672 2283 3681 2317
rect 3629 2238 3681 2283
rect 3629 2231 3638 2238
rect 3672 2231 3681 2238
rect 3629 2166 3681 2179
rect 3629 2080 3681 2114
rect 3629 2046 3638 2080
rect 3672 2046 3681 2080
tri 3522 2008 3554 2040 sw
rect 3629 2034 3681 2046
rect 3788 2867 3834 2879
rect 3788 2833 3794 2867
rect 3828 2833 3834 2867
rect 3788 2792 3834 2833
rect 3788 2758 3794 2792
rect 3828 2758 3834 2792
rect 3788 2717 3834 2758
rect 3788 2683 3794 2717
rect 3828 2683 3834 2717
rect 3788 2642 3834 2683
rect 3788 2608 3794 2642
rect 3828 2608 3834 2642
rect 3788 2567 3834 2608
rect 3788 2533 3794 2567
rect 3828 2533 3834 2567
rect 3788 2492 3834 2533
rect 3788 2458 3794 2492
rect 3828 2458 3834 2492
rect 3788 2417 3834 2458
rect 3788 2383 3794 2417
rect 3828 2383 3834 2417
rect 3788 2342 3834 2383
rect 3788 2308 3794 2342
rect 3828 2308 3834 2342
rect 3788 2267 3834 2308
rect 3788 2233 3794 2267
rect 3828 2233 3834 2267
rect 3788 2192 3834 2233
rect 3788 2158 3794 2192
rect 3828 2158 3834 2192
rect 3788 2117 3834 2158
rect 3788 2083 3794 2117
rect 3828 2083 3834 2117
rect 3788 2042 3834 2083
rect 3941 2867 3993 2879
rect 3941 2833 3950 2867
rect 3984 2833 3993 2867
rect 3941 2790 3993 2833
rect 3941 2756 3950 2790
rect 3984 2756 3993 2790
rect 3941 2712 3993 2756
rect 3941 2678 3950 2712
rect 3984 2678 3993 2712
rect 3941 2634 3993 2678
rect 3941 2600 3950 2634
rect 3984 2600 3993 2634
rect 3941 2556 3993 2600
rect 3941 2522 3950 2556
rect 3984 2522 3993 2556
rect 3941 2478 3993 2522
rect 3941 2444 3950 2478
rect 3984 2444 3993 2478
rect 3941 2400 3993 2444
rect 3941 2366 3950 2400
rect 3984 2366 3993 2400
rect 3941 2322 3993 2366
rect 3941 2288 3950 2322
rect 3984 2288 3993 2322
rect 3941 2244 3993 2288
rect 3941 2231 3950 2244
rect 3984 2231 3993 2244
rect 3941 2166 3993 2179
rect 3941 2088 3993 2114
rect 3941 2054 3950 2088
rect 3984 2054 3993 2088
rect 3941 2042 3993 2054
rect 4097 2867 4149 2879
rect 4097 2833 4106 2867
rect 4140 2833 4149 2867
rect 4664 2867 4673 2901
rect 4707 2867 4716 2901
rect 4097 2792 4149 2833
rect 4097 2758 4106 2792
rect 4140 2758 4149 2792
rect 4097 2717 4149 2758
rect 4097 2683 4106 2717
rect 4140 2683 4149 2717
rect 4097 2642 4149 2683
rect 4097 2608 4106 2642
rect 4140 2608 4149 2642
rect 4097 2567 4149 2608
rect 4097 2533 4106 2567
rect 4140 2533 4149 2567
rect 4292 2857 4344 2863
rect 4292 2793 4344 2805
rect 4292 2642 4344 2741
rect 4664 2827 4716 2867
rect 4664 2793 4673 2827
rect 4707 2793 4716 2827
rect 4664 2753 4716 2793
rect 4664 2719 4673 2753
rect 4707 2719 4716 2753
rect 4664 2679 4716 2719
rect 4664 2645 4673 2679
rect 4707 2645 4716 2679
tri 4344 2642 4345 2643 sw
rect 4292 2609 4345 2642
tri 4345 2609 4378 2642 sw
rect 4292 2603 4517 2609
rect 4292 2569 4304 2603
rect 4338 2569 4388 2603
rect 4422 2569 4471 2603
rect 4505 2569 4517 2603
rect 4292 2563 4517 2569
rect 4664 2605 4716 2645
rect 4664 2571 4673 2605
rect 4707 2571 4716 2605
rect 4097 2492 4149 2533
rect 4097 2458 4106 2492
rect 4140 2458 4149 2492
rect 4664 2531 4716 2571
rect 4664 2497 4673 2531
rect 4707 2497 4716 2531
rect 4097 2417 4149 2458
rect 4097 2383 4106 2417
rect 4140 2383 4149 2417
rect 4097 2342 4149 2383
rect 4097 2308 4106 2342
rect 4140 2308 4149 2342
rect 4097 2267 4149 2308
rect 4097 2233 4106 2267
rect 4140 2233 4149 2267
rect 4097 2192 4149 2233
rect 4097 2158 4106 2192
rect 4140 2158 4149 2192
rect 4097 2117 4149 2158
rect 4097 2083 4106 2117
rect 4140 2083 4149 2117
tri 4091 2042 4097 2048 se
rect 4097 2042 4149 2083
tri 3782 2034 3788 2040 se
rect 3788 2034 3794 2042
tri 3756 2008 3782 2034 se
rect 3782 2008 3794 2034
rect 3828 2008 3834 2042
tri 4090 2041 4091 2042 se
rect 4091 2041 4106 2042
tri 3834 2008 3867 2041 sw
tri 4057 2008 4090 2041 se
rect 4090 2008 4106 2041
rect 4140 2008 4149 2042
rect 3476 2006 3554 2008
tri 3554 2006 3556 2008 sw
tri 3754 2006 3756 2008 se
rect 3756 2006 3867 2008
tri 3867 2006 3869 2008 sw
tri 4055 2006 4057 2008 se
rect 4057 2006 4149 2008
rect 3476 1967 4149 2006
rect 3476 1933 3482 1967
rect 3516 1933 3794 1967
rect 3828 1933 4106 1967
rect 4140 1933 4149 1967
rect 3476 1921 4149 1933
rect 4210 2459 4256 2471
rect 4210 2425 4216 2459
rect 4250 2425 4256 2459
rect 4210 2377 4256 2425
rect 4210 2343 4216 2377
rect 4250 2343 4256 2377
rect 4210 2295 4256 2343
rect 4210 2261 4216 2295
rect 4250 2261 4256 2295
rect 4210 2213 4256 2261
rect 4210 2179 4216 2213
rect 4250 2179 4256 2213
rect 4210 2131 4256 2179
rect 4210 2097 4216 2131
rect 4250 2097 4256 2131
rect 4210 2049 4256 2097
rect 4210 2015 4216 2049
rect 4250 2015 4256 2049
rect 4210 1967 4256 2015
rect 4210 1933 4216 1967
rect 4250 1933 4256 1967
tri 3516 1913 3524 1921 ne
rect 3524 1913 3625 1921
tri 1500 1902 1511 1913 sw
tri 3524 1902 3535 1913 ne
rect 3535 1902 3625 1913
tri 3625 1902 3644 1921 nw
tri 4199 1902 4210 1913 se
rect 4210 1908 4256 1933
rect 4361 2459 4413 2471
rect 4361 2425 4372 2459
rect 4406 2425 4413 2459
rect 4361 2377 4413 2425
rect 4361 2343 4372 2377
rect 4406 2343 4413 2377
rect 4361 2295 4413 2343
rect 4361 2261 4372 2295
rect 4406 2261 4413 2295
rect 4361 2231 4413 2261
rect 4361 2166 4413 2179
rect 4361 2097 4372 2114
rect 4406 2097 4413 2114
rect 4361 2049 4413 2097
rect 4361 2015 4372 2049
rect 4406 2015 4413 2049
rect 4361 1967 4413 2015
rect 4361 1933 4372 1967
rect 4406 1933 4413 1967
rect 4361 1921 4413 1933
rect 4522 2459 4568 2471
rect 4522 2425 4528 2459
rect 4562 2425 4568 2459
rect 4522 2377 4568 2425
rect 4522 2343 4528 2377
rect 4562 2343 4568 2377
rect 4522 2295 4568 2343
rect 4522 2261 4528 2295
rect 4562 2261 4568 2295
rect 4522 2213 4568 2261
rect 4522 2179 4528 2213
rect 4562 2179 4568 2213
rect 4522 2131 4568 2179
rect 4522 2097 4528 2131
rect 4562 2097 4568 2131
rect 4522 2049 4568 2097
rect 4522 2015 4528 2049
rect 4562 2015 4568 2049
rect 4522 1967 4568 2015
rect 4522 1933 4528 1967
rect 4562 1933 4568 1967
tri 4256 1908 4261 1913 sw
rect 4210 1902 4261 1908
tri 4261 1902 4267 1908 sw
tri 4516 1902 4522 1908 se
rect 4522 1902 4568 1933
rect 705 1896 770 1902
tri 770 1896 776 1902 sw
tri 1429 1896 1435 1902 se
rect 1435 1896 1511 1902
tri 1511 1896 1517 1902 sw
tri 3535 1896 3541 1902 ne
rect 3541 1896 3619 1902
tri 3619 1896 3625 1902 nw
tri 4193 1896 4199 1902 se
rect 4199 1896 4267 1902
tri 4267 1896 4273 1902 sw
tri 4510 1896 4516 1902 se
rect 4516 1896 4568 1902
rect 705 1888 776 1896
tri 776 1888 784 1896 sw
tri 1421 1888 1429 1896 se
rect 1429 1888 1517 1896
tri 1517 1888 1525 1896 sw
tri 3541 1888 3549 1896 ne
rect 3549 1888 3611 1896
tri 3611 1888 3619 1896 nw
tri 4185 1888 4193 1896 se
rect 4193 1888 4273 1896
tri 4273 1888 4281 1896 sw
tri 4502 1888 4510 1896 se
rect 4510 1888 4568 1896
rect 705 1881 784 1888
tri 784 1881 791 1888 sw
tri 1414 1881 1421 1888 se
rect 1421 1887 1525 1888
tri 1525 1887 1526 1888 sw
tri 3549 1887 3550 1888 ne
rect 1421 1882 1526 1887
tri 1526 1882 1531 1887 sw
rect 1421 1881 1531 1882
tri 1531 1881 1532 1882 sw
rect 705 1879 791 1881
tri 791 1879 793 1881 sw
tri 1412 1879 1414 1881 se
rect 1414 1879 1532 1881
tri 1532 1879 1534 1881 sw
rect 705 1873 2016 1879
rect 705 1839 717 1873
rect 751 1839 817 1873
rect 851 1839 917 1873
rect 951 1839 1245 1873
rect 1279 1839 1318 1873
rect 1352 1839 1391 1873
rect 1425 1839 1464 1873
rect 1498 1839 1537 1873
rect 1571 1839 1610 1873
rect 1644 1839 1682 1873
rect 1716 1839 1754 1873
rect 1788 1839 1826 1873
rect 1860 1839 1898 1873
rect 1932 1839 1970 1873
rect 2004 1839 2016 1873
rect 705 1833 2016 1839
rect 2154 1873 2225 1882
rect 2154 1839 2166 1873
rect 2200 1839 2225 1873
rect 2154 1830 2225 1839
rect 2277 1830 2289 1882
rect 2341 1873 2575 1882
rect 2346 1839 2385 1873
rect 2419 1839 2457 1873
rect 2491 1839 2529 1873
rect 2563 1839 2575 1873
rect 2341 1830 2575 1839
rect 2750 1830 2756 1882
rect 2808 1830 2820 1882
rect 2872 1873 3304 1882
rect 2879 1839 2928 1873
rect 2962 1839 3011 1873
rect 3045 1839 3094 1873
rect 3128 1839 3176 1873
rect 3210 1839 3258 1873
rect 3292 1839 3304 1873
rect 2872 1830 3304 1839
rect 424 1788 476 1828
rect 424 1754 433 1788
rect 467 1754 476 1788
rect 424 1752 476 1754
tri 476 1752 478 1754 sw
rect 424 1744 478 1752
tri 478 1744 486 1752 sw
rect 424 1735 486 1744
tri 486 1735 495 1744 sw
rect 424 1729 495 1735
tri 495 1729 501 1735 sw
rect 821 1729 827 1781
rect 879 1729 891 1781
rect 943 1729 949 1781
rect 424 1720 501 1729
tri 501 1720 510 1729 sw
rect 424 1674 516 1720
rect 1029 1714 2207 1720
rect 1029 1680 1067 1714
rect 1101 1680 1144 1714
rect 1178 1680 1221 1714
rect 1255 1680 1298 1714
rect 1332 1680 1375 1714
rect 1409 1680 1451 1714
rect 1485 1680 1527 1714
rect 1561 1680 1603 1714
rect 1637 1680 1679 1714
rect 1713 1680 1755 1714
rect 1789 1680 1831 1714
rect 1865 1680 1907 1714
rect 1941 1680 1983 1714
rect 2017 1680 2059 1714
rect 2093 1680 2135 1714
rect 2169 1680 2207 1714
rect 1029 1674 2207 1680
rect 2358 1714 3506 1720
rect 2358 1680 2396 1714
rect 2430 1680 2476 1714
rect 2510 1680 2556 1714
rect 2590 1680 2636 1714
rect 2670 1680 2716 1714
rect 2750 1680 2795 1714
rect 2829 1680 2874 1714
rect 2908 1680 2984 1714
rect 3018 1680 3059 1714
rect 3093 1680 3134 1714
rect 3168 1680 3209 1714
rect 3243 1680 3284 1714
rect 3318 1680 3359 1714
rect 3393 1680 3434 1714
rect 3468 1680 3506 1714
rect 2358 1674 3506 1680
tri 158 1638 176 1656 sw
rect 3550 1649 3610 1888
tri 3610 1887 3611 1888 nw
tri 4184 1887 4185 1888 se
rect 4185 1887 4281 1888
tri 4281 1887 4282 1888 sw
tri 4501 1887 4502 1888 se
rect 4502 1887 4568 1888
tri 4178 1881 4184 1887 se
rect 4184 1881 4282 1887
tri 4282 1881 4288 1887 sw
tri 4495 1881 4501 1887 se
rect 4501 1881 4568 1887
tri 4176 1879 4178 1881 se
rect 4178 1879 4288 1881
tri 4288 1879 4290 1881 sw
tri 4493 1879 4495 1881 se
rect 4495 1879 4568 1881
rect 3649 1873 4568 1879
rect 3649 1839 3661 1873
rect 3695 1839 3734 1873
rect 3768 1839 3807 1873
rect 3841 1839 3880 1873
rect 3914 1839 3953 1873
rect 3987 1839 4025 1873
rect 4059 1839 4568 1873
rect 3649 1833 4568 1839
rect 4664 2457 4716 2497
rect 4664 2423 4673 2457
rect 4707 2423 4716 2457
rect 4664 2383 4716 2423
rect 4664 2349 4673 2383
rect 4707 2349 4716 2383
rect 4664 2309 4716 2349
rect 4664 2275 4673 2309
rect 4707 2275 4716 2309
rect 4664 2235 4716 2275
rect 4664 2231 4673 2235
rect 4707 2231 4716 2235
rect 4664 2166 4716 2179
rect 4664 2086 4716 2114
rect 4664 2052 4673 2086
rect 4707 2052 4716 2086
rect 4664 2011 4716 2052
rect 4664 1977 4673 2011
rect 4707 1977 4716 2011
rect 4890 3016 4896 3050
rect 4930 3016 5098 3050
rect 5132 3016 5138 3050
rect 5348 3049 6700 3055
tri 6858 3054 6859 3055 ne
rect 6859 3054 7039 3055
tri 6859 3052 6861 3054 ne
rect 6861 3052 6999 3054
rect 4890 2976 5138 3016
rect 4890 2942 4896 2976
rect 4930 2942 5098 2976
rect 5132 2942 5138 2976
rect 4890 2902 5138 2942
rect 4890 2868 4896 2902
rect 4930 2868 5098 2902
rect 5132 2868 5138 2902
rect 4890 2828 5138 2868
rect 4890 2794 4896 2828
rect 4930 2794 5098 2828
rect 5132 2794 5138 2828
rect 4890 2754 5138 2794
rect 4890 2720 4896 2754
rect 4930 2720 5098 2754
rect 5132 2720 5138 2754
rect 4890 2680 5138 2720
rect 4890 2646 4896 2680
rect 4930 2646 5098 2680
rect 5132 2646 5138 2680
rect 4890 2606 5138 2646
rect 4890 2572 4896 2606
rect 4930 2572 5098 2606
rect 5132 2572 5138 2606
rect 4890 2532 5138 2572
rect 4890 2498 4896 2532
rect 4930 2498 5098 2532
rect 5132 2498 5138 2532
rect 4890 2458 5138 2498
rect 4890 2424 4896 2458
rect 4930 2424 5098 2458
rect 5132 2424 5138 2458
rect 4890 2384 5138 2424
rect 4890 2350 4896 2384
rect 4930 2350 5098 2384
rect 5132 2350 5138 2384
rect 4890 2310 5138 2350
rect 4890 2276 4896 2310
rect 4930 2276 5098 2310
rect 5132 2276 5138 2310
rect 4890 2236 5138 2276
rect 4890 2202 4896 2236
rect 4930 2202 5098 2236
rect 5132 2202 5138 2236
rect 4890 2162 5138 2202
rect 4890 2161 5098 2162
rect 4890 2127 4896 2161
rect 4930 2128 5098 2161
rect 5132 2128 5138 2162
rect 4930 2127 5138 2128
rect 4890 2088 5138 2127
rect 4890 2086 5098 2088
rect 4890 2052 4896 2086
rect 4930 2054 5098 2086
rect 5132 2054 5138 2088
rect 4930 2052 5138 2054
rect 4890 2013 5138 2052
rect 4890 2011 5098 2013
rect 4664 1936 4716 1977
rect 4664 1902 4673 1936
rect 4707 1902 4716 1936
rect 4664 1861 4716 1902
tri 4020 1827 4026 1833 ne
rect 4026 1827 4128 1833
tri 4128 1827 4134 1833 nw
rect 4664 1827 4673 1861
rect 4707 1827 4716 1861
tri 4026 1824 4029 1827 ne
rect 4029 1824 4125 1827
tri 4125 1824 4128 1827 nw
tri 4029 1816 4037 1824 ne
rect 4037 1816 4117 1824
tri 4117 1816 4125 1824 nw
tri 4037 1808 4045 1816 ne
rect 4045 1808 4109 1816
tri 4109 1808 4117 1816 nw
tri 4045 1799 4054 1808 ne
tri 4033 1714 4054 1735 se
rect 4054 1714 4100 1808
tri 4100 1799 4109 1808 nw
rect 4664 1786 4716 1827
tri 4662 1752 4664 1754 se
rect 4664 1752 4673 1786
rect 4707 1752 4716 1786
tri 4654 1744 4662 1752 se
rect 4662 1744 4716 1752
tri 4645 1735 4654 1744 se
rect 4654 1735 4716 1744
tri 4630 1720 4645 1735 se
rect 4645 1720 4716 1735
tri 4020 1701 4033 1714 se
rect 4033 1701 4100 1714
tri 3610 1649 3616 1655 sw
rect 3972 1649 3978 1701
rect 4030 1649 4042 1701
rect 4094 1649 4100 1701
rect 4135 1714 4716 1720
rect 4135 1680 4173 1714
rect 4207 1680 4257 1714
rect 4291 1680 4341 1714
rect 4375 1680 4424 1714
rect 4458 1680 4507 1714
rect 4541 1680 4590 1714
rect 4624 1680 4716 1714
rect 4135 1674 4716 1680
rect 4787 1994 4839 2000
rect 4787 1930 4839 1942
rect 3550 1639 3616 1649
tri 3616 1639 3626 1649 sw
rect 3550 1638 3626 1639
tri 3626 1638 3627 1639 sw
tri 4786 1638 4787 1639 se
rect 4787 1638 4839 1878
tri 95 1636 97 1638 se
rect 97 1636 176 1638
tri 176 1636 178 1638 sw
rect 3550 1636 3627 1638
tri 3627 1636 3629 1638 sw
tri 4784 1636 4786 1638 se
rect 4786 1636 4839 1638
tri 80 1621 95 1636 se
rect 95 1621 178 1636
tri 178 1621 193 1636 sw
rect 3550 1621 3629 1636
tri 3629 1621 3644 1636 sw
tri 4769 1621 4784 1636 se
rect 4784 1621 4839 1636
rect 3550 1569 3556 1621
rect 3608 1569 3620 1621
rect 3672 1569 3678 1621
tri 4753 1605 4769 1621 se
rect 4769 1605 4839 1621
rect 3960 1559 4839 1605
rect 4890 1977 4896 2011
rect 4930 1979 5098 2011
rect 5132 1979 5138 2013
rect 4930 1977 5138 1979
rect 4890 1938 5138 1977
rect 4890 1936 5098 1938
rect 4890 1902 4896 1936
rect 4930 1904 5098 1936
rect 5132 1904 5138 1938
rect 4930 1902 5138 1904
rect 4890 1863 5138 1902
rect 5196 3013 5299 3019
rect 5196 2961 5221 3013
rect 5273 2961 5299 3013
rect 5196 2949 5299 2961
rect 5196 2897 5221 2949
rect 5273 2897 5299 2949
rect 5196 2701 5299 2897
rect 5196 2649 5221 2701
rect 5273 2649 5299 2701
rect 5196 2637 5299 2649
rect 5196 2585 5221 2637
rect 5273 2585 5299 2637
rect 5196 1902 5299 2585
rect 5348 3015 5443 3049
rect 5477 3015 5530 3049
rect 5564 3015 5640 3049
rect 5674 3015 5712 3049
rect 5746 3015 5784 3049
rect 5818 3015 5856 3049
rect 5890 3015 5928 3049
rect 5962 3015 6001 3049
rect 6035 3015 6074 3049
rect 6108 3015 6147 3049
rect 6181 3015 6220 3049
rect 6254 3015 6293 3049
rect 6327 3015 6366 3049
rect 6400 3015 6439 3049
rect 6473 3015 6512 3049
rect 6546 3015 6585 3049
rect 6619 3015 6700 3049
tri 6861 3042 6871 3052 ne
rect 5348 3009 6700 3015
rect 5348 2982 5407 3009
tri 5407 2982 5434 3009 nw
tri 6614 2982 6641 3009 ne
rect 6641 2982 6700 3009
rect 5348 2981 5406 2982
tri 5406 2981 5407 2982 nw
tri 6641 2981 6642 2982 ne
rect 6642 2981 6700 2982
rect 5348 2978 5403 2981
tri 5403 2978 5406 2981 nw
tri 6642 2978 6645 2981 ne
rect 6645 2978 6700 2981
rect 5348 2977 5400 2978
rect 5348 2943 5357 2977
rect 5391 2943 5400 2977
tri 5400 2975 5403 2978 nw
tri 6645 2975 6648 2978 ne
rect 6648 2975 6700 2978
rect 5348 2902 5400 2943
rect 5348 2868 5357 2902
rect 5391 2868 5400 2902
rect 5620 2891 5626 2943
rect 5678 2891 5690 2943
rect 5742 2891 5748 2943
rect 6648 2941 6657 2975
rect 6691 2941 6700 2975
rect 6648 2901 6700 2941
tri 5620 2879 5632 2891 ne
rect 5632 2879 5720 2891
tri 5720 2879 5732 2891 nw
rect 5348 2827 5400 2868
rect 5348 2793 5357 2827
rect 5391 2793 5400 2827
rect 5348 2752 5400 2793
rect 5348 2718 5357 2752
rect 5391 2718 5400 2752
rect 5348 2701 5400 2718
rect 5348 2643 5357 2649
rect 5391 2643 5400 2649
rect 5348 2637 5400 2643
rect 5348 2568 5357 2585
rect 5391 2568 5400 2585
rect 5348 2528 5400 2568
rect 5348 2494 5357 2528
rect 5391 2494 5400 2528
rect 5348 2454 5400 2494
rect 5348 2420 5357 2454
rect 5391 2420 5400 2454
rect 5348 2380 5400 2420
rect 5348 2346 5357 2380
rect 5391 2346 5400 2380
rect 5348 2306 5400 2346
rect 5348 2272 5357 2306
rect 5391 2272 5400 2306
rect 5348 2232 5400 2272
rect 5348 2198 5357 2232
rect 5391 2198 5400 2232
rect 5348 2158 5400 2198
rect 5348 2124 5357 2158
rect 5391 2124 5400 2158
rect 5348 2084 5400 2124
rect 5348 2050 5357 2084
rect 5391 2050 5400 2084
rect 5348 2010 5400 2050
rect 5348 1976 5357 2010
rect 5391 1976 5400 2010
rect 5348 1936 5400 1976
tri 5299 1902 5307 1910 sw
rect 5348 1902 5357 1936
rect 5391 1902 5400 1936
rect 5493 2867 5545 2879
tri 5632 2867 5644 2879 ne
rect 5644 2867 5708 2879
tri 5708 2867 5720 2879 nw
rect 5803 2867 5855 2879
rect 5493 2833 5502 2867
rect 5536 2833 5545 2867
tri 5644 2859 5652 2867 ne
rect 5493 2792 5545 2833
rect 5493 2758 5502 2792
rect 5536 2758 5545 2792
rect 5493 2717 5545 2758
rect 5493 2701 5502 2717
rect 5536 2701 5545 2717
rect 5493 2642 5545 2649
rect 5493 2637 5502 2642
rect 5536 2637 5545 2642
rect 5493 2567 5545 2585
rect 5493 2533 5502 2567
rect 5536 2533 5545 2567
rect 5493 2492 5545 2533
rect 5493 2458 5502 2492
rect 5536 2458 5545 2492
rect 5493 2417 5545 2458
rect 5493 2383 5502 2417
rect 5536 2383 5545 2417
rect 5493 2342 5545 2383
rect 5493 2308 5502 2342
rect 5536 2308 5545 2342
rect 5493 2267 5545 2308
rect 5493 2233 5502 2267
rect 5536 2233 5545 2267
rect 5493 2192 5545 2233
rect 5493 2158 5502 2192
rect 5536 2158 5545 2192
rect 5493 2117 5545 2158
rect 5493 2083 5502 2117
rect 5536 2083 5545 2117
rect 5652 2833 5658 2867
rect 5692 2833 5698 2867
tri 5698 2857 5708 2867 nw
rect 5652 2788 5698 2833
rect 5652 2754 5658 2788
rect 5692 2754 5698 2788
rect 5652 2709 5698 2754
rect 5652 2675 5658 2709
rect 5692 2675 5698 2709
rect 5652 2630 5698 2675
rect 5652 2596 5658 2630
rect 5692 2596 5698 2630
rect 5652 2551 5698 2596
rect 5652 2517 5658 2551
rect 5692 2517 5698 2551
rect 5652 2472 5698 2517
rect 5652 2438 5658 2472
rect 5692 2438 5698 2472
rect 5652 2393 5698 2438
rect 5652 2359 5658 2393
rect 5692 2359 5698 2393
rect 5652 2314 5698 2359
rect 5652 2280 5658 2314
rect 5692 2280 5698 2314
rect 5652 2234 5698 2280
rect 5652 2200 5658 2234
rect 5692 2200 5698 2234
rect 5652 2154 5698 2200
rect 5652 2120 5658 2154
rect 5692 2120 5698 2154
rect 5652 2108 5698 2120
rect 5803 2833 5812 2867
rect 5846 2833 5855 2867
rect 5803 2792 5855 2833
rect 5803 2758 5812 2792
rect 5846 2758 5855 2792
rect 5803 2717 5855 2758
rect 5803 2701 5812 2717
rect 5846 2701 5855 2717
rect 5803 2642 5855 2649
rect 5803 2637 5812 2642
rect 5846 2637 5855 2642
rect 5803 2567 5855 2585
rect 5803 2533 5812 2567
rect 5846 2533 5855 2567
rect 5803 2492 5855 2533
rect 5803 2458 5812 2492
rect 5846 2458 5855 2492
rect 5803 2417 5855 2458
rect 5803 2383 5812 2417
rect 5846 2383 5855 2417
rect 5803 2342 5855 2383
rect 5803 2308 5812 2342
rect 5846 2308 5855 2342
rect 5803 2267 5855 2308
rect 5803 2233 5812 2267
rect 5846 2233 5855 2267
rect 5803 2192 5855 2233
rect 5803 2158 5812 2192
rect 5846 2158 5855 2192
rect 5803 2117 5855 2158
rect 5493 2042 5545 2083
rect 5803 2083 5812 2117
rect 5846 2083 5855 2117
rect 5493 2008 5502 2042
rect 5536 2008 5545 2042
rect 5493 1967 5545 2008
rect 5493 1933 5502 1967
rect 5536 1933 5545 1967
rect 5493 1921 5545 1933
rect 5613 2028 5619 2080
rect 5671 2028 5683 2080
rect 5735 2028 5741 2080
tri 5602 1902 5613 1913 se
rect 5613 1902 5741 2028
rect 5803 2042 5855 2083
rect 5803 2008 5812 2042
rect 5846 2008 5855 2042
rect 5803 1967 5855 2008
rect 5803 1933 5812 1967
rect 5846 1933 5855 1967
rect 5803 1921 5855 1933
rect 6021 2867 6073 2879
rect 6021 2857 6030 2867
rect 6064 2857 6073 2867
rect 6021 2793 6073 2805
rect 6021 2717 6073 2741
rect 6021 2683 6030 2717
rect 6064 2683 6073 2717
rect 6021 2642 6073 2683
rect 6021 2608 6030 2642
rect 6064 2608 6073 2642
rect 6021 2567 6073 2608
rect 6021 2533 6030 2567
rect 6064 2533 6073 2567
rect 6021 2492 6073 2533
rect 6021 2458 6030 2492
rect 6064 2458 6073 2492
rect 6021 2417 6073 2458
rect 6021 2383 6030 2417
rect 6064 2383 6073 2417
rect 6021 2342 6073 2383
rect 6021 2308 6030 2342
rect 6064 2308 6073 2342
rect 6021 2267 6073 2308
rect 6021 2233 6030 2267
rect 6064 2233 6073 2267
rect 6021 2192 6073 2233
rect 6021 2158 6030 2192
rect 6064 2158 6073 2192
rect 6021 2117 6073 2158
rect 6021 2083 6030 2117
rect 6064 2083 6073 2117
rect 6021 2042 6073 2083
rect 6021 2008 6030 2042
rect 6064 2008 6073 2042
rect 6021 1967 6073 2008
rect 6021 1933 6030 1967
rect 6064 1933 6073 1967
rect 6021 1921 6073 1933
rect 6237 2867 6289 2879
rect 6237 2833 6246 2867
rect 6280 2833 6289 2867
rect 6506 2867 6558 2880
rect 6237 2792 6289 2833
rect 6237 2758 6246 2792
rect 6280 2758 6289 2792
rect 6237 2717 6289 2758
rect 6237 2701 6246 2717
rect 6280 2701 6289 2717
rect 6237 2642 6289 2649
rect 6237 2637 6246 2642
rect 6280 2637 6289 2642
rect 6237 2567 6289 2585
rect 6237 2533 6246 2567
rect 6280 2533 6289 2567
rect 6237 2492 6289 2533
rect 6424 2857 6476 2863
rect 6424 2793 6476 2805
rect 6237 2458 6246 2492
rect 6280 2458 6289 2492
rect 6237 2417 6289 2458
rect 6237 2383 6246 2417
rect 6280 2383 6289 2417
rect 6237 2342 6289 2383
rect 6237 2308 6246 2342
rect 6280 2308 6289 2342
rect 6237 2267 6289 2308
rect 6237 2233 6246 2267
rect 6280 2233 6289 2267
rect 6237 2192 6289 2233
rect 6237 2158 6246 2192
rect 6280 2158 6289 2192
rect 6237 2117 6289 2158
rect 6237 2083 6246 2117
rect 6280 2083 6289 2117
rect 6237 2042 6289 2083
rect 6237 2008 6246 2042
rect 6280 2008 6289 2042
rect 6237 1967 6289 2008
rect 6237 1933 6246 1967
rect 6280 1933 6289 1967
rect 6237 1921 6289 1933
rect 6350 2509 6396 2521
rect 6350 2475 6356 2509
rect 6390 2475 6396 2509
rect 6350 2389 6396 2475
rect 6350 2355 6356 2389
rect 6390 2355 6396 2389
tri 5741 1902 5752 1913 sw
tri 5191 1896 5196 1901 se
rect 5196 1896 5307 1902
tri 5307 1896 5313 1902 sw
rect 4890 1861 5098 1863
rect 4890 1827 4896 1861
rect 4930 1829 5098 1861
rect 5132 1829 5138 1863
tri 5188 1893 5191 1896 se
rect 5191 1893 5313 1896
tri 5313 1893 5316 1896 sw
rect 5188 1841 5194 1893
rect 5246 1841 5258 1893
rect 5310 1841 5316 1893
tri 5188 1833 5196 1841 ne
rect 5196 1833 5308 1841
tri 5308 1833 5316 1841 nw
rect 5348 1862 5400 1902
tri 5596 1896 5602 1902 se
rect 5602 1896 5752 1902
tri 5752 1896 5758 1902 sw
tri 5588 1888 5596 1896 se
rect 5596 1888 5758 1896
tri 5758 1888 5766 1896 sw
tri 5581 1881 5588 1888 se
rect 5588 1881 5766 1888
tri 5766 1881 5773 1888 sw
tri 5579 1879 5581 1881 se
rect 5581 1879 5773 1881
tri 5773 1879 5775 1881 sw
rect 4930 1827 5138 1829
rect 4890 1788 5138 1827
rect 5196 1828 5303 1833
tri 5303 1828 5308 1833 nw
rect 5348 1828 5357 1862
rect 5391 1828 5400 1862
rect 5551 1873 5779 1879
rect 5551 1839 5563 1873
rect 5597 1839 5648 1873
rect 5682 1839 5733 1873
rect 5767 1839 5779 1873
rect 5551 1833 5779 1839
rect 5867 1873 6232 1879
rect 5867 1839 5879 1873
rect 5913 1839 5956 1873
rect 5990 1839 6033 1873
rect 6067 1839 6110 1873
rect 6144 1839 6186 1873
rect 6220 1839 6232 1873
rect 5867 1833 6232 1839
rect 5196 1827 5302 1828
tri 5302 1827 5303 1828 nw
rect 5196 1810 5299 1827
tri 5299 1824 5302 1827 nw
rect 4890 1786 5098 1788
rect 4890 1752 4896 1786
rect 4930 1754 5098 1786
rect 5132 1754 5138 1788
rect 4930 1752 5138 1754
rect 4890 1713 5138 1752
rect 4890 1711 5098 1713
rect 4890 1677 4896 1711
rect 4930 1679 5098 1711
rect 5132 1679 5138 1713
rect 4930 1677 5138 1679
rect 4890 1638 5138 1677
rect 5348 1788 5400 1828
tri 5908 1827 5914 1833 ne
rect 5914 1827 6098 1833
tri 6098 1827 6104 1833 nw
tri 5914 1824 5917 1827 ne
rect 5917 1824 6095 1827
tri 6095 1824 6098 1827 nw
tri 5917 1816 5925 1824 ne
rect 5925 1816 6087 1824
tri 6087 1816 6095 1824 nw
tri 5925 1808 5933 1816 ne
rect 5933 1808 6079 1816
tri 6079 1808 6087 1816 nw
tri 5933 1799 5942 1808 ne
rect 5348 1754 5357 1788
rect 5391 1754 5400 1788
rect 5348 1752 5400 1754
tri 5400 1752 5402 1754 sw
rect 5348 1744 5402 1752
tri 5402 1744 5410 1752 sw
rect 5348 1735 5410 1744
tri 5410 1735 5419 1744 sw
rect 5348 1720 5419 1735
tri 5419 1720 5434 1735 sw
rect 5348 1714 5826 1720
rect 5348 1680 5429 1714
rect 5463 1680 5511 1714
rect 5545 1680 5592 1714
rect 5626 1680 5673 1714
rect 5707 1680 5754 1714
rect 5788 1680 5826 1714
rect 5348 1674 5826 1680
rect 4890 1636 5098 1638
rect 4890 1602 4896 1636
rect 4930 1604 5098 1636
rect 5132 1604 5138 1638
rect 4930 1602 5138 1604
rect 4890 1563 5138 1602
rect 4890 1561 5098 1563
rect 3960 1527 4008 1559
tri 4008 1527 4040 1559 nw
rect 4890 1527 4896 1561
rect 4930 1529 5098 1561
rect 5132 1529 5138 1563
rect 4930 1527 5138 1529
rect 945 1490 2189 1496
rect 945 1456 957 1490
rect 991 1456 1031 1490
rect 1065 1456 1105 1490
rect 1139 1456 1179 1490
rect 1213 1456 1253 1490
rect 1287 1456 1327 1490
rect 1361 1456 1401 1490
rect 1435 1456 1475 1490
rect 1509 1456 1549 1490
rect 1583 1456 1623 1490
rect 1657 1456 1697 1490
rect 1731 1456 1771 1490
rect 1805 1456 1845 1490
rect 1879 1456 1919 1490
rect 1953 1456 1993 1490
rect 2027 1456 2068 1490
rect 2102 1456 2143 1490
rect 2177 1456 2189 1490
rect 945 1450 2189 1456
rect 2363 1490 3911 1496
rect 2363 1456 2375 1490
rect 2409 1456 2449 1490
rect 2483 1456 2523 1490
rect 2557 1456 2597 1490
rect 2631 1456 2671 1490
rect 2705 1456 2745 1490
rect 2779 1456 2819 1490
rect 2853 1456 2893 1490
rect 2927 1456 2967 1490
rect 3001 1456 3041 1490
rect 3075 1456 3115 1490
rect 3149 1456 3190 1490
rect 3224 1456 3265 1490
rect 3299 1456 3340 1490
rect 3374 1456 3415 1490
rect 3449 1456 3490 1490
rect 3524 1456 3565 1490
rect 3599 1456 3640 1490
rect 3674 1456 3715 1490
rect 3749 1456 3790 1490
rect 3824 1456 3865 1490
rect 3899 1456 3911 1490
rect 2363 1450 3911 1456
tri 2784 1230 2803 1249 ne
rect 2803 1230 2888 1249
tri 2888 1230 2907 1249 nw
tri 2803 1214 2819 1230 ne
rect 2005 1072 2026 1076
rect 1601 1066 2342 1072
rect 1601 1032 1613 1066
rect 1647 1032 1689 1066
rect 1723 1032 1765 1066
rect 1799 1032 1841 1066
rect 1875 1032 1917 1066
rect 1951 1032 1993 1066
rect 2027 1032 2069 1066
rect 2103 1032 2145 1066
rect 2179 1032 2221 1066
rect 2255 1032 2296 1066
rect 2330 1032 2342 1066
rect 1601 1026 2342 1032
rect 1812 908 1946 1026
rect 2005 873 2026 1026
rect 2819 843 2872 1230
tri 2872 1214 2888 1230 nw
tri 3928 1158 3960 1190 se
rect 3960 1158 4006 1527
tri 4006 1525 4008 1527 nw
rect 4890 1497 5138 1527
rect 5942 1541 6070 1808
tri 6070 1799 6079 1808 nw
tri 6329 1714 6350 1735 se
rect 6350 1714 6396 2355
rect 6424 2309 6476 2741
rect 6506 2833 6512 2867
rect 6546 2833 6558 2867
rect 6506 2788 6558 2833
rect 6506 2754 6512 2788
rect 6546 2754 6558 2788
rect 6506 2709 6558 2754
rect 6506 2701 6512 2709
rect 6546 2701 6558 2709
rect 6506 2637 6558 2649
rect 6506 2549 6558 2585
rect 6506 2515 6512 2549
rect 6546 2515 6558 2549
rect 6506 2469 6558 2515
rect 6506 2435 6512 2469
rect 6546 2435 6558 2469
rect 6506 2389 6558 2435
rect 6506 2355 6512 2389
rect 6546 2355 6558 2389
rect 6506 2343 6558 2355
rect 6648 2867 6657 2901
rect 6691 2867 6700 2901
rect 6648 2827 6700 2867
rect 6648 2793 6657 2827
rect 6691 2793 6700 2827
rect 6648 2753 6700 2793
rect 6648 2719 6657 2753
rect 6691 2719 6700 2753
rect 6648 2701 6700 2719
rect 6648 2645 6657 2649
rect 6691 2645 6700 2649
rect 6648 2637 6700 2645
rect 6648 2571 6657 2585
rect 6691 2571 6700 2585
rect 6648 2531 6700 2571
rect 6648 2497 6657 2531
rect 6691 2497 6700 2531
rect 6648 2457 6700 2497
rect 6648 2423 6657 2457
rect 6691 2423 6700 2457
rect 6648 2383 6700 2423
rect 6648 2349 6657 2383
rect 6691 2349 6700 2383
tri 6476 2309 6480 2313 sw
rect 6648 2309 6700 2349
rect 6424 2279 6480 2309
tri 6480 2279 6510 2309 sw
rect 6424 2273 6554 2279
rect 6424 2239 6436 2273
rect 6470 2239 6508 2273
rect 6542 2239 6554 2273
rect 6424 2233 6554 2239
rect 6648 2275 6657 2309
rect 6691 2275 6700 2309
rect 6648 2235 6700 2275
rect 6648 2201 6657 2235
rect 6691 2201 6700 2235
rect 6648 2161 6700 2201
rect 6648 2127 6657 2161
rect 6691 2127 6700 2161
rect 6648 2086 6700 2127
rect 6648 2052 6657 2086
rect 6691 2052 6700 2086
rect 6648 2011 6700 2052
rect 6648 1977 6657 2011
rect 6691 1977 6700 2011
rect 6648 1936 6700 1977
rect 6648 1902 6657 1936
rect 6691 1902 6700 1936
rect 6648 1861 6700 1902
rect 6648 1827 6657 1861
rect 6691 1827 6700 1861
rect 6648 1786 6700 1827
tri 6646 1752 6648 1754 se
rect 6648 1752 6657 1786
rect 6691 1752 6700 1786
tri 6638 1744 6646 1752 se
rect 6646 1744 6700 1752
tri 6629 1735 6638 1744 se
rect 6638 1735 6700 1744
tri 6614 1720 6629 1735 se
rect 6629 1720 6700 1735
tri 6316 1701 6329 1714 se
rect 6329 1701 6396 1714
rect 6268 1649 6274 1701
rect 6326 1649 6338 1701
rect 6390 1649 6396 1701
rect 6509 1714 6700 1720
rect 6509 1680 6566 1714
rect 6600 1680 6700 1714
rect 6509 1674 6700 1680
rect 6871 3018 6877 3052
rect 6911 3020 6999 3052
rect 7033 3020 7039 3054
rect 6911 3018 7039 3020
rect 6871 2981 7039 3018
rect 6871 2978 6999 2981
rect 6871 2944 6877 2978
rect 6911 2947 6999 2978
rect 7033 2947 7039 2981
rect 6911 2944 7039 2947
rect 6871 2908 7039 2944
rect 6871 2904 6999 2908
rect 6871 2870 6877 2904
rect 6911 2874 6999 2904
rect 7033 2874 7039 2908
rect 6911 2870 7039 2874
rect 6871 2835 7039 2870
rect 6871 2830 6999 2835
rect 6871 2796 6877 2830
rect 6911 2801 6999 2830
rect 7033 2801 7039 2835
rect 6911 2796 7039 2801
rect 6871 2762 7039 2796
rect 6871 2757 6999 2762
rect 6871 2723 6877 2757
rect 6911 2728 6999 2757
rect 7033 2728 7039 2762
rect 6911 2723 7039 2728
rect 6871 2689 7039 2723
rect 6871 2684 6999 2689
rect 6871 2650 6877 2684
rect 6911 2655 6999 2684
rect 7033 2655 7039 2689
rect 6911 2650 7039 2655
rect 6871 2616 7039 2650
rect 6871 2611 6999 2616
rect 6871 2577 6877 2611
rect 6911 2582 6999 2611
rect 7033 2582 7039 2616
rect 6911 2577 7039 2582
rect 6871 2543 7039 2577
rect 6871 2538 6999 2543
rect 6871 2504 6877 2538
rect 6911 2509 6999 2538
rect 7033 2509 7039 2543
rect 6911 2504 7039 2509
rect 6871 2470 7039 2504
rect 6871 2465 6999 2470
rect 6871 2431 6877 2465
rect 6911 2436 6999 2465
rect 7033 2436 7039 2470
rect 6911 2431 7039 2436
rect 6871 2397 7039 2431
rect 6871 2392 6999 2397
rect 6871 2358 6877 2392
rect 6911 2363 6999 2392
rect 7033 2363 7039 2397
rect 6911 2358 7039 2363
rect 6871 2324 7039 2358
rect 6871 2319 6999 2324
rect 6871 2285 6877 2319
rect 6911 2290 6999 2319
rect 7033 2290 7039 2324
rect 6911 2285 7039 2290
rect 6871 2251 7039 2285
rect 6871 2246 6999 2251
rect 6871 2212 6877 2246
rect 6911 2217 6999 2246
rect 7033 2217 7039 2251
rect 6911 2212 7039 2217
rect 6871 2178 7039 2212
rect 6871 2173 6999 2178
rect 6871 2139 6877 2173
rect 6911 2144 6999 2173
rect 7033 2144 7039 2178
rect 6911 2139 7039 2144
rect 6871 2105 7039 2139
rect 6871 2100 6999 2105
rect 6871 2066 6877 2100
rect 6911 2071 6999 2100
rect 7033 2071 7039 2105
rect 6911 2066 7039 2071
rect 6871 2032 7039 2066
rect 6871 2027 6999 2032
rect 6871 1993 6877 2027
rect 6911 1998 6999 2027
rect 7033 1998 7039 2032
rect 6911 1993 7039 1998
rect 6871 1960 7039 1993
rect 6871 1954 6999 1960
rect 6871 1920 6877 1954
rect 6911 1926 6999 1954
rect 7033 1926 7039 1960
rect 6911 1920 7039 1926
rect 6871 1888 7039 1920
rect 6871 1881 6999 1888
rect 6871 1847 6877 1881
rect 6911 1854 6999 1881
rect 7033 1854 7039 1888
rect 6911 1847 7039 1854
rect 6871 1816 7039 1847
rect 6871 1808 6999 1816
rect 6871 1774 6877 1808
rect 6911 1782 6999 1808
rect 7033 1782 7039 1816
rect 6911 1774 7039 1782
rect 6871 1744 7039 1774
rect 6871 1735 6999 1744
rect 6871 1701 6877 1735
rect 6911 1710 6999 1735
rect 7033 1710 7039 1744
rect 7216 3049 8838 3055
rect 7216 3015 7302 3049
rect 7336 3015 7380 3049
rect 7414 3015 7458 3049
rect 7492 3015 7536 3049
rect 7570 3015 7646 3049
rect 7680 3015 7722 3049
rect 7756 3015 7799 3049
rect 7833 3015 7876 3049
rect 7910 3015 7953 3049
rect 7987 3015 8030 3049
rect 8064 3015 8107 3049
rect 8141 3015 8184 3049
rect 8218 3015 8261 3049
rect 8295 3015 8338 3049
rect 8372 3015 8415 3049
rect 8449 3015 8492 3049
rect 8526 3015 8569 3049
rect 8603 3015 8646 3049
rect 8680 3015 8723 3049
rect 8757 3015 8838 3049
rect 7216 3009 8838 3015
rect 7216 2982 7275 3009
tri 7275 2982 7302 3009 nw
tri 8752 2982 8779 3009 ne
rect 8779 2982 8838 3009
rect 7216 2977 7269 2982
rect 7216 2943 7225 2977
rect 7259 2976 7269 2977
tri 7269 2976 7275 2982 nw
tri 8779 2976 8785 2982 ne
rect 8785 2976 8838 2982
rect 7259 2943 7268 2976
tri 7268 2975 7269 2976 nw
tri 8785 2975 8786 2976 ne
rect 8786 2975 8838 2976
rect 7216 2903 7268 2943
rect 7216 2869 7225 2903
rect 7259 2869 7268 2903
rect 8009 2912 8061 2924
rect 8131 2914 8137 2966
rect 8189 2914 8210 2966
rect 8262 2914 8283 2966
rect 8335 2914 8356 2966
rect 8408 2914 8429 2966
rect 8481 2914 8502 2966
rect 8554 2914 8560 2966
rect 7216 2829 7268 2869
rect 7216 2795 7225 2829
rect 7259 2795 7268 2829
rect 7216 2755 7268 2795
rect 7216 2721 7225 2755
rect 7259 2721 7268 2755
rect 7216 2700 7268 2721
rect 7216 2636 7268 2648
rect 7216 2575 7225 2584
rect 7259 2575 7268 2584
rect 7216 2536 7268 2575
rect 7216 2502 7225 2536
rect 7259 2502 7268 2536
rect 7216 2463 7268 2502
rect 7216 2429 7225 2463
rect 7259 2429 7268 2463
rect 7216 2390 7268 2429
rect 7216 2356 7225 2390
rect 7259 2356 7268 2390
rect 7216 2317 7268 2356
rect 7216 2283 7225 2317
rect 7259 2283 7268 2317
rect 7216 2244 7268 2283
rect 7216 2210 7225 2244
rect 7259 2210 7268 2244
rect 7216 2171 7268 2210
rect 7216 2137 7225 2171
rect 7259 2137 7268 2171
rect 7216 2098 7268 2137
rect 7216 2064 7225 2098
rect 7259 2064 7268 2098
rect 7216 2025 7268 2064
rect 7216 1991 7225 2025
rect 7259 1991 7268 2025
rect 7216 1952 7268 1991
rect 7216 1918 7225 1952
rect 7259 1918 7268 1952
rect 7361 2867 7413 2879
rect 7361 2857 7370 2867
rect 7404 2857 7413 2867
rect 7361 2793 7413 2805
rect 7361 2717 7413 2741
rect 7361 2683 7370 2717
rect 7404 2683 7413 2717
rect 7361 2642 7413 2683
rect 7361 2608 7370 2642
rect 7404 2608 7413 2642
rect 7361 2567 7413 2608
rect 7361 2533 7370 2567
rect 7404 2533 7413 2567
rect 7361 2492 7413 2533
rect 7361 2458 7370 2492
rect 7404 2458 7413 2492
rect 7361 2417 7413 2458
rect 7361 2383 7370 2417
rect 7404 2383 7413 2417
rect 7361 2342 7413 2383
rect 7361 2308 7370 2342
rect 7404 2308 7413 2342
rect 7361 2267 7413 2308
rect 7361 2233 7370 2267
rect 7404 2233 7413 2267
rect 7361 2192 7413 2233
rect 7361 2158 7370 2192
rect 7404 2158 7413 2192
rect 7361 2117 7413 2158
rect 7361 2083 7370 2117
rect 7404 2083 7413 2117
rect 7361 2042 7413 2083
rect 7361 2008 7370 2042
rect 7404 2008 7413 2042
rect 7361 1967 7413 2008
rect 7361 1933 7370 1967
rect 7404 1933 7413 1967
rect 7361 1921 7413 1933
rect 7577 2867 7629 2879
rect 7577 2833 7586 2867
rect 7620 2833 7629 2867
rect 7577 2792 7629 2833
rect 7577 2758 7586 2792
rect 7620 2758 7629 2792
rect 7577 2717 7629 2758
rect 7577 2700 7586 2717
rect 7620 2700 7629 2717
rect 7577 2642 7629 2648
rect 7577 2630 7586 2642
rect 7620 2630 7629 2642
rect 7577 2567 7629 2578
rect 7577 2560 7586 2567
rect 7620 2560 7629 2567
rect 7577 2492 7629 2508
rect 7577 2458 7586 2492
rect 7620 2458 7629 2492
rect 7577 2417 7629 2458
rect 7577 2383 7586 2417
rect 7620 2383 7629 2417
rect 7577 2342 7629 2383
rect 7577 2308 7586 2342
rect 7620 2308 7629 2342
rect 7577 2267 7629 2308
rect 7577 2233 7586 2267
rect 7620 2233 7629 2267
rect 7577 2192 7629 2233
rect 7577 2158 7586 2192
rect 7620 2158 7629 2192
rect 7577 2117 7629 2158
rect 7577 2083 7586 2117
rect 7620 2083 7629 2117
rect 7577 2042 7629 2083
rect 7577 2008 7586 2042
rect 7620 2008 7629 2042
rect 7577 1967 7629 2008
rect 7577 1933 7586 1967
rect 7620 1933 7629 1967
rect 7577 1921 7629 1933
rect 7793 2867 7845 2879
rect 7793 2857 7802 2867
rect 7836 2857 7845 2867
rect 7793 2793 7845 2805
rect 7793 2717 7845 2741
rect 7793 2683 7802 2717
rect 7836 2683 7845 2717
rect 7793 2642 7845 2683
rect 7793 2608 7802 2642
rect 7836 2608 7845 2642
rect 7793 2567 7845 2608
rect 7793 2533 7802 2567
rect 7836 2533 7845 2567
rect 7793 2492 7845 2533
rect 7793 2458 7802 2492
rect 7836 2458 7845 2492
rect 7793 2417 7845 2458
rect 7793 2383 7802 2417
rect 7836 2383 7845 2417
rect 7793 2342 7845 2383
rect 7793 2308 7802 2342
rect 7836 2308 7845 2342
rect 7793 2267 7845 2308
rect 7793 2233 7802 2267
rect 7836 2233 7845 2267
rect 7793 2192 7845 2233
rect 7793 2158 7802 2192
rect 7836 2158 7845 2192
rect 7793 2117 7845 2158
rect 7793 2083 7802 2117
rect 7836 2083 7845 2117
rect 7793 2042 7845 2083
rect 7793 2008 7802 2042
rect 7836 2008 7845 2042
rect 7793 1967 7845 2008
rect 7793 1933 7802 1967
rect 7836 1933 7845 1967
rect 7793 1921 7845 1933
rect 8009 2878 8018 2912
rect 8052 2878 8061 2912
tri 8134 2909 8139 2914 ne
rect 8139 2909 8243 2914
tri 8243 2909 8248 2914 nw
tri 8446 2909 8451 2914 ne
rect 8451 2909 8555 2914
tri 8555 2909 8560 2914 nw
rect 8786 2941 8795 2975
rect 8829 2941 8838 2975
tri 8139 2902 8146 2909 ne
rect 8146 2902 8236 2909
tri 8236 2902 8243 2909 nw
tri 8451 2902 8458 2909 ne
rect 8458 2902 8548 2909
tri 8548 2902 8555 2909 nw
tri 8146 2901 8147 2902 ne
rect 8147 2901 8235 2902
tri 8235 2901 8236 2902 nw
tri 8458 2901 8459 2902 ne
rect 8459 2901 8547 2902
tri 8547 2901 8548 2902 nw
rect 8786 2901 8838 2941
tri 8147 2880 8168 2901 ne
rect 8009 2840 8061 2878
rect 8009 2806 8018 2840
rect 8052 2806 8061 2840
rect 8009 2768 8061 2806
rect 8009 2734 8018 2768
rect 8052 2734 8061 2768
rect 8009 2700 8061 2734
rect 8009 2630 8061 2648
rect 8009 2560 8061 2578
rect 8009 2478 8061 2508
rect 8009 2444 8018 2478
rect 8052 2444 8061 2478
rect 8009 2405 8061 2444
rect 8009 2371 8018 2405
rect 8052 2371 8061 2405
rect 8009 2332 8061 2371
rect 8009 2298 8018 2332
rect 8052 2298 8061 2332
rect 8009 2259 8061 2298
rect 8009 2225 8018 2259
rect 8052 2225 8061 2259
rect 8009 2186 8061 2225
rect 8009 2152 8018 2186
rect 8052 2152 8061 2186
rect 8009 2113 8061 2152
rect 8009 2079 8018 2113
rect 8052 2079 8061 2113
rect 8168 2867 8214 2901
tri 8214 2880 8235 2901 nw
tri 8459 2880 8480 2901 ne
rect 8168 2833 8174 2867
rect 8208 2833 8214 2867
rect 8168 2788 8214 2833
rect 8168 2754 8174 2788
rect 8208 2754 8214 2788
rect 8168 2709 8214 2754
rect 8168 2675 8174 2709
rect 8208 2675 8214 2709
rect 8168 2630 8214 2675
rect 8168 2596 8174 2630
rect 8208 2596 8214 2630
rect 8168 2551 8214 2596
rect 8168 2517 8174 2551
rect 8208 2517 8214 2551
rect 8168 2472 8214 2517
rect 8168 2438 8174 2472
rect 8208 2438 8214 2472
rect 8168 2393 8214 2438
rect 8168 2359 8174 2393
rect 8208 2359 8214 2393
rect 8168 2314 8214 2359
rect 8168 2280 8174 2314
rect 8208 2280 8214 2314
rect 8168 2234 8214 2280
rect 8168 2200 8174 2234
rect 8208 2200 8214 2234
rect 8168 2154 8214 2200
rect 8168 2120 8174 2154
rect 8208 2120 8214 2154
rect 8168 2108 8214 2120
rect 8321 2867 8373 2879
rect 8321 2833 8330 2867
rect 8364 2833 8373 2867
rect 8321 2792 8373 2833
rect 8321 2758 8330 2792
rect 8364 2758 8373 2792
rect 8321 2717 8373 2758
rect 8321 2700 8330 2717
rect 8364 2700 8373 2717
rect 8321 2642 8373 2648
rect 8321 2630 8330 2642
rect 8364 2630 8373 2642
rect 8321 2567 8373 2578
rect 8321 2560 8330 2567
rect 8364 2560 8373 2567
rect 8321 2492 8373 2508
rect 8321 2458 8330 2492
rect 8364 2458 8373 2492
rect 8321 2417 8373 2458
rect 8321 2383 8330 2417
rect 8364 2383 8373 2417
rect 8321 2342 8373 2383
rect 8321 2308 8330 2342
rect 8364 2308 8373 2342
rect 8321 2267 8373 2308
rect 8321 2233 8330 2267
rect 8364 2233 8373 2267
rect 8321 2192 8373 2233
rect 8321 2158 8330 2192
rect 8364 2158 8373 2192
rect 8321 2117 8373 2158
rect 8321 2083 8330 2117
rect 8364 2083 8373 2117
rect 8480 2867 8526 2901
tri 8526 2880 8547 2901 nw
rect 8480 2833 8486 2867
rect 8520 2833 8526 2867
rect 8480 2788 8526 2833
rect 8480 2754 8486 2788
rect 8520 2754 8526 2788
rect 8480 2709 8526 2754
rect 8636 2867 8682 2879
rect 8636 2833 8642 2867
rect 8676 2833 8682 2867
rect 8636 2792 8682 2833
rect 8636 2758 8642 2792
rect 8676 2758 8682 2792
rect 8636 2717 8682 2758
rect 8480 2675 8486 2709
rect 8520 2675 8526 2709
rect 8480 2630 8526 2675
rect 8480 2596 8486 2630
rect 8520 2596 8526 2630
rect 8480 2551 8526 2596
rect 8480 2517 8486 2551
rect 8520 2517 8526 2551
rect 8480 2472 8526 2517
tri 8633 2706 8636 2709 se
rect 8636 2706 8642 2717
rect 8633 2700 8642 2706
rect 8676 2706 8682 2717
rect 8786 2867 8795 2901
rect 8829 2867 8838 2901
rect 8786 2827 8838 2867
rect 8786 2793 8795 2827
rect 8829 2793 8838 2827
rect 8786 2753 8838 2793
rect 8786 2719 8795 2753
rect 8829 2719 8838 2753
tri 8682 2706 8685 2709 sw
rect 8676 2700 8685 2706
rect 8633 2642 8685 2648
rect 8633 2630 8642 2642
rect 8676 2630 8685 2642
rect 8633 2567 8685 2578
rect 8633 2560 8642 2567
rect 8676 2560 8685 2567
rect 8633 2502 8685 2508
tri 8633 2499 8636 2502 ne
rect 8480 2438 8486 2472
rect 8520 2438 8526 2472
rect 8480 2393 8526 2438
rect 8480 2359 8486 2393
rect 8520 2359 8526 2393
rect 8480 2314 8526 2359
rect 8480 2280 8486 2314
rect 8520 2280 8526 2314
rect 8480 2234 8526 2280
rect 8480 2200 8486 2234
rect 8520 2200 8526 2234
rect 8480 2154 8526 2200
rect 8480 2120 8486 2154
rect 8520 2120 8526 2154
rect 8480 2108 8526 2120
rect 8636 2492 8682 2502
tri 8682 2499 8685 2502 nw
rect 8786 2700 8838 2719
rect 8786 2645 8795 2648
rect 8829 2645 8838 2648
rect 8786 2630 8838 2645
rect 8786 2571 8795 2578
rect 8829 2571 8838 2578
rect 8786 2560 8838 2571
rect 8636 2458 8642 2492
rect 8676 2458 8682 2492
rect 8636 2417 8682 2458
rect 8636 2383 8642 2417
rect 8676 2383 8682 2417
rect 8636 2342 8682 2383
rect 8636 2308 8642 2342
rect 8676 2308 8682 2342
rect 8636 2267 8682 2308
rect 8636 2233 8642 2267
rect 8676 2233 8682 2267
rect 8636 2192 8682 2233
rect 8636 2158 8642 2192
rect 8676 2158 8682 2192
rect 8636 2117 8682 2158
rect 8009 2040 8061 2079
rect 8009 2006 8018 2040
rect 8052 2006 8061 2040
rect 8127 2028 8133 2080
rect 8185 2028 8197 2080
rect 8249 2028 8255 2080
rect 8321 2042 8373 2083
rect 8636 2083 8642 2117
rect 8676 2083 8682 2117
tri 8128 2008 8148 2028 ne
rect 8148 2008 8230 2028
tri 8230 2008 8250 2028 nw
rect 8321 2008 8330 2042
rect 8364 2008 8373 2042
rect 8439 2028 8445 2080
rect 8497 2028 8509 2080
rect 8561 2028 8567 2080
rect 8636 2042 8682 2083
tri 8440 2008 8460 2028 ne
rect 8460 2008 8542 2028
tri 8542 2008 8562 2028 nw
rect 8636 2008 8642 2042
rect 8676 2008 8682 2042
rect 8009 1967 8061 2006
tri 8148 1994 8162 2008 ne
rect 8009 1933 8018 1967
rect 8052 1933 8061 1967
rect 8009 1921 8061 1933
rect 7216 1879 7268 1918
tri 8151 1902 8162 1913 se
rect 8162 1902 8216 2008
tri 8216 1994 8230 2008 nw
rect 8321 1967 8373 2008
tri 8460 1994 8474 2008 ne
rect 8321 1933 8330 1967
rect 8364 1933 8373 1967
rect 8321 1921 8373 1933
tri 8216 1902 8227 1913 sw
tri 8463 1902 8474 1913 se
rect 8474 1902 8528 2008
tri 8528 1994 8542 2008 nw
rect 8636 1967 8682 2008
rect 8636 1933 8642 1967
rect 8676 1933 8682 1967
rect 8636 1921 8682 1933
rect 8786 2497 8795 2508
rect 8829 2497 8838 2508
rect 8786 2457 8838 2497
rect 8786 2423 8795 2457
rect 8829 2423 8838 2457
rect 8786 2383 8838 2423
rect 8786 2349 8795 2383
rect 8829 2349 8838 2383
rect 8786 2309 8838 2349
rect 8786 2275 8795 2309
rect 8829 2275 8838 2309
rect 8786 2235 8838 2275
rect 8786 2201 8795 2235
rect 8829 2201 8838 2235
rect 8786 2161 8838 2201
rect 8786 2127 8795 2161
rect 8829 2127 8838 2161
rect 8786 2086 8838 2127
rect 8786 2052 8795 2086
rect 8829 2052 8838 2086
rect 8786 2011 8838 2052
rect 8786 1977 8795 2011
rect 8829 1977 8838 2011
rect 8786 1936 8838 1977
tri 8528 1902 8539 1913 sw
rect 8786 1902 8795 1936
rect 8829 1902 8838 1936
tri 8145 1896 8151 1902 se
rect 8151 1896 8227 1902
tri 8227 1896 8233 1902 sw
tri 8457 1896 8463 1902 se
rect 8463 1896 8539 1902
tri 8539 1896 8545 1902 sw
tri 8128 1879 8145 1896 se
rect 8145 1879 8233 1896
tri 8233 1879 8250 1896 sw
tri 8440 1879 8457 1896 se
rect 8457 1879 8545 1896
tri 8545 1879 8562 1896 sw
rect 7216 1845 7225 1879
rect 7259 1845 7268 1879
rect 7216 1806 7268 1845
rect 7439 1873 7960 1879
rect 7439 1839 7451 1873
rect 7485 1839 7529 1873
rect 7563 1839 7606 1873
rect 7640 1839 7683 1873
rect 7717 1839 7760 1873
rect 7794 1839 7837 1873
rect 7871 1839 7914 1873
rect 7948 1839 7960 1873
rect 7439 1833 7960 1839
rect 8089 1873 8613 1879
rect 8089 1839 8101 1873
rect 8135 1839 8179 1873
rect 8213 1839 8257 1873
rect 8291 1839 8335 1873
rect 8369 1839 8413 1873
rect 8447 1839 8490 1873
rect 8524 1839 8567 1873
rect 8601 1839 8613 1873
rect 8089 1833 8613 1839
rect 8786 1861 8838 1902
tri 7522 1827 7528 1833 ne
rect 7528 1827 7712 1833
tri 7712 1827 7718 1833 nw
rect 8786 1827 8795 1861
rect 8829 1827 8838 1861
tri 7528 1824 7531 1827 ne
rect 7531 1824 7709 1827
tri 7709 1824 7712 1827 nw
rect 7216 1772 7225 1806
rect 7259 1772 7268 1806
tri 7531 1799 7556 1824 ne
rect 7216 1734 7268 1772
rect 6911 1701 7039 1710
rect 6871 1672 7039 1701
rect 6871 1662 6999 1672
rect 4890 1495 5860 1497
rect 4074 1491 5860 1495
rect 4074 1489 5170 1491
rect 4074 1455 4112 1489
rect 4146 1455 4191 1489
rect 4225 1455 4270 1489
rect 4304 1455 4349 1489
rect 4383 1455 4428 1489
rect 4462 1455 4506 1489
rect 4540 1455 4584 1489
rect 4618 1455 4662 1489
rect 4696 1455 4740 1489
rect 4774 1455 4818 1489
rect 4852 1457 5170 1489
rect 5204 1457 5242 1491
rect 5276 1457 5314 1491
rect 5348 1457 5386 1491
rect 5420 1457 5458 1491
rect 5492 1457 5530 1491
rect 5564 1457 5602 1491
rect 5636 1457 5675 1491
rect 5709 1457 5748 1491
rect 5782 1457 5860 1491
rect 5942 1489 5948 1541
rect 6000 1489 6012 1541
rect 6064 1489 6070 1541
rect 6871 1628 6877 1662
rect 6911 1638 6999 1662
rect 7033 1638 7039 1672
rect 7211 1649 7217 1701
rect 7269 1649 7281 1701
rect 7333 1649 7339 1701
tri 7244 1638 7255 1649 ne
rect 7255 1638 7339 1649
rect 6911 1628 7039 1638
rect 6871 1600 7039 1628
tri 7255 1621 7272 1638 ne
rect 7272 1621 7339 1638
tri 7272 1614 7279 1621 ne
rect 6871 1589 6999 1600
rect 6871 1555 6877 1589
rect 6911 1566 6999 1589
rect 7033 1566 7039 1600
rect 6911 1555 7039 1566
rect 6871 1528 7039 1555
rect 6871 1498 6999 1528
rect 6157 1494 6999 1498
rect 7033 1494 7039 1528
rect 6157 1492 7039 1494
rect 4852 1455 5860 1457
rect 4074 1451 5860 1455
rect 4074 1449 5096 1451
rect 5814 1427 5860 1451
rect 6157 1458 6241 1492
rect 6275 1458 6319 1492
rect 6353 1458 6397 1492
rect 6431 1458 6476 1492
rect 6510 1458 6555 1492
rect 6589 1458 6634 1492
rect 6668 1458 6713 1492
rect 6747 1458 6792 1492
rect 6826 1458 6871 1492
rect 6905 1458 7039 1492
rect 6157 1456 7039 1458
rect 6157 1452 6993 1456
rect 6157 1427 6203 1452
rect 5814 1421 6203 1427
rect 5814 1387 5910 1421
rect 5944 1387 6000 1421
rect 6034 1387 6091 1421
rect 6125 1387 6203 1421
rect 5814 1381 6203 1387
tri 7245 1236 7279 1270 se
rect 7279 1236 7339 1621
rect 6726 1230 6856 1236
rect 6726 1196 6738 1230
rect 6772 1196 6810 1230
rect 6844 1196 6856 1230
rect 6726 1190 6856 1196
rect 7017 1230 7147 1236
rect 7017 1196 7029 1230
rect 7063 1196 7101 1230
rect 7135 1196 7147 1230
rect 7017 1190 7147 1196
rect 7209 1230 7339 1236
rect 7209 1196 7221 1230
rect 7255 1196 7293 1230
rect 7327 1196 7339 1230
tri 3926 1156 3928 1158 se
rect 3928 1156 4006 1158
rect 3794 1104 3800 1156
rect 3852 1104 3864 1156
rect 3916 1146 4006 1156
rect 3916 1112 3972 1146
tri 3972 1112 4006 1146 nw
rect 5894 1146 6592 1158
rect 5894 1112 6116 1146
rect 6150 1112 6548 1146
rect 6582 1112 6592 1146
rect 3916 1104 3964 1112
tri 3964 1104 3972 1112 nw
rect 5894 1106 6592 1112
rect 5894 1104 5957 1106
tri 5957 1104 5959 1106 nw
tri 6076 1104 6078 1106 ne
rect 6078 1104 6184 1106
rect 5894 1100 5953 1104
tri 5953 1100 5957 1104 nw
tri 6078 1100 6082 1104 ne
rect 6082 1100 6184 1104
tri 6184 1100 6190 1106 nw
tri 6506 1100 6512 1106 ne
rect 6512 1100 6592 1106
rect 5894 1094 5947 1100
tri 5947 1094 5953 1100 nw
tri 6082 1094 6088 1100 ne
rect 6088 1094 6158 1100
rect 4039 1082 4091 1094
rect 3431 1076 3711 1079
tri 3711 1076 3714 1079 sw
rect 3431 1074 3714 1076
tri 3714 1074 3716 1076 sw
rect 2954 1068 3429 1074
rect 2954 1034 2966 1068
rect 3000 1034 3049 1068
rect 3083 1034 3132 1068
rect 3166 1034 3215 1068
rect 3249 1034 3299 1068
rect 3333 1034 3383 1068
rect 3417 1034 3429 1068
rect 2954 1028 3429 1034
rect 3431 1048 3716 1074
tri 3716 1048 3742 1074 sw
rect 4039 1048 4048 1082
rect 4082 1048 4091 1082
rect 3431 1028 3742 1048
tri 3742 1028 3762 1048 sw
rect 3431 1026 3762 1028
tri 3762 1026 3764 1028 sw
rect 3431 1020 3764 1026
tri 3764 1020 3770 1026 sw
rect 3431 1019 3770 1020
tri 3770 1019 3771 1020 sw
rect 3933 1019 3985 1031
rect 3431 985 3771 1019
tri 3771 985 3805 1019 sw
rect 3933 985 3942 1019
rect 3976 985 3985 1019
rect 3431 984 3805 985
tri 3805 984 3806 985 sw
rect 3431 876 3806 984
tri 3637 873 3640 876 ne
rect 3640 873 3806 876
tri 2872 843 2902 873 sw
tri 3640 843 3670 873 ne
rect 3670 843 3806 873
rect 2254 832 2362 838
tri 2362 832 2368 838 sw
rect 2254 831 2368 832
tri 2368 831 2369 832 sw
rect 2819 831 3212 843
tri 3670 839 3674 843 ne
rect 3674 839 3806 843
tri 3674 838 3675 839 ne
rect 3675 838 3806 839
tri 3675 832 3681 838 ne
rect 3681 832 3806 838
rect 2254 826 2369 831
rect 2254 792 2260 826
rect 2294 823 2369 826
tri 2369 823 2377 831 sw
rect 2294 821 2377 823
tri 2377 821 2379 823 sw
rect 2294 797 2379 821
tri 2379 797 2403 821 sw
rect 2819 814 3172 831
tri 2819 797 2836 814 ne
rect 2836 797 3172 814
rect 3206 797 3212 831
tri 3681 825 3688 832 ne
rect 3688 825 3806 832
tri 3688 823 3690 825 ne
rect 2294 792 2403 797
rect 2254 766 2403 792
tri 2403 766 2434 797 sw
tri 2836 773 2860 797 ne
rect 2860 773 3212 797
tri 3117 766 3124 773 ne
rect 3124 766 3212 773
rect 2254 760 2434 766
tri 2434 760 2440 766 sw
tri 3124 760 3130 766 ne
rect 3130 760 3212 766
rect 2254 759 2440 760
tri 2440 759 2441 760 sw
tri 3130 759 3131 760 ne
rect 3131 759 3212 760
rect 2254 754 2441 759
rect 2254 720 2260 754
rect 2294 725 2441 754
tri 2441 725 2475 759 sw
tri 3131 725 3165 759 ne
rect 3165 725 3172 759
rect 3206 725 3212 759
rect 2294 720 2475 725
rect 2254 708 2475 720
tri 2475 708 2492 725 sw
tri 3165 724 3166 725 ne
rect 3166 713 3212 725
rect 2254 707 2492 708
tri 2353 693 2367 707 ne
rect 2367 693 2492 707
tri 2492 693 2507 708 sw
tri 2367 688 2372 693 ne
rect 2372 688 2507 693
tri 2507 688 2512 693 sw
tri 2372 685 2375 688 ne
rect 2375 685 2512 688
tri 2512 685 2515 688 sw
rect 472 678 2220 685
tri 2220 678 2227 685 sw
tri 2375 681 2379 685 ne
rect 2379 681 2515 685
tri 2515 681 2519 685 sw
tri 2379 678 2382 681 ne
rect 2382 678 3622 681
tri 3622 678 3625 681 sw
rect 472 663 2227 678
tri 2227 663 2242 678 sw
tri 2382 663 2397 678 ne
rect 2397 663 3625 678
tri 3625 663 3640 678 sw
rect 472 658 2242 663
tri 2242 658 2247 663 sw
tri 2397 658 2402 663 ne
rect 2402 658 3640 663
tri 3640 658 3645 663 sw
rect 472 654 2247 658
tri 2247 654 2251 658 sw
tri 2402 654 2406 658 ne
rect 2406 654 3645 658
tri 3645 654 3649 658 sw
rect 472 636 2251 654
tri 2251 636 2269 654 sw
tri 2406 650 2410 654 ne
rect 2410 650 3649 654
tri 3649 650 3653 654 sw
rect 472 633 2269 636
tri 2197 620 2210 633 ne
rect 2210 620 2269 633
tri 2410 629 2431 650 ne
rect 2431 629 3653 650
tri 3567 620 3576 629 ne
rect 3576 620 3653 629
tri 2210 616 2214 620 ne
rect 2214 616 2269 620
tri 3576 616 3580 620 ne
rect 3580 616 3653 620
tri 2214 609 2221 616 ne
rect 1886 593 1938 599
rect 1886 526 1938 541
rect 1679 448 1725 460
rect 1679 414 1685 448
rect 1719 414 1725 448
rect 1679 376 1725 414
rect 1886 456 1938 474
rect 2221 473 2269 616
tri 3580 606 3590 616 ne
rect 3590 606 3653 616
tri 3590 595 3601 606 ne
rect 3504 560 3556 566
tri 2269 473 2298 502 sw
rect 3504 485 3556 508
rect 2221 465 3125 473
tri 2221 461 2225 465 ne
rect 2225 461 3125 465
rect 1886 422 1895 456
rect 1929 422 1938 456
rect 1679 342 1685 376
rect 1719 342 1725 376
rect 1679 330 1725 342
rect 1783 399 1829 411
rect 1783 365 1789 399
rect 1823 365 1829 399
rect 1783 331 1829 365
rect 1886 383 1938 422
rect 1886 349 1895 383
rect 1929 349 1938 383
tri 1829 331 1841 343 sw
rect 1886 340 1938 349
rect 2145 449 2191 461
tri 2225 458 2228 461 ne
rect 2228 458 3125 461
tri 2228 455 2231 458 ne
rect 2231 455 3125 458
rect 2145 415 2151 449
rect 2185 415 2191 449
tri 2231 421 2265 455 ne
rect 2265 421 3085 455
rect 3119 421 3125 455
tri 2265 419 2267 421 ne
rect 2267 419 3125 421
rect 2145 377 2191 415
tri 3051 399 3071 419 ne
rect 3071 399 3125 419
tri 3071 397 3073 399 ne
rect 3073 397 3125 399
tri 3073 391 3079 397 ne
rect 2145 343 2151 377
rect 2185 343 2191 377
tri 1886 337 1889 340 ne
rect 1889 337 1935 340
tri 1935 337 1938 340 nw
tri 2139 337 2145 343 se
rect 2145 337 2191 343
rect 3079 383 3125 397
rect 3079 349 3085 383
rect 3119 349 3125 383
rect 3248 471 3300 477
rect 3248 407 3300 419
rect 3248 352 3257 355
rect 3291 352 3300 355
rect 3248 349 3300 352
rect 3504 410 3556 433
rect 3079 337 3125 349
rect 3251 340 3297 349
tri 2133 331 2139 337 se
rect 2139 331 2191 337
rect 1783 327 1841 331
rect 1783 293 1789 327
rect 1823 325 1841 327
tri 1841 325 1847 331 sw
tri 2127 325 2133 331 se
rect 2133 325 2191 331
rect 1823 324 1847 325
tri 1847 324 1848 325 sw
tri 2126 324 2127 325 se
rect 2127 324 2191 325
rect 1823 316 1848 324
tri 1848 316 1856 324 sw
tri 2118 316 2126 324 se
rect 2126 316 2191 324
rect 1823 309 1856 316
tri 1856 309 1863 316 sw
tri 2111 309 2118 316 se
rect 2118 309 2191 316
rect 1823 293 2191 309
rect 1783 281 2191 293
rect 3504 334 3556 358
rect 2000 230 2054 253
rect 1580 178 1586 230
rect 1638 178 1656 230
rect 1708 178 1726 230
rect 1778 178 1796 230
rect 1848 178 1866 230
rect 1918 178 1936 230
rect 1988 178 2006 230
rect 2058 178 2076 230
rect 2128 178 2146 230
rect 2198 178 2216 230
rect 2268 178 2285 230
rect 2337 178 2343 230
rect 1580 160 2343 178
rect 1580 108 1586 160
rect 1638 108 1656 160
rect 1708 108 1726 160
rect 1778 108 1796 160
rect 1848 108 1866 160
rect 1918 108 1936 160
rect 1988 108 2006 160
rect 2058 108 2076 160
rect 2128 108 2146 160
rect 2198 108 2216 160
rect 2268 108 2285 160
rect 2337 108 2343 160
rect 1580 90 2343 108
rect 1580 38 1586 90
rect 1638 82 1656 90
rect 1708 82 1726 90
rect 1778 82 1796 90
rect 1848 82 1866 90
rect 1918 82 1936 90
rect 1988 82 2006 90
rect 2058 82 2076 90
rect 2128 82 2146 90
rect 2198 82 2216 90
rect 1988 48 1992 82
rect 2058 48 2066 82
rect 2128 48 2140 82
rect 2198 48 2214 82
rect 1638 38 1656 48
rect 1708 38 1726 48
rect 1778 38 1796 48
rect 1848 38 1866 48
rect 1918 38 1936 48
rect 1988 38 2006 48
rect 2058 38 2076 48
rect 2128 38 2146 48
rect 2198 38 2216 48
rect 2268 38 2285 90
rect 2337 38 2343 90
rect 2953 178 2959 230
rect 3011 178 3029 230
rect 3081 178 3098 230
rect 3150 178 3167 230
rect 3219 178 3236 230
rect 3288 178 3305 230
rect 3357 178 3374 230
rect 3426 178 3432 230
rect 2953 160 3432 178
rect 2953 108 2959 160
rect 3011 108 3029 160
rect 3081 108 3098 160
rect 3150 108 3167 160
rect 3219 108 3236 160
rect 3288 108 3305 160
rect 3357 108 3374 160
rect 3426 108 3432 160
rect 2953 90 3432 108
rect 2953 38 2959 90
rect 3011 82 3029 90
rect 3081 82 3098 90
rect 3150 82 3167 90
rect 3219 82 3236 90
rect 3288 82 3305 90
rect 3357 82 3374 90
rect 3025 48 3029 82
rect 3357 48 3363 82
rect 3011 38 3029 48
rect 3081 38 3098 48
rect 3150 38 3167 48
rect 3219 38 3236 48
rect 3288 38 3305 48
rect 3357 38 3374 48
rect 3426 38 3432 90
rect 3504 132 3556 282
rect 3601 212 3653 606
rect 3690 560 3806 825
rect 3742 508 3754 560
rect 3690 485 3806 508
rect 3742 433 3754 485
rect 3690 410 3806 433
rect 3742 358 3754 410
rect 3690 334 3806 358
rect 3742 282 3754 334
rect 3690 276 3806 282
rect 3933 946 3985 985
rect 3933 912 3942 946
rect 3976 912 3985 946
rect 3933 873 3985 912
rect 3933 839 3942 873
rect 3976 839 3985 873
rect 3933 800 3985 839
rect 3933 766 3942 800
rect 3976 766 3985 800
rect 3933 727 3985 766
rect 3933 693 3942 727
rect 3976 693 3985 727
rect 3933 654 3985 693
rect 3933 620 3942 654
rect 3976 620 3985 654
rect 3933 581 3985 620
rect 3933 560 3942 581
rect 3976 560 3985 581
rect 3933 507 3985 508
rect 3933 484 3942 507
rect 3976 484 3985 507
rect 3933 409 3942 432
rect 3976 409 3985 432
rect 3933 334 3942 357
rect 3976 334 3985 357
rect 3933 251 3942 282
rect 3976 251 3985 282
rect 3933 239 3985 251
rect 4039 1010 4091 1048
rect 4039 976 4048 1010
rect 4082 976 4091 1010
rect 4039 949 4091 976
rect 4039 873 4091 897
rect 4039 798 4091 821
rect 4039 723 4091 746
rect 4039 650 4091 671
rect 4039 616 4048 650
rect 4082 616 4091 650
rect 4039 577 4091 616
rect 4039 543 4048 577
rect 4082 543 4091 577
rect 4039 504 4091 543
rect 4039 470 4048 504
rect 4082 470 4091 504
rect 4039 431 4091 470
rect 4039 397 4048 431
rect 4082 397 4091 431
rect 4039 358 4091 397
rect 4039 324 4048 358
rect 4082 324 4091 358
rect 4039 285 4091 324
rect 4039 251 4048 285
rect 4082 251 4091 285
rect 4039 239 4091 251
rect 4145 1082 4197 1094
rect 4145 1048 4154 1082
rect 4188 1048 4197 1082
rect 4145 1010 4197 1048
rect 4145 976 4154 1010
rect 4188 976 4197 1010
rect 4145 938 4197 976
rect 4145 904 4154 938
rect 4188 904 4197 938
rect 4145 866 4197 904
rect 4145 832 4154 866
rect 4188 832 4197 866
rect 4145 794 4197 832
rect 4145 760 4154 794
rect 4188 760 4197 794
rect 4145 722 4197 760
rect 4145 688 4154 722
rect 4188 688 4197 722
rect 4145 650 4197 688
rect 4145 616 4154 650
rect 4188 616 4197 650
rect 4145 577 4197 616
rect 4145 560 4154 577
rect 4188 560 4197 577
rect 4145 504 4197 508
rect 4145 484 4154 504
rect 4188 484 4197 504
rect 4145 431 4197 432
rect 4145 409 4154 431
rect 4188 409 4197 431
rect 4145 334 4154 357
rect 4188 334 4197 357
rect 4145 251 4154 282
rect 4188 251 4197 282
rect 4145 239 4197 251
rect 4251 1082 4303 1094
rect 4251 1048 4260 1082
rect 4294 1048 4303 1082
rect 4251 1010 4303 1048
rect 4251 976 4260 1010
rect 4294 976 4303 1010
rect 4251 949 4303 976
rect 4251 873 4303 897
rect 4251 798 4303 821
rect 4251 723 4303 746
rect 4251 650 4303 671
rect 4251 616 4260 650
rect 4294 616 4303 650
rect 4251 577 4303 616
rect 4251 543 4260 577
rect 4294 543 4303 577
rect 4251 504 4303 543
rect 4251 470 4260 504
rect 4294 470 4303 504
rect 4251 431 4303 470
rect 4251 397 4260 431
rect 4294 397 4303 431
rect 4251 358 4303 397
rect 4251 324 4260 358
rect 4294 324 4303 358
rect 4251 285 4303 324
rect 4251 251 4260 285
rect 4294 251 4303 285
rect 4251 239 4303 251
rect 4357 1082 4409 1094
rect 4357 1048 4366 1082
rect 4400 1048 4409 1082
rect 4357 1010 4409 1048
rect 4357 976 4366 1010
rect 4400 976 4409 1010
rect 4357 938 4409 976
rect 4357 904 4366 938
rect 4400 904 4409 938
rect 4357 866 4409 904
rect 4357 832 4366 866
rect 4400 832 4409 866
rect 4357 794 4409 832
rect 4357 760 4366 794
rect 4400 760 4409 794
rect 4357 722 4409 760
rect 4357 688 4366 722
rect 4400 688 4409 722
rect 4357 650 4409 688
rect 4357 616 4366 650
rect 4400 616 4409 650
rect 4357 577 4409 616
rect 4357 560 4366 577
rect 4400 560 4409 577
rect 4357 504 4409 508
rect 4357 484 4366 504
rect 4400 484 4409 504
rect 4357 431 4409 432
rect 4357 409 4366 431
rect 4400 409 4409 431
rect 4357 334 4366 357
rect 4400 334 4409 357
rect 4357 251 4366 282
rect 4400 251 4409 282
rect 4357 239 4409 251
rect 4463 1082 4515 1094
rect 4463 1048 4472 1082
rect 4506 1048 4515 1082
rect 4463 1010 4515 1048
rect 4463 976 4472 1010
rect 4506 976 4515 1010
rect 4463 949 4515 976
rect 4463 873 4515 897
rect 4463 798 4515 821
rect 4463 723 4515 746
rect 4463 650 4515 671
rect 4463 616 4472 650
rect 4506 616 4515 650
rect 4463 577 4515 616
rect 4463 543 4472 577
rect 4506 543 4515 577
rect 4463 504 4515 543
rect 4463 470 4472 504
rect 4506 470 4515 504
rect 4463 431 4515 470
rect 4463 397 4472 431
rect 4506 397 4515 431
rect 4463 358 4515 397
rect 4463 324 4472 358
rect 4506 324 4515 358
rect 4463 285 4515 324
rect 4463 251 4472 285
rect 4506 251 4515 285
rect 4463 239 4515 251
rect 4569 1082 4621 1094
rect 4569 1048 4578 1082
rect 4612 1048 4621 1082
rect 4569 1010 4621 1048
rect 4569 976 4578 1010
rect 4612 976 4621 1010
rect 4569 938 4621 976
rect 4569 904 4578 938
rect 4612 904 4621 938
rect 4569 866 4621 904
rect 4569 832 4578 866
rect 4612 832 4621 866
rect 4569 794 4621 832
rect 4569 760 4578 794
rect 4612 760 4621 794
rect 4569 722 4621 760
rect 4569 688 4578 722
rect 4612 688 4621 722
rect 4569 650 4621 688
rect 4569 616 4578 650
rect 4612 616 4621 650
rect 4569 577 4621 616
rect 4569 560 4578 577
rect 4612 560 4621 577
rect 4569 504 4621 508
rect 4569 484 4578 504
rect 4612 484 4621 504
rect 4569 431 4621 432
rect 4569 409 4578 431
rect 4612 409 4621 431
rect 4569 334 4578 357
rect 4612 334 4621 357
rect 4569 251 4578 282
rect 4612 251 4621 282
rect 4569 239 4621 251
rect 4675 1082 4727 1094
rect 4675 1048 4684 1082
rect 4718 1048 4727 1082
rect 4675 1010 4727 1048
rect 4675 976 4684 1010
rect 4718 976 4727 1010
rect 4675 949 4727 976
rect 4675 873 4727 897
rect 4675 798 4727 821
rect 4675 723 4727 746
rect 4675 650 4727 671
rect 4675 616 4684 650
rect 4718 616 4727 650
rect 4675 577 4727 616
rect 4675 543 4684 577
rect 4718 543 4727 577
rect 4675 504 4727 543
rect 4675 470 4684 504
rect 4718 470 4727 504
rect 4675 431 4727 470
rect 4675 397 4684 431
rect 4718 397 4727 431
rect 4675 358 4727 397
rect 4675 324 4684 358
rect 4718 324 4727 358
rect 4675 285 4727 324
rect 4675 251 4684 285
rect 4718 251 4727 285
rect 4675 239 4727 251
rect 4781 1082 4833 1094
rect 4781 1048 4790 1082
rect 4824 1048 4833 1082
rect 4781 1010 4833 1048
rect 4781 976 4790 1010
rect 4824 976 4833 1010
rect 4781 938 4833 976
rect 4781 904 4790 938
rect 4824 904 4833 938
rect 4781 866 4833 904
rect 4781 832 4790 866
rect 4824 832 4833 866
rect 4781 794 4833 832
rect 4781 760 4790 794
rect 4824 760 4833 794
rect 4781 722 4833 760
rect 4781 688 4790 722
rect 4824 688 4833 722
rect 4781 650 4833 688
rect 4781 616 4790 650
rect 4824 616 4833 650
rect 4781 577 4833 616
rect 4781 560 4790 577
rect 4824 560 4833 577
rect 4781 504 4833 508
rect 4781 484 4790 504
rect 4824 484 4833 504
rect 4781 431 4833 432
rect 4781 409 4790 431
rect 4824 409 4833 431
rect 4781 334 4790 357
rect 4824 334 4833 357
rect 4781 251 4790 282
rect 4824 251 4833 282
rect 4781 239 4833 251
rect 4887 1082 4939 1094
rect 4887 1048 4896 1082
rect 4930 1048 4939 1082
rect 4887 1010 4939 1048
rect 4887 976 4896 1010
rect 4930 976 4939 1010
rect 4887 949 4939 976
rect 4887 873 4939 897
rect 4887 798 4939 821
rect 4887 723 4939 746
rect 4887 650 4939 671
rect 4887 616 4896 650
rect 4930 616 4939 650
rect 4887 577 4939 616
rect 4887 543 4896 577
rect 4930 543 4939 577
rect 4887 504 4939 543
rect 4887 470 4896 504
rect 4930 470 4939 504
rect 4887 431 4939 470
rect 4887 397 4896 431
rect 4930 397 4939 431
rect 4887 358 4939 397
rect 4887 324 4896 358
rect 4930 324 4939 358
rect 4887 285 4939 324
rect 4887 251 4896 285
rect 4930 251 4939 285
rect 4887 239 4939 251
rect 4993 1082 5045 1094
rect 4993 1048 5002 1082
rect 5036 1048 5045 1082
rect 4993 1010 5045 1048
rect 4993 976 5002 1010
rect 5036 976 5045 1010
rect 4993 938 5045 976
rect 4993 904 5002 938
rect 5036 904 5045 938
rect 4993 866 5045 904
rect 4993 832 5002 866
rect 5036 832 5045 866
rect 4993 794 5045 832
rect 4993 760 5002 794
rect 5036 760 5045 794
rect 4993 722 5045 760
rect 4993 688 5002 722
rect 5036 688 5045 722
rect 4993 650 5045 688
rect 4993 616 5002 650
rect 5036 616 5045 650
rect 4993 577 5045 616
rect 4993 560 5002 577
rect 5036 560 5045 577
rect 4993 504 5045 508
rect 4993 484 5002 504
rect 5036 484 5045 504
rect 4993 431 5045 432
rect 4993 409 5002 431
rect 5036 409 5045 431
rect 4993 334 5002 357
rect 5036 334 5045 357
rect 4993 251 5002 282
rect 5036 251 5045 282
rect 4993 239 5045 251
rect 5099 1082 5151 1094
rect 5099 1048 5108 1082
rect 5142 1048 5151 1082
rect 5099 1010 5151 1048
rect 5099 976 5108 1010
rect 5142 976 5151 1010
rect 5099 949 5151 976
rect 5099 873 5151 897
rect 5099 798 5151 821
rect 5099 723 5151 746
rect 5099 650 5151 671
rect 5099 616 5108 650
rect 5142 616 5151 650
rect 5099 577 5151 616
rect 5099 543 5108 577
rect 5142 543 5151 577
rect 5099 504 5151 543
rect 5099 470 5108 504
rect 5142 470 5151 504
rect 5099 431 5151 470
rect 5099 397 5108 431
rect 5142 397 5151 431
rect 5099 358 5151 397
rect 5099 324 5108 358
rect 5142 324 5151 358
rect 5099 285 5151 324
rect 5099 251 5108 285
rect 5142 251 5151 285
rect 5099 239 5151 251
rect 5205 1082 5257 1094
rect 5205 1048 5214 1082
rect 5248 1048 5257 1082
rect 5205 1010 5257 1048
rect 5205 976 5214 1010
rect 5248 976 5257 1010
rect 5205 938 5257 976
rect 5205 904 5214 938
rect 5248 904 5257 938
rect 5205 866 5257 904
rect 5205 832 5214 866
rect 5248 832 5257 866
rect 5205 794 5257 832
rect 5205 760 5214 794
rect 5248 760 5257 794
rect 5205 722 5257 760
rect 5205 688 5214 722
rect 5248 688 5257 722
rect 5205 650 5257 688
rect 5205 616 5214 650
rect 5248 616 5257 650
rect 5205 577 5257 616
rect 5205 560 5214 577
rect 5248 560 5257 577
rect 5205 504 5257 508
rect 5205 484 5214 504
rect 5248 484 5257 504
rect 5205 431 5257 432
rect 5205 409 5214 431
rect 5248 409 5257 431
rect 5205 334 5214 357
rect 5248 334 5257 357
rect 5205 251 5214 282
rect 5248 251 5257 282
rect 5205 239 5257 251
rect 5311 1082 5363 1094
rect 5311 1048 5320 1082
rect 5354 1048 5363 1082
rect 5311 1010 5363 1048
rect 5311 976 5320 1010
rect 5354 976 5363 1010
rect 5311 949 5363 976
rect 5311 873 5363 897
rect 5311 798 5363 821
rect 5311 723 5363 746
rect 5311 650 5363 671
rect 5311 616 5320 650
rect 5354 616 5363 650
rect 5311 577 5363 616
rect 5311 543 5320 577
rect 5354 543 5363 577
rect 5311 504 5363 543
rect 5311 470 5320 504
rect 5354 470 5363 504
rect 5311 431 5363 470
rect 5311 397 5320 431
rect 5354 397 5363 431
rect 5311 358 5363 397
rect 5311 324 5320 358
rect 5354 324 5363 358
rect 5311 285 5363 324
rect 5311 251 5320 285
rect 5354 251 5363 285
rect 5311 239 5363 251
rect 5417 1082 5469 1094
rect 5417 1048 5426 1082
rect 5460 1048 5469 1082
rect 5417 1010 5469 1048
rect 5417 976 5426 1010
rect 5460 976 5469 1010
rect 5417 938 5469 976
rect 5417 904 5426 938
rect 5460 904 5469 938
rect 5417 866 5469 904
rect 5417 832 5426 866
rect 5460 832 5469 866
rect 5417 794 5469 832
rect 5417 760 5426 794
rect 5460 760 5469 794
rect 5417 722 5469 760
rect 5417 688 5426 722
rect 5460 688 5469 722
rect 5417 650 5469 688
rect 5417 616 5426 650
rect 5460 616 5469 650
rect 5417 577 5469 616
rect 5417 560 5426 577
rect 5460 560 5469 577
rect 5417 504 5469 508
rect 5417 484 5426 504
rect 5460 484 5469 504
rect 5417 431 5469 432
rect 5417 409 5426 431
rect 5460 409 5469 431
rect 5417 334 5426 357
rect 5460 334 5469 357
rect 5417 251 5426 282
rect 5460 251 5469 282
rect 5417 239 5469 251
rect 5523 1082 5575 1094
rect 5523 1048 5532 1082
rect 5566 1048 5575 1082
rect 5523 1010 5575 1048
rect 5523 976 5532 1010
rect 5566 976 5575 1010
rect 5523 949 5575 976
rect 5523 873 5575 897
rect 5523 798 5575 821
rect 5523 723 5575 746
rect 5523 650 5575 671
rect 5523 616 5532 650
rect 5566 616 5575 650
rect 5523 577 5575 616
rect 5523 543 5532 577
rect 5566 543 5575 577
rect 5523 504 5575 543
rect 5523 470 5532 504
rect 5566 470 5575 504
rect 5523 431 5575 470
rect 5523 397 5532 431
rect 5566 397 5575 431
rect 5523 358 5575 397
rect 5523 324 5532 358
rect 5566 324 5575 358
rect 5523 285 5575 324
rect 5523 251 5532 285
rect 5566 251 5575 285
rect 5523 239 5575 251
rect 5629 1082 5681 1094
rect 5629 1048 5638 1082
rect 5672 1048 5681 1082
rect 5629 1010 5681 1048
rect 5894 1054 5940 1094
tri 5940 1087 5947 1094 nw
tri 6088 1087 6095 1094 ne
rect 6095 1087 6158 1094
tri 6095 1074 6108 1087 ne
rect 6108 1074 6158 1087
tri 6158 1074 6184 1100 nw
tri 6512 1074 6538 1100 ne
rect 6538 1074 6592 1100
tri 6108 1072 6110 1074 ne
tri 5892 1020 5894 1022 se
rect 5894 1020 5900 1054
rect 5934 1020 5940 1054
rect 6110 1040 6116 1074
rect 6150 1040 6156 1074
tri 6156 1072 6158 1074 nw
tri 6538 1072 6540 1074 ne
rect 6110 1028 6156 1040
rect 6327 1054 6373 1066
tri 5940 1020 5942 1022 sw
tri 6325 1020 6327 1022 se
rect 6327 1020 6333 1054
rect 6367 1020 6373 1054
rect 6540 1040 6548 1074
rect 6582 1040 6592 1074
rect 5629 976 5638 1010
rect 5672 976 5681 1010
tri 5865 993 5892 1020 se
rect 5892 993 5942 1020
tri 5942 993 5969 1020 sw
tri 6298 993 6325 1020 se
rect 6325 993 6373 1020
tri 6373 993 6402 1022 sw
tri 5860 988 5865 993 se
rect 5865 988 5969 993
tri 5969 988 5974 993 sw
tri 6293 988 6298 993 se
rect 6298 988 6402 993
tri 6402 988 6407 993 sw
tri 5777 986 5779 988 se
rect 5779 986 6501 988
tri 5773 982 5777 986 se
rect 5777 982 6501 986
rect 5629 938 5681 976
tri 5739 948 5773 982 se
rect 5773 948 5900 982
rect 5934 948 6333 982
rect 6367 948 6501 982
rect 5629 904 5638 938
rect 5672 904 5681 938
rect 5629 866 5681 904
rect 5629 832 5638 866
rect 5672 832 5681 866
rect 5629 794 5681 832
rect 5629 760 5638 794
rect 5672 760 5681 794
rect 5629 722 5681 760
rect 5629 688 5638 722
rect 5672 688 5681 722
rect 5629 650 5681 688
rect 5629 616 5638 650
rect 5672 616 5681 650
rect 5629 577 5681 616
rect 5629 560 5638 577
rect 5672 560 5681 577
rect 5629 504 5681 508
rect 5629 484 5638 504
rect 5672 484 5681 504
rect 5629 431 5681 432
rect 5629 409 5638 431
rect 5672 409 5681 431
rect 5629 334 5638 357
rect 5672 334 5681 357
rect 5629 251 5638 282
rect 5672 251 5681 282
rect 5629 239 5681 251
tri 5730 939 5739 948 se
rect 5739 939 6501 948
rect 5730 900 6501 939
rect 5730 866 5957 900
rect 5991 866 6040 900
rect 6074 866 6123 900
rect 6157 866 6206 900
rect 6240 866 6289 900
rect 6323 866 6372 900
rect 6406 866 6455 900
rect 6489 866 6501 900
rect 5730 804 6501 866
rect 5730 770 5900 804
rect 5934 770 6333 804
rect 6367 770 6501 804
rect 5730 764 6501 770
rect 5730 744 5788 764
tri 5788 744 5808 764 nw
tri 5867 744 5887 764 ne
rect 5887 744 5954 764
tri 5954 744 5974 764 nw
tri 6293 744 6313 764 ne
rect 6313 744 6387 764
tri 6387 744 6407 764 nw
rect 5730 334 5782 744
tri 5782 738 5788 744 nw
tri 5887 738 5893 744 ne
rect 5893 738 5942 744
tri 5893 737 5894 738 ne
rect 5894 732 5942 738
tri 5942 732 5954 744 nw
tri 6313 732 6325 744 ne
rect 6325 732 6375 744
tri 6375 732 6387 744 nw
rect 5894 698 5900 732
rect 5934 698 5940 732
tri 5940 730 5942 732 nw
tri 6325 730 6327 732 ne
rect 5894 663 5940 698
rect 6110 712 6156 724
tri 6108 678 6110 680 se
rect 6110 678 6116 712
rect 6150 678 6156 712
rect 6327 698 6333 732
rect 6367 698 6373 732
tri 6373 730 6375 732 nw
rect 6327 686 6373 698
rect 6540 712 6592 1040
tri 6156 678 6158 680 sw
tri 6538 678 6540 680 se
rect 6540 678 6548 712
rect 6582 678 6592 712
tri 6094 664 6108 678 se
rect 6108 664 6158 678
tri 5940 663 5941 664 sw
tri 6093 663 6094 664 se
rect 6094 663 6158 664
tri 6158 663 6173 678 sw
tri 6523 663 6538 678 se
rect 6538 663 6592 678
rect 5894 658 5941 663
tri 5941 658 5946 663 sw
tri 6088 658 6093 663 se
rect 6093 658 6173 663
tri 6173 658 6178 663 sw
tri 6518 658 6523 663 se
rect 6523 658 6592 663
rect 5894 646 5946 658
tri 5946 646 5958 658 sw
tri 6076 646 6088 658 se
rect 6088 646 6178 658
tri 6178 646 6190 658 sw
tri 6506 646 6518 658 se
rect 6518 646 6592 658
rect 5894 640 6592 646
rect 5894 606 6116 640
rect 6150 606 6548 640
rect 6582 606 6592 640
rect 5894 594 6592 606
rect 6652 1100 6698 1112
rect 6652 1066 6658 1100
rect 6692 1066 6698 1100
rect 6652 1027 6698 1066
rect 6652 993 6658 1027
rect 6692 993 6698 1027
rect 6652 954 6698 993
rect 6652 920 6658 954
rect 6692 920 6698 954
rect 6726 1048 6778 1190
tri 6778 1156 6812 1190 nw
tri 7175 1112 7209 1146 se
rect 7209 1112 7339 1196
rect 6726 984 6778 996
rect 6726 926 6778 932
rect 6808 1100 7339 1112
rect 6808 1066 6814 1100
rect 6848 1066 7126 1100
rect 7160 1066 7339 1100
rect 6808 1052 7339 1066
rect 7386 1569 7392 1621
rect 7444 1569 7456 1621
rect 7508 1569 7514 1621
rect 7386 1563 7475 1569
tri 7475 1563 7481 1569 nw
rect 7386 1529 7441 1563
tri 7441 1529 7475 1563 nw
rect 7556 1541 7684 1824
tri 7684 1799 7709 1824 nw
rect 8786 1786 8838 1827
tri 8784 1752 8786 1754 se
rect 8786 1752 8795 1786
rect 8829 1752 8838 1786
tri 8754 1722 8784 1752 se
rect 8784 1722 8838 1752
tri 8752 1720 8754 1722 se
rect 8754 1720 8838 1722
rect 7742 1714 8838 1720
rect 7742 1680 7780 1714
rect 7814 1680 7853 1714
rect 7887 1680 7926 1714
rect 7960 1680 7999 1714
rect 8033 1680 8072 1714
rect 8106 1680 8145 1714
rect 8179 1680 8218 1714
rect 8252 1680 8291 1714
rect 8325 1680 8363 1714
rect 8397 1680 8435 1714
rect 8469 1680 8507 1714
rect 8541 1680 8579 1714
rect 8613 1680 8651 1714
rect 8685 1680 8723 1714
rect 8757 1680 8838 1714
rect 7742 1674 8838 1680
rect 9012 3050 9058 3090
rect 9012 3016 9018 3050
rect 9052 3016 9058 3050
rect 9012 2976 9058 3016
rect 9012 2942 9018 2976
rect 9052 2942 9058 2976
rect 9012 2902 9058 2942
rect 9012 2868 9018 2902
rect 9052 2868 9058 2902
rect 9012 2828 9058 2868
rect 9497 3245 9503 3297
rect 9555 3245 9639 3297
rect 9691 3245 9775 3297
rect 9827 3245 9911 3297
rect 9963 3245 10047 3297
rect 10099 3245 10183 3297
rect 10235 3245 10319 3297
rect 10371 3245 10455 3297
rect 10507 3245 10591 3297
rect 10643 3245 10727 3297
rect 10779 3245 10863 3297
rect 10915 3245 10999 3297
rect 11051 3245 11135 3297
rect 11187 3245 11271 3297
rect 11323 3245 11407 3297
rect 11459 3245 11542 3297
rect 11594 3245 11677 3297
rect 11729 3245 11735 3297
rect 9497 3187 11735 3245
rect 9497 3135 9503 3187
rect 9555 3135 9639 3187
rect 9691 3135 9775 3187
rect 9827 3135 9911 3187
rect 9963 3135 10047 3187
rect 10099 3135 10183 3187
rect 10235 3135 10319 3187
rect 10371 3135 10455 3187
rect 10507 3135 10591 3187
rect 10643 3135 10727 3187
rect 10779 3135 10863 3187
rect 10915 3135 10999 3187
rect 11051 3135 11135 3187
rect 11187 3135 11271 3187
rect 11323 3135 11407 3187
rect 11459 3135 11542 3187
rect 11594 3135 11677 3187
rect 11729 3135 11735 3187
rect 9497 3088 11735 3135
rect 9497 3054 9588 3088
rect 9622 3054 9673 3088
rect 9707 3054 9759 3088
rect 9793 3054 9845 3088
rect 9879 3054 9931 3088
rect 9965 3054 10041 3088
rect 10075 3054 10116 3088
rect 10150 3054 10191 3088
rect 10225 3054 10266 3088
rect 10300 3054 10341 3088
rect 10375 3054 10416 3088
rect 10450 3054 10491 3088
rect 10525 3054 10566 3088
rect 10600 3054 10641 3088
rect 10675 3054 10716 3088
rect 10750 3054 10791 3088
rect 10825 3054 10866 3088
rect 10900 3054 10941 3088
rect 10975 3054 11016 3088
rect 11050 3054 11091 3088
rect 11125 3054 11167 3088
rect 11201 3054 11243 3088
rect 11277 3054 11319 3088
rect 11353 3054 11395 3088
rect 11429 3054 11471 3088
rect 11505 3054 11547 3088
rect 11581 3054 11623 3088
rect 11657 3054 11735 3088
rect 9497 3016 11735 3054
rect 9497 2982 9503 3016
rect 9537 2982 11695 3016
rect 11729 2982 11735 3016
rect 9497 2944 11735 2982
rect 9497 2943 11695 2944
rect 9497 2909 9503 2943
rect 9537 2910 11695 2943
rect 11729 2910 11735 2944
rect 9537 2909 11735 2910
rect 9497 2875 9648 2909
rect 9682 2875 9960 2909
rect 9994 2875 10272 2909
rect 10306 2875 10584 2909
rect 10618 2875 10896 2909
rect 10930 2875 11208 2909
rect 11242 2875 11520 2909
rect 11554 2875 11735 2909
rect 9497 2872 11735 2875
rect 9497 2870 11695 2872
rect 9012 2794 9018 2828
rect 9052 2794 9058 2828
rect 9012 2754 9058 2794
rect 9012 2720 9018 2754
rect 9052 2720 9058 2754
rect 9012 2680 9058 2720
rect 9012 2646 9018 2680
rect 9052 2646 9058 2680
rect 9012 2606 9058 2646
rect 9012 2572 9018 2606
rect 9052 2572 9058 2606
rect 9012 2532 9058 2572
rect 9012 2498 9018 2532
rect 9052 2498 9058 2532
rect 9012 2458 9058 2498
rect 9012 2424 9018 2458
rect 9052 2424 9058 2458
rect 9012 2384 9058 2424
rect 9012 2350 9018 2384
rect 9052 2350 9058 2384
rect 9012 2310 9058 2350
rect 9012 2276 9018 2310
rect 9052 2276 9058 2310
rect 9012 2236 9058 2276
rect 9012 2202 9018 2236
rect 9052 2202 9058 2236
rect 9012 2162 9058 2202
rect 9012 2128 9018 2162
rect 9052 2128 9058 2162
rect 9012 2088 9058 2128
rect 9012 2054 9018 2088
rect 9052 2054 9058 2088
rect 9012 2013 9058 2054
rect 9012 1979 9018 2013
rect 9052 1979 9058 2013
rect 9012 1938 9058 1979
rect 9012 1904 9018 1938
rect 9052 1904 9058 1938
rect 9012 1863 9058 1904
rect 9012 1829 9018 1863
rect 9052 1829 9058 1863
rect 9012 1788 9058 1829
rect 9012 1754 9018 1788
rect 9052 1754 9058 1788
rect 9012 1713 9058 1754
rect 9012 1679 9018 1713
rect 9052 1679 9058 1713
rect 7386 1082 7432 1529
tri 7432 1520 7441 1529 nw
rect 7556 1489 7562 1541
rect 7614 1489 7626 1541
rect 7678 1489 7684 1541
rect 9012 1638 9058 1679
rect 9012 1604 9018 1638
rect 9052 1604 9058 1638
rect 9012 1563 9058 1604
tri 9010 1529 9012 1531 se
rect 9012 1529 9018 1563
rect 9052 1529 9058 1563
tri 8978 1497 9010 1529 se
rect 9010 1497 9058 1529
rect 7761 1491 9058 1497
rect 7761 1457 7799 1491
rect 7833 1457 7876 1491
rect 7910 1457 7953 1491
rect 7987 1457 8030 1491
rect 8064 1457 8106 1491
rect 8140 1457 8182 1491
rect 8216 1457 8258 1491
rect 8292 1457 8334 1491
rect 8368 1457 8410 1491
rect 8444 1457 8486 1491
rect 8520 1457 8562 1491
rect 8596 1457 8638 1491
rect 8672 1457 8714 1491
rect 8748 1457 8790 1491
rect 8824 1457 8866 1491
rect 8900 1457 8942 1491
rect 8976 1457 9058 1491
rect 7761 1451 9058 1457
rect 9097 2811 9103 2863
rect 9155 2811 9181 2863
rect 9233 2811 9239 2863
rect 9097 2787 9239 2811
rect 9097 2735 9103 2787
rect 9155 2735 9181 2787
rect 9233 2735 9239 2787
tri 9049 1337 9097 1385 se
rect 9097 1337 9239 2735
rect 9497 2836 9503 2870
rect 9537 2850 11695 2870
rect 9537 2838 9710 2850
tri 9710 2838 9722 2850 nw
tri 9920 2838 9932 2850 ne
rect 9932 2838 10022 2850
tri 10022 2838 10034 2850 nw
tri 10232 2838 10244 2850 ne
rect 10244 2838 10334 2850
tri 10334 2838 10346 2850 nw
tri 10544 2838 10556 2850 ne
rect 10556 2838 10646 2850
tri 10646 2838 10658 2850 nw
tri 10856 2838 10868 2850 ne
rect 10868 2838 10958 2850
tri 10958 2838 10970 2850 nw
tri 11168 2838 11180 2850 ne
rect 11180 2838 11270 2850
tri 11270 2838 11282 2850 nw
tri 11480 2838 11492 2850 ne
rect 11492 2838 11582 2850
tri 11582 2838 11594 2850 nw
tri 11655 2838 11667 2850 ne
rect 11667 2838 11695 2850
rect 11729 2838 11735 2872
rect 9537 2837 9709 2838
tri 9709 2837 9710 2838 nw
tri 9932 2837 9933 2838 ne
rect 9933 2837 10021 2838
tri 10021 2837 10022 2838 nw
tri 10244 2837 10245 2838 ne
rect 10245 2837 10333 2838
tri 10333 2837 10334 2838 nw
tri 10556 2837 10557 2838 ne
rect 10557 2837 10645 2838
tri 10645 2837 10646 2838 nw
tri 10868 2837 10869 2838 ne
rect 10869 2837 10957 2838
tri 10957 2837 10958 2838 nw
tri 11180 2837 11181 2838 ne
rect 11181 2837 11269 2838
tri 11269 2837 11270 2838 nw
tri 11492 2837 11493 2838 ne
rect 11493 2837 11560 2838
rect 9537 2836 9648 2837
rect 9497 2803 9648 2836
rect 9682 2803 9688 2837
tri 9688 2816 9709 2837 nw
tri 9933 2816 9954 2837 ne
rect 9497 2797 9688 2803
rect 9497 2763 9503 2797
rect 9537 2765 9688 2797
rect 9954 2803 9960 2837
rect 9994 2803 10000 2837
tri 10000 2816 10021 2837 nw
tri 10245 2816 10266 2837 ne
rect 9537 2763 9648 2765
rect 9497 2731 9648 2763
rect 9682 2731 9688 2765
rect 9497 2724 9688 2731
rect 9497 2690 9503 2724
rect 9537 2693 9688 2724
rect 9537 2690 9648 2693
rect 9497 2659 9648 2690
rect 9682 2659 9688 2693
rect 9497 2651 9688 2659
rect 9497 2617 9503 2651
rect 9537 2621 9688 2651
rect 9537 2617 9648 2621
rect 9497 2587 9648 2617
rect 9682 2587 9688 2621
rect 9497 2578 9688 2587
rect 9497 2544 9503 2578
rect 9537 2549 9688 2578
rect 9537 2544 9648 2549
rect 9497 2515 9648 2544
rect 9682 2515 9688 2549
rect 9497 2506 9688 2515
rect 8180 1273 9239 1337
rect 9270 2422 9276 2474
rect 9328 2422 9340 2474
rect 9392 2422 9398 2474
rect 9497 2472 9503 2506
rect 9537 2477 9688 2506
rect 9537 2472 9648 2477
rect 9497 2443 9648 2472
rect 9682 2443 9688 2477
rect 9497 2434 9688 2443
rect 9270 2400 9334 2422
tri 9334 2400 9356 2422 nw
rect 9497 2400 9503 2434
rect 9537 2405 9688 2434
rect 9537 2400 9648 2405
rect 8180 1270 8353 1273
tri 8353 1270 8356 1273 nw
tri 8146 1236 8180 1270 se
rect 8180 1236 8322 1270
tri 8322 1239 8353 1270 nw
rect 7580 1230 8322 1236
rect 7580 1196 7592 1230
rect 7626 1196 7668 1230
rect 7702 1196 7744 1230
rect 7778 1196 7820 1230
rect 7854 1196 7896 1230
rect 7930 1196 7972 1230
rect 8006 1196 8048 1230
rect 8082 1196 8124 1230
rect 8158 1196 8200 1230
rect 8234 1196 8276 1230
rect 8310 1196 8322 1230
rect 7580 1190 8322 1196
rect 8371 1230 8567 1236
rect 8371 1196 8383 1230
rect 8417 1196 8521 1230
rect 8555 1196 8567 1230
rect 8371 1190 8567 1196
tri 8146 1181 8155 1190 ne
rect 8155 1181 8322 1190
tri 8155 1156 8180 1181 ne
rect 6808 1048 6884 1052
tri 6884 1048 6888 1052 nw
tri 7086 1048 7090 1052 ne
rect 7090 1048 7196 1052
tri 7196 1048 7200 1052 nw
rect 7386 1048 7392 1082
rect 7426 1048 7432 1082
rect 6808 1020 6856 1048
tri 6856 1020 6884 1048 nw
tri 7090 1020 7118 1048 ne
rect 7118 1020 7167 1048
rect 6808 986 6814 1020
rect 6848 986 6854 1020
tri 6854 1018 6856 1020 nw
tri 7118 1018 7120 1020 ne
rect 6808 940 6854 986
rect 6652 880 6698 920
rect 6652 846 6658 880
rect 6692 846 6698 880
rect 6652 806 6698 846
rect 6652 772 6658 806
rect 6692 772 6698 806
rect 6652 732 6698 772
rect 6652 698 6658 732
rect 6692 698 6698 732
rect 6652 658 6698 698
rect 6652 624 6658 658
rect 6692 624 6698 658
rect 6652 584 6698 624
rect 6652 550 6658 584
rect 6692 550 6698 584
rect 6808 906 6814 940
rect 6848 906 6854 940
rect 6808 859 6854 906
rect 6808 825 6814 859
rect 6848 825 6854 859
rect 6808 778 6854 825
rect 6808 744 6814 778
rect 6848 744 6854 778
rect 6808 697 6854 744
rect 6808 663 6814 697
rect 6848 663 6854 697
rect 6808 616 6854 663
rect 6808 582 6814 616
rect 6848 582 6854 616
rect 6808 570 6854 582
rect 6964 986 7010 998
rect 6964 952 6970 986
rect 7004 952 7010 986
rect 6964 908 7010 952
rect 6964 874 6970 908
rect 7004 874 7010 908
rect 6964 830 7010 874
rect 6964 796 6970 830
rect 7004 796 7010 830
rect 6964 752 7010 796
rect 6964 718 6970 752
rect 7004 718 7010 752
rect 6964 674 7010 718
rect 6964 640 6970 674
rect 7004 640 7010 674
rect 6964 595 7010 640
rect 5860 528 6501 534
rect 5860 494 5957 528
rect 5991 494 6040 528
rect 6074 494 6123 528
rect 6157 494 6206 528
rect 6240 494 6289 528
rect 6323 494 6372 528
rect 6406 494 6455 528
rect 6489 494 6501 528
rect 5860 450 6501 494
rect 5860 416 5900 450
rect 5934 416 6332 450
rect 6366 416 6501 450
rect 5860 410 6501 416
rect 6652 510 6698 550
rect 6652 476 6658 510
rect 6692 482 6698 510
rect 6964 561 6970 595
rect 7004 561 7010 595
rect 7120 986 7126 1020
rect 7160 1019 7167 1020
tri 7167 1019 7196 1048 nw
rect 7160 986 7166 1019
tri 7166 1018 7167 1019 nw
rect 7386 1004 7432 1048
rect 7120 940 7166 986
rect 7120 906 7126 940
rect 7160 906 7166 940
rect 7120 859 7166 906
rect 7120 825 7126 859
rect 7160 825 7166 859
rect 7120 778 7166 825
rect 7120 744 7126 778
rect 7160 744 7166 778
rect 7120 697 7166 744
rect 7120 663 7126 697
rect 7160 663 7166 697
rect 7120 616 7166 663
rect 7120 582 7126 616
rect 7160 582 7166 616
rect 7120 570 7166 582
rect 7227 986 7279 999
rect 7227 952 7236 986
rect 7270 952 7279 986
rect 7227 912 7279 952
rect 7227 878 7236 912
rect 7270 878 7279 912
rect 7227 838 7279 878
rect 7227 804 7236 838
rect 7270 804 7279 838
rect 7227 764 7279 804
rect 7227 730 7236 764
rect 7270 730 7279 764
rect 7227 690 7279 730
rect 7227 656 7236 690
rect 7270 656 7279 690
rect 7227 616 7279 656
rect 7227 582 7236 616
rect 7270 582 7279 616
rect 6964 516 7010 561
tri 6698 482 6720 504 sw
tri 6942 482 6964 504 se
rect 6964 482 6970 516
rect 7004 502 7010 516
rect 7227 541 7279 582
rect 7227 507 7236 541
rect 7270 507 7279 541
tri 7010 502 7012 504 sw
tri 7225 502 7227 504 se
rect 7227 502 7279 507
rect 7004 494 7012 502
tri 7012 494 7020 502 sw
tri 7217 494 7225 502 se
rect 7225 494 7279 502
rect 7004 482 7020 494
rect 6692 476 6720 482
rect 6652 470 6720 476
tri 6720 470 6732 482 sw
tri 6930 470 6942 482 se
rect 6942 470 7020 482
tri 7020 470 7044 494 sw
tri 7193 470 7217 494 se
rect 7217 470 7279 494
rect 6652 466 7279 470
rect 6652 437 7236 466
rect 6652 436 6970 437
tri 5860 402 5868 410 ne
rect 5868 402 5966 410
tri 5966 402 5974 410 nw
tri 6292 402 6300 410 ne
rect 6300 402 6398 410
tri 6398 402 6406 410 nw
rect 6652 402 6658 436
rect 6692 403 6970 436
rect 7004 432 7236 437
rect 7270 432 7279 466
rect 7004 403 7279 432
rect 6692 402 7279 403
tri 5868 391 5879 402 ne
rect 5879 391 5955 402
tri 5955 391 5966 402 nw
tri 6300 391 6311 402 ne
rect 6311 391 6387 402
tri 6387 391 6398 402 nw
rect 6652 391 7279 402
tri 5879 390 5880 391 ne
rect 5880 390 5954 391
tri 5954 390 5955 391 nw
tri 6311 390 6312 391 ne
rect 6312 390 6386 391
tri 6386 390 6387 391 nw
rect 6652 390 7236 391
tri 5880 378 5892 390 ne
rect 5892 378 5942 390
tri 5942 378 5954 390 nw
tri 6312 378 6324 390 ne
rect 6324 378 6372 390
tri 5892 376 5894 378 ne
rect 5730 270 5782 282
rect 5894 344 5900 378
rect 5934 344 5940 378
tri 5940 376 5942 378 nw
tri 6324 376 6326 378 ne
rect 5894 326 5940 344
rect 6110 358 6156 370
tri 5940 326 5941 327 sw
rect 5894 324 5941 326
tri 5941 324 5943 326 sw
tri 6108 324 6110 326 se
rect 6110 324 6116 358
rect 6150 324 6156 358
rect 6326 344 6332 378
rect 6366 344 6372 378
tri 6372 376 6386 390 nw
tri 7193 376 7207 390 ne
rect 7207 376 7236 390
tri 7207 370 7213 376 ne
rect 7213 370 7236 376
rect 6326 332 6372 344
rect 6542 364 6594 370
tri 6156 324 6158 326 sw
tri 6540 324 6542 326 se
tri 7213 357 7226 370 ne
rect 7226 357 7236 370
rect 7270 357 7279 391
tri 7226 356 7227 357 ne
rect 5894 316 5943 324
tri 5943 316 5951 324 sw
tri 6100 316 6108 324 se
rect 6108 316 6158 324
tri 6158 316 6166 324 sw
tri 6532 316 6540 324 se
rect 6540 316 6542 324
rect 5894 292 5951 316
tri 5951 292 5975 316 sw
tri 6076 292 6100 316 se
rect 6100 292 6166 316
tri 6166 292 6190 316 sw
tri 6508 292 6532 316 se
rect 6532 312 6542 316
tri 6750 316 6769 335 se
rect 6769 316 6791 335
rect 6532 300 6594 312
rect 6532 292 6542 300
rect 5894 286 6542 292
rect 5894 252 6116 286
rect 6150 252 6542 286
tri 6717 283 6750 316 se
rect 6750 283 6791 316
rect 6843 283 6855 335
rect 6907 283 6913 335
rect 7227 316 7279 357
tri 6716 282 6717 283 se
rect 6717 282 6790 283
tri 6790 282 6791 283 nw
rect 7227 282 7236 316
rect 7270 282 7279 316
tri 6703 269 6716 282 se
rect 6716 269 6777 282
tri 6777 269 6790 282 nw
tri 6701 267 6703 269 se
rect 6703 267 6775 269
tri 6775 267 6777 269 nw
rect 5894 248 6542 252
rect 5894 240 6594 248
tri 6675 241 6701 267 se
rect 6701 241 6749 267
tri 6749 241 6775 267 nw
rect 7227 241 7279 282
tri 6674 240 6675 241 se
rect 6675 240 6748 241
tri 6748 240 6749 241 nw
tri 3653 212 3657 216 sw
rect 5730 212 5782 218
tri 6646 212 6674 240 se
rect 6674 212 6720 240
tri 6720 212 6748 240 nw
rect 7227 224 7236 241
rect 7270 224 7279 241
rect 3601 207 3657 212
tri 3657 207 3662 212 sw
tri 6641 207 6646 212 se
rect 6646 207 6715 212
tri 6715 207 6720 212 nw
rect 3601 195 3662 207
tri 3662 195 3674 207 sw
tri 6629 195 6641 207 se
rect 6641 195 6703 207
tri 6703 195 6715 207 nw
rect 3601 194 3674 195
tri 3601 188 3607 194 ne
rect 3607 188 3674 194
tri 3674 188 3681 195 sw
tri 6622 188 6629 195 se
rect 6629 188 6696 195
tri 6696 188 6703 195 nw
tri 3607 173 3622 188 ne
rect 3622 173 3681 188
tri 3681 173 3696 188 sw
tri 6607 173 6622 188 se
rect 6622 173 6674 188
tri 3622 166 3629 173 ne
rect 3629 166 6674 173
tri 6674 166 6696 188 nw
rect 7386 970 7392 1004
rect 7426 970 7432 1004
rect 7386 926 7432 970
rect 7386 892 7392 926
rect 7426 892 7432 926
rect 7386 848 7432 892
rect 7386 814 7392 848
rect 7426 814 7432 848
rect 7386 770 7432 814
rect 7386 736 7392 770
rect 7426 736 7432 770
rect 7386 692 7432 736
rect 7386 658 7392 692
rect 7426 658 7432 692
rect 7386 614 7432 658
rect 7386 580 7392 614
rect 7426 580 7432 614
rect 7386 536 7432 580
rect 7386 502 7392 536
rect 7426 502 7432 536
rect 7386 458 7432 502
rect 7386 424 7392 458
rect 7426 424 7432 458
rect 7386 380 7432 424
rect 7386 346 7392 380
rect 7426 346 7432 380
rect 7386 301 7432 346
rect 7386 267 7392 301
rect 7426 267 7432 301
rect 7386 222 7432 267
rect 7386 188 7392 222
rect 7426 188 7432 222
rect 7386 176 7432 188
rect 7493 1094 7545 1106
rect 7493 1060 7502 1094
rect 7536 1060 7545 1094
rect 7493 1019 7545 1060
rect 7925 1094 7977 1106
rect 7925 1060 7934 1094
rect 7968 1060 7977 1094
rect 7493 985 7502 1019
rect 7536 985 7545 1019
rect 7493 944 7545 985
rect 7493 910 7502 944
rect 7536 910 7545 944
rect 7493 869 7545 910
rect 7493 835 7502 869
rect 7536 835 7545 869
rect 7493 794 7545 835
rect 7493 760 7502 794
rect 7536 760 7545 794
rect 7493 736 7545 760
rect 7493 672 7545 684
rect 7493 610 7502 620
rect 7536 610 7545 620
rect 7493 569 7545 610
rect 7493 535 7502 569
rect 7536 535 7545 569
rect 7493 494 7545 535
rect 7493 460 7502 494
rect 7536 460 7545 494
rect 7493 419 7545 460
rect 7493 385 7502 419
rect 7536 385 7545 419
rect 7493 344 7545 385
rect 7493 310 7502 344
rect 7536 310 7545 344
rect 7493 269 7545 310
rect 7493 235 7502 269
rect 7536 235 7545 269
rect 7493 194 7545 235
rect 7227 166 7279 172
tri 3556 132 3590 166 sw
tri 3629 142 3653 166 ne
rect 3653 142 6640 166
tri 3653 132 3663 142 ne
rect 3663 132 6640 142
tri 6640 132 6674 166 nw
rect 7227 160 7236 166
rect 7270 160 7279 166
rect 7493 160 7502 194
rect 7536 160 7545 194
rect 7493 148 7545 160
rect 7709 1008 7761 1020
rect 7709 974 7718 1008
rect 7752 974 7761 1008
rect 7709 934 7761 974
rect 7709 900 7718 934
rect 7752 900 7761 934
rect 7709 892 7761 900
rect 7709 828 7718 840
rect 7752 828 7761 840
rect 7709 752 7718 776
rect 7752 752 7761 776
rect 7709 712 7761 752
rect 7709 678 7718 712
rect 7752 678 7761 712
rect 7709 638 7761 678
rect 7709 604 7718 638
rect 7752 604 7761 638
rect 7709 564 7761 604
rect 7709 530 7718 564
rect 7752 530 7761 564
rect 7709 490 7761 530
rect 7709 456 7718 490
rect 7752 456 7761 490
rect 7709 416 7761 456
rect 7709 382 7718 416
rect 7752 382 7761 416
rect 7709 342 7761 382
rect 7709 308 7718 342
rect 7752 308 7761 342
rect 7709 268 7761 308
rect 7709 234 7718 268
rect 7752 234 7761 268
rect 7709 194 7761 234
rect 7709 160 7718 194
rect 7752 160 7761 194
rect 7709 148 7761 160
rect 7925 1019 7977 1060
rect 7925 985 7934 1019
rect 7968 985 7977 1019
rect 7925 944 7977 985
rect 7925 910 7934 944
rect 7968 910 7977 944
rect 8180 1054 8322 1181
tri 9235 1146 9270 1181 se
rect 9270 1146 9322 2400
tri 9322 2388 9334 2400 nw
rect 9398 2388 9458 2394
rect 9398 2336 9402 2388
rect 9454 2336 9458 2388
rect 9398 2324 9458 2336
rect 9398 2272 9402 2324
rect 9454 2272 9458 2324
tri 9376 1230 9398 1252 se
rect 9398 1230 9458 2272
rect 9497 2371 9648 2400
rect 9682 2371 9688 2405
rect 9497 2362 9688 2371
rect 9497 2328 9503 2362
rect 9537 2332 9688 2362
rect 9537 2328 9648 2332
rect 9497 2298 9648 2328
rect 9682 2298 9688 2332
rect 9497 2290 9688 2298
rect 9497 2256 9503 2290
rect 9537 2259 9688 2290
rect 9537 2256 9648 2259
rect 9497 2225 9648 2256
rect 9682 2225 9688 2259
rect 9497 2218 9688 2225
rect 9497 2184 9503 2218
rect 9537 2186 9688 2218
rect 9537 2184 9648 2186
rect 9497 2152 9648 2184
rect 9682 2152 9688 2186
rect 9497 2146 9688 2152
rect 9497 2112 9503 2146
rect 9537 2113 9688 2146
rect 9537 2112 9648 2113
rect 9497 2079 9648 2112
rect 9682 2079 9688 2113
rect 9497 2074 9688 2079
rect 9497 2040 9503 2074
rect 9537 2040 9688 2074
rect 9497 2006 9648 2040
rect 9682 2006 9688 2040
rect 9497 2002 9688 2006
rect 9497 1968 9503 2002
rect 9537 1968 9688 2002
rect 9497 1967 9688 1968
rect 9497 1933 9648 1967
rect 9682 1933 9688 1967
rect 9497 1930 9688 1933
rect 9497 1896 9503 1930
rect 9537 1921 9688 1930
rect 9795 2782 9847 2794
rect 9795 2748 9803 2782
rect 9837 2748 9847 2782
rect 9795 2708 9847 2748
rect 9795 2674 9803 2708
rect 9837 2674 9847 2708
rect 9795 2634 9847 2674
rect 9795 2600 9803 2634
rect 9837 2600 9847 2634
rect 9795 2560 9847 2600
rect 9795 2526 9803 2560
rect 9837 2526 9847 2560
rect 9795 2486 9847 2526
rect 9795 2452 9803 2486
rect 9837 2452 9847 2486
rect 9795 2412 9847 2452
rect 9795 2388 9803 2412
rect 9837 2388 9847 2412
rect 9795 2324 9803 2336
rect 9837 2324 9847 2336
rect 9795 2264 9847 2272
rect 9795 2230 9803 2264
rect 9837 2230 9847 2264
rect 9795 2190 9847 2230
rect 9795 2156 9803 2190
rect 9837 2156 9847 2190
rect 9795 2116 9847 2156
rect 9795 2082 9803 2116
rect 9837 2082 9847 2116
rect 9795 2042 9847 2082
rect 9795 2008 9803 2042
rect 9837 2008 9847 2042
rect 9795 1967 9847 2008
rect 9795 1933 9803 1967
rect 9837 1933 9847 1967
rect 9795 1921 9847 1933
rect 9954 2765 10000 2803
rect 10266 2803 10272 2837
rect 10306 2803 10312 2837
tri 10312 2816 10333 2837 nw
tri 10557 2816 10578 2837 ne
rect 9954 2731 9960 2765
rect 9994 2731 10000 2765
rect 9954 2693 10000 2731
rect 9954 2659 9960 2693
rect 9994 2659 10000 2693
rect 9954 2621 10000 2659
rect 9954 2587 9960 2621
rect 9994 2587 10000 2621
rect 9954 2549 10000 2587
rect 9954 2515 9960 2549
rect 9994 2515 10000 2549
rect 9954 2477 10000 2515
rect 10110 2782 10156 2794
rect 10110 2748 10116 2782
rect 10150 2748 10156 2782
rect 10110 2705 10156 2748
rect 10110 2671 10116 2705
rect 10150 2671 10156 2705
rect 10110 2628 10156 2671
rect 10110 2594 10116 2628
rect 10150 2594 10156 2628
rect 10110 2551 10156 2594
rect 10110 2517 10116 2551
rect 10150 2517 10156 2551
tri 10108 2506 10110 2508 se
rect 10110 2506 10156 2517
rect 10266 2765 10312 2803
rect 10578 2803 10584 2837
rect 10618 2822 10630 2837
tri 10630 2822 10645 2837 nw
tri 10869 2822 10884 2837 ne
rect 10884 2822 10896 2837
rect 10618 2803 10624 2822
tri 10624 2816 10630 2822 nw
rect 10266 2731 10272 2765
rect 10306 2731 10312 2765
rect 10266 2693 10312 2731
rect 10266 2659 10272 2693
rect 10306 2659 10312 2693
rect 10266 2621 10312 2659
rect 10266 2587 10272 2621
rect 10306 2587 10312 2621
rect 10266 2549 10312 2587
rect 10266 2515 10272 2549
rect 10306 2515 10312 2549
tri 10156 2506 10158 2508 sw
tri 10104 2502 10108 2506 se
rect 10108 2502 10158 2506
tri 10158 2502 10162 2506 sw
tri 10093 2491 10104 2502 se
rect 10104 2491 10162 2502
tri 10162 2491 10173 2502 sw
tri 10079 2477 10093 2491 se
rect 10093 2477 10173 2491
tri 10173 2477 10187 2491 sw
rect 10266 2477 10312 2515
rect 9954 2443 9960 2477
rect 9994 2443 10000 2477
tri 10076 2474 10079 2477 se
rect 10079 2474 10187 2477
tri 10187 2474 10190 2477 sw
rect 9954 2405 10000 2443
rect 10068 2422 10074 2474
rect 10126 2422 10138 2440
rect 10190 2422 10196 2474
rect 10266 2443 10272 2477
rect 10306 2443 10312 2477
tri 10076 2411 10087 2422 ne
rect 10087 2411 10179 2422
tri 10179 2411 10190 2422 nw
tri 10087 2405 10093 2411 ne
rect 10093 2405 10173 2411
tri 10173 2405 10179 2411 nw
rect 10266 2405 10312 2443
rect 9954 2371 9960 2405
rect 9994 2371 10000 2405
tri 10093 2397 10101 2405 ne
rect 10101 2397 10156 2405
tri 10101 2388 10110 2397 ne
rect 9954 2332 10000 2371
rect 9954 2298 9960 2332
rect 9994 2298 10000 2332
rect 9954 2259 10000 2298
rect 9954 2225 9960 2259
rect 9994 2225 10000 2259
rect 9954 2186 10000 2225
rect 9954 2152 9960 2186
rect 9994 2152 10000 2186
rect 9954 2113 10000 2152
rect 9954 2079 9960 2113
rect 9994 2079 10000 2113
rect 9954 2040 10000 2079
rect 10110 2363 10116 2397
rect 10150 2363 10156 2397
tri 10156 2388 10173 2405 nw
rect 10110 2320 10156 2363
rect 10110 2286 10116 2320
rect 10150 2286 10156 2320
rect 10110 2243 10156 2286
rect 10110 2209 10116 2243
rect 10150 2209 10156 2243
rect 10110 2166 10156 2209
rect 10110 2132 10116 2166
rect 10150 2132 10156 2166
rect 10110 2088 10156 2132
rect 10110 2054 10116 2088
rect 10150 2054 10156 2088
rect 10110 2042 10156 2054
rect 10266 2371 10272 2405
rect 10306 2371 10312 2405
rect 10266 2332 10312 2371
rect 10266 2298 10272 2332
rect 10306 2298 10312 2332
rect 10266 2259 10312 2298
rect 10266 2225 10272 2259
rect 10306 2225 10312 2259
rect 10266 2186 10312 2225
rect 10266 2152 10272 2186
rect 10306 2152 10312 2186
rect 10266 2113 10312 2152
rect 10266 2079 10272 2113
rect 10306 2079 10312 2113
rect 9954 2006 9960 2040
rect 9994 2006 10000 2040
rect 9954 1967 10000 2006
rect 9954 1933 9960 1967
rect 9994 1933 10000 1967
rect 9954 1921 10000 1933
rect 10266 2040 10312 2079
rect 10419 2782 10471 2794
rect 10419 2748 10428 2782
rect 10462 2748 10471 2782
rect 10419 2705 10471 2748
rect 10419 2671 10428 2705
rect 10462 2671 10471 2705
rect 10419 2628 10471 2671
rect 10419 2594 10428 2628
rect 10462 2594 10471 2628
rect 10419 2551 10471 2594
rect 10419 2517 10428 2551
rect 10462 2517 10471 2551
rect 10419 2474 10471 2517
rect 10419 2440 10428 2474
rect 10462 2440 10471 2474
rect 10419 2397 10471 2440
rect 10419 2363 10428 2397
rect 10462 2363 10471 2397
rect 10419 2320 10471 2363
rect 10419 2286 10428 2320
rect 10462 2286 10471 2320
rect 10419 2243 10471 2286
rect 10419 2231 10428 2243
rect 10462 2231 10471 2243
rect 10419 2166 10471 2179
rect 10419 2088 10471 2114
rect 10419 2054 10428 2088
rect 10462 2054 10471 2088
rect 10419 2042 10471 2054
rect 10578 2765 10624 2803
rect 10578 2731 10584 2765
rect 10618 2731 10624 2765
rect 10578 2693 10624 2731
rect 10578 2659 10584 2693
rect 10618 2659 10624 2693
rect 10578 2621 10624 2659
rect 10578 2587 10584 2621
rect 10618 2587 10624 2621
rect 10578 2549 10624 2587
rect 10578 2515 10584 2549
rect 10618 2515 10624 2549
rect 10578 2477 10624 2515
rect 10578 2443 10584 2477
rect 10618 2443 10624 2477
rect 10578 2405 10624 2443
rect 10578 2371 10584 2405
rect 10618 2371 10624 2405
rect 10578 2332 10624 2371
rect 10578 2298 10584 2332
rect 10618 2298 10624 2332
rect 10578 2259 10624 2298
rect 10578 2225 10584 2259
rect 10618 2225 10624 2259
rect 10578 2186 10624 2225
rect 10578 2152 10584 2186
rect 10618 2152 10624 2186
rect 10578 2113 10624 2152
rect 10578 2079 10584 2113
rect 10618 2079 10624 2113
rect 10266 2006 10272 2040
rect 10306 2006 10312 2040
rect 10266 1967 10312 2006
rect 10266 1933 10272 1967
rect 10306 1933 10312 1967
rect 10266 1921 10312 1933
rect 10578 2040 10624 2079
rect 10731 2810 10783 2822
tri 10884 2816 10890 2822 ne
rect 10731 2776 10740 2810
rect 10774 2776 10783 2810
rect 10731 2731 10783 2776
rect 10731 2700 10740 2731
rect 10774 2700 10783 2731
rect 10731 2630 10740 2648
rect 10774 2630 10783 2648
rect 10731 2571 10783 2578
rect 10731 2560 10740 2571
rect 10774 2560 10783 2571
rect 10731 2491 10783 2508
rect 10731 2457 10740 2491
rect 10774 2457 10783 2491
rect 10731 2411 10783 2457
rect 10731 2377 10740 2411
rect 10774 2377 10783 2411
rect 10731 2331 10783 2377
rect 10731 2297 10740 2331
rect 10774 2297 10783 2331
rect 10731 2251 10783 2297
rect 10731 2217 10740 2251
rect 10774 2217 10783 2251
rect 10731 2171 10783 2217
rect 10731 2137 10740 2171
rect 10774 2137 10783 2171
rect 10731 2091 10783 2137
rect 10731 2057 10740 2091
rect 10774 2057 10783 2091
rect 10731 2045 10783 2057
rect 10890 2803 10896 2822
rect 10930 2822 10942 2837
tri 10942 2822 10957 2837 nw
tri 11181 2822 11196 2837 ne
rect 11196 2822 11208 2837
rect 10930 2803 10936 2822
tri 10936 2816 10942 2822 nw
rect 10890 2765 10936 2803
rect 10890 2731 10896 2765
rect 10930 2731 10936 2765
rect 10890 2693 10936 2731
rect 10890 2659 10896 2693
rect 10930 2659 10936 2693
rect 10890 2621 10936 2659
rect 10890 2587 10896 2621
rect 10930 2587 10936 2621
rect 10890 2549 10936 2587
rect 10890 2515 10896 2549
rect 10930 2515 10936 2549
rect 10890 2477 10936 2515
rect 10890 2443 10896 2477
rect 10930 2443 10936 2477
rect 10890 2405 10936 2443
rect 10890 2371 10896 2405
rect 10930 2371 10936 2405
rect 10890 2332 10936 2371
rect 10890 2298 10896 2332
rect 10930 2298 10936 2332
rect 10890 2259 10936 2298
rect 10890 2225 10896 2259
rect 10930 2225 10936 2259
rect 10890 2186 10936 2225
rect 10890 2152 10896 2186
rect 10930 2152 10936 2186
rect 10890 2113 10936 2152
rect 10890 2079 10896 2113
rect 10930 2079 10936 2113
rect 10578 2006 10584 2040
rect 10618 2006 10624 2040
rect 10578 1967 10624 2006
rect 10890 2040 10936 2079
rect 10890 2006 10896 2040
rect 10930 2006 10936 2040
rect 10578 1933 10584 1967
rect 10618 1933 10624 1967
rect 10578 1921 10624 1933
rect 10692 1948 10698 2000
rect 10750 1948 10762 2000
rect 10814 1948 10820 2000
rect 9537 1913 9569 1921
tri 9569 1913 9577 1921 nw
rect 9537 1898 9554 1913
tri 9554 1898 9569 1913 nw
tri 10677 1898 10692 1913 se
rect 10692 1898 10820 1948
rect 10890 1967 10936 2006
rect 10890 1933 10896 1967
rect 10930 1933 10936 1967
rect 10890 1921 10936 1933
rect 11043 2810 11095 2822
tri 11196 2816 11202 2822 ne
rect 11043 2776 11052 2810
rect 11086 2776 11095 2810
rect 11043 2734 11095 2776
rect 11043 2700 11052 2734
rect 11086 2700 11095 2734
rect 11043 2658 11095 2700
rect 11043 2624 11052 2658
rect 11086 2624 11095 2658
rect 11043 2582 11095 2624
rect 11043 2548 11052 2582
rect 11086 2548 11095 2582
rect 11043 2506 11095 2548
rect 11043 2472 11052 2506
rect 11086 2472 11095 2506
rect 11043 2429 11095 2472
rect 11043 2426 11052 2429
rect 11086 2426 11095 2429
rect 11043 2362 11095 2374
rect 11043 2275 11095 2310
rect 11043 2241 11052 2275
rect 11086 2241 11095 2275
rect 11043 2198 11095 2241
rect 11043 2164 11052 2198
rect 11086 2164 11095 2198
rect 11043 2121 11095 2164
rect 11043 2087 11052 2121
rect 11086 2087 11095 2121
rect 11043 2044 11095 2087
rect 11043 2010 11052 2044
rect 11086 2010 11095 2044
rect 11043 1967 11095 2010
rect 11043 1933 11052 1967
rect 11086 1933 11095 1967
rect 11043 1921 11095 1933
rect 11202 2803 11208 2822
rect 11242 2803 11248 2837
tri 11248 2816 11269 2837 nw
tri 11493 2816 11514 2837 ne
rect 11202 2765 11248 2803
rect 11514 2803 11520 2837
rect 11554 2803 11560 2837
tri 11560 2816 11582 2838 nw
tri 11667 2816 11689 2838 ne
rect 11202 2731 11208 2765
rect 11242 2731 11248 2765
rect 11310 2742 11316 2794
rect 11368 2782 11380 2794
rect 11368 2742 11380 2748
rect 11432 2742 11438 2794
tri 11324 2731 11335 2742 ne
rect 11335 2731 11427 2742
tri 11427 2731 11438 2742 nw
rect 11514 2765 11560 2803
rect 11514 2731 11520 2765
rect 11554 2731 11560 2765
rect 11202 2693 11248 2731
tri 11335 2728 11338 2731 ne
rect 11338 2728 11424 2731
tri 11424 2728 11427 2731 nw
tri 11338 2708 11358 2728 ne
rect 11358 2708 11404 2728
tri 11404 2708 11424 2728 nw
rect 11202 2659 11208 2693
rect 11242 2659 11248 2693
rect 11202 2621 11248 2659
rect 11202 2587 11208 2621
rect 11242 2587 11248 2621
rect 11202 2549 11248 2587
rect 11202 2515 11208 2549
rect 11242 2515 11248 2549
rect 11202 2477 11248 2515
rect 11202 2443 11208 2477
rect 11242 2443 11248 2477
rect 11202 2405 11248 2443
rect 11202 2371 11208 2405
rect 11242 2371 11248 2405
rect 11202 2332 11248 2371
rect 11202 2298 11208 2332
rect 11242 2298 11248 2332
rect 11202 2259 11248 2298
rect 11202 2225 11208 2259
rect 11242 2225 11248 2259
rect 11202 2186 11248 2225
rect 11202 2152 11208 2186
rect 11242 2152 11248 2186
rect 11202 2113 11248 2152
rect 11202 2079 11208 2113
rect 11242 2079 11248 2113
rect 11202 2040 11248 2079
rect 11202 2006 11208 2040
rect 11242 2006 11248 2040
rect 11202 1967 11248 2006
rect 11202 1933 11208 1967
rect 11242 1933 11248 1967
rect 11202 1921 11248 1933
rect 11358 2674 11364 2708
rect 11398 2674 11404 2708
rect 11358 2634 11404 2674
rect 11358 2600 11364 2634
rect 11398 2600 11404 2634
rect 11358 2560 11404 2600
rect 11358 2526 11364 2560
rect 11398 2526 11404 2560
rect 11358 2486 11404 2526
rect 11358 2452 11364 2486
rect 11398 2452 11404 2486
rect 11358 2412 11404 2452
rect 11358 2378 11364 2412
rect 11398 2378 11404 2412
rect 11358 2338 11404 2378
rect 11358 2304 11364 2338
rect 11398 2304 11404 2338
rect 11358 2264 11404 2304
rect 11358 2230 11364 2264
rect 11398 2230 11404 2264
rect 11358 2190 11404 2230
rect 11358 2156 11364 2190
rect 11398 2156 11404 2190
rect 11358 2116 11404 2156
rect 11358 2082 11364 2116
rect 11398 2082 11404 2116
rect 11358 2042 11404 2082
rect 11358 2008 11364 2042
rect 11398 2008 11404 2042
rect 11358 1967 11404 2008
rect 11358 1933 11364 1967
rect 11398 1933 11404 1967
rect 11358 1921 11404 1933
rect 11514 2693 11560 2731
rect 11514 2659 11520 2693
rect 11554 2659 11560 2693
rect 11514 2621 11560 2659
rect 11514 2587 11520 2621
rect 11554 2587 11560 2621
rect 11514 2549 11560 2587
rect 11514 2515 11520 2549
rect 11554 2515 11560 2549
rect 11514 2477 11560 2515
rect 11514 2443 11520 2477
rect 11554 2443 11560 2477
rect 11514 2405 11560 2443
rect 11514 2371 11520 2405
rect 11554 2371 11560 2405
rect 11514 2332 11560 2371
rect 11514 2298 11520 2332
rect 11554 2298 11560 2332
rect 11514 2259 11560 2298
rect 11514 2225 11520 2259
rect 11554 2225 11560 2259
rect 11514 2186 11560 2225
rect 11514 2152 11520 2186
rect 11554 2152 11560 2186
rect 11514 2113 11560 2152
rect 11514 2079 11520 2113
rect 11554 2079 11560 2113
rect 11514 2040 11560 2079
rect 11514 2006 11520 2040
rect 11554 2006 11560 2040
rect 11514 1967 11560 2006
rect 11514 1933 11520 1967
rect 11554 1933 11560 1967
rect 11514 1921 11560 1933
rect 11689 2800 11735 2838
rect 11689 2766 11695 2800
rect 11729 2766 11735 2800
rect 11689 2728 11735 2766
rect 11689 2694 11695 2728
rect 11729 2694 11735 2728
rect 11689 2656 11735 2694
rect 11689 2622 11695 2656
rect 11729 2622 11735 2656
rect 11689 2584 11735 2622
rect 11689 2550 11695 2584
rect 11729 2550 11735 2584
rect 11689 2512 11735 2550
rect 11689 2478 11695 2512
rect 11729 2478 11735 2512
rect 11689 2440 11735 2478
rect 11689 2406 11695 2440
rect 11729 2406 11735 2440
rect 11689 2368 11735 2406
rect 11689 2334 11695 2368
rect 11729 2334 11735 2368
rect 11689 2296 11735 2334
rect 11689 2262 11695 2296
rect 11729 2262 11735 2296
rect 11689 2224 11735 2262
rect 11689 2190 11695 2224
rect 11729 2190 11735 2224
rect 11689 2151 11735 2190
rect 11689 2117 11695 2151
rect 11729 2117 11735 2151
rect 11689 2078 11735 2117
rect 11689 2044 11695 2078
rect 11729 2044 11735 2078
rect 11689 2005 11735 2044
rect 11689 1971 11695 2005
rect 11729 1971 11735 2005
rect 11689 1932 11735 1971
tri 10820 1898 10835 1913 sw
rect 11689 1898 11695 1932
rect 11729 1898 11735 1932
rect 9537 1896 9543 1898
rect 9497 1858 9543 1896
tri 9543 1887 9554 1898 nw
tri 10666 1887 10677 1898 se
rect 10677 1887 10835 1898
tri 10658 1879 10666 1887 se
rect 10666 1882 10835 1887
tri 10835 1882 10851 1898 sw
rect 10666 1879 10851 1882
tri 10851 1879 10854 1882 sw
rect 9497 1824 9503 1858
rect 9537 1824 9543 1858
rect 9497 1786 9543 1824
rect 9497 1752 9503 1786
rect 9537 1752 9543 1786
rect 9699 1873 9927 1879
rect 9699 1839 9711 1873
rect 9745 1839 9796 1873
rect 9830 1839 9881 1873
rect 9915 1839 9927 1873
rect 9699 1833 9927 1839
rect 10274 1873 10858 1879
rect 10274 1839 10286 1873
rect 10320 1839 10362 1873
rect 10396 1839 10437 1873
rect 10471 1839 10512 1873
rect 10546 1839 10587 1873
rect 10621 1839 10662 1873
rect 10696 1839 10737 1873
rect 10771 1839 10812 1873
rect 10846 1839 10858 1873
rect 10274 1833 10858 1839
rect 9699 1830 9782 1833
tri 9782 1830 9785 1833 nw
rect 10942 1830 10948 1882
rect 11000 1830 11012 1882
rect 11064 1873 11503 1882
rect 11081 1839 11140 1873
rect 11174 1839 11271 1873
rect 11305 1839 11364 1873
rect 11398 1839 11457 1873
rect 11491 1839 11503 1873
rect 11064 1830 11503 1839
rect 11689 1859 11735 1898
rect 9699 1825 9777 1830
tri 9777 1825 9782 1830 nw
rect 11689 1825 11695 1859
rect 11729 1825 11735 1859
tri 9543 1752 9545 1754 sw
rect 9497 1722 9545 1752
tri 9545 1722 9575 1752 sw
rect 9497 1720 9575 1722
tri 9575 1720 9577 1722 sw
rect 9497 1714 9604 1720
rect 9497 1680 9517 1714
rect 9551 1680 9604 1714
rect 9497 1674 9604 1680
tri 9691 1650 9699 1658 se
rect 9699 1650 9751 1825
tri 9751 1799 9777 1825 nw
rect 11689 1786 11735 1825
tri 11687 1752 11689 1754 se
rect 11689 1752 11695 1786
rect 11729 1752 11735 1786
tri 11657 1722 11687 1752 se
rect 11687 1722 11735 1752
tri 11655 1720 11657 1722 se
rect 11657 1720 11735 1722
rect 10240 1714 11735 1720
rect 10240 1680 10278 1714
rect 10312 1680 10353 1714
rect 10387 1680 10428 1714
rect 10462 1680 10503 1714
rect 10537 1680 10578 1714
rect 10612 1680 10653 1714
rect 10687 1680 10728 1714
rect 10762 1680 10803 1714
rect 10837 1680 10878 1714
rect 10912 1680 10953 1714
rect 10987 1680 11028 1714
rect 11062 1680 11103 1714
rect 11137 1680 11177 1714
rect 11211 1680 11251 1714
rect 11285 1680 11325 1714
rect 11359 1680 11399 1714
rect 11433 1680 11473 1714
rect 11507 1680 11547 1714
rect 11581 1680 11621 1714
rect 11655 1680 11735 1714
rect 10240 1674 11735 1680
rect 11916 3297 17128 3298
rect 11916 3245 11922 3297
rect 11974 3245 11987 3297
rect 12039 3245 12052 3297
rect 12104 3245 12117 3297
rect 12169 3245 12182 3297
rect 12234 3245 12247 3297
rect 12299 3245 12312 3297
rect 12364 3245 12377 3297
rect 12429 3245 12442 3297
rect 12494 3245 12507 3297
rect 12559 3245 12572 3297
rect 12624 3245 12637 3297
rect 12689 3245 12702 3297
rect 12754 3245 12767 3297
rect 12819 3245 12832 3297
rect 12884 3245 12897 3297
rect 12949 3245 12962 3297
rect 13014 3245 13027 3297
rect 13079 3245 13092 3297
rect 13144 3245 13157 3297
rect 13209 3245 13222 3297
rect 13274 3245 13287 3297
rect 13339 3245 13352 3297
rect 13404 3245 13417 3297
rect 13469 3245 13482 3297
rect 13534 3245 13547 3297
rect 13599 3245 13612 3297
rect 13664 3245 13677 3297
rect 13729 3245 13742 3297
rect 13794 3245 13806 3297
rect 13858 3245 13870 3297
rect 13922 3245 13934 3297
rect 13986 3245 13998 3297
rect 14050 3245 14062 3297
rect 14114 3245 14126 3297
rect 14178 3245 14190 3297
rect 14242 3245 14254 3297
rect 14306 3245 14318 3297
rect 14370 3245 14382 3297
rect 14434 3245 14446 3297
rect 14498 3245 14510 3297
rect 14562 3245 14574 3297
rect 14626 3245 14638 3297
rect 14690 3245 14702 3297
rect 14754 3245 14766 3297
rect 14818 3245 14830 3297
rect 14882 3245 14894 3297
rect 14946 3245 14958 3297
rect 15010 3245 15022 3297
rect 15074 3245 15086 3297
rect 15138 3245 15150 3297
rect 15202 3245 15214 3297
rect 15266 3245 15278 3297
rect 15330 3245 15342 3297
rect 15394 3245 15406 3297
rect 15458 3245 15470 3297
rect 15522 3245 15534 3297
rect 15586 3245 15598 3297
rect 15650 3245 15662 3297
rect 15714 3245 15726 3297
rect 15778 3245 15790 3297
rect 15842 3245 15854 3297
rect 15906 3245 15918 3297
rect 15970 3245 15982 3297
rect 16034 3245 16046 3297
rect 16098 3245 16110 3297
rect 16162 3245 16174 3297
rect 16226 3245 16238 3297
rect 16290 3245 16302 3297
rect 16354 3245 16366 3297
rect 16418 3245 16430 3297
rect 16482 3245 16494 3297
rect 16546 3245 16558 3297
rect 16610 3245 16622 3297
rect 16674 3245 16686 3297
rect 16738 3245 16750 3297
rect 16802 3245 16814 3297
rect 16866 3245 16878 3297
rect 16930 3245 16942 3297
rect 16994 3245 17006 3297
rect 17058 3245 17070 3297
rect 17122 3245 17128 3297
rect 11916 3187 17128 3245
rect 11916 3135 11922 3187
rect 11974 3135 11987 3187
rect 12039 3135 12052 3187
rect 12104 3135 12117 3187
rect 12169 3135 12182 3187
rect 12234 3135 12247 3187
rect 12299 3135 12312 3187
rect 12364 3135 12377 3187
rect 12429 3135 12442 3187
rect 12494 3135 12507 3187
rect 12559 3135 12572 3187
rect 12624 3135 12637 3187
rect 12689 3135 12702 3187
rect 12754 3135 12767 3187
rect 12819 3135 12832 3187
rect 12884 3135 12897 3187
rect 12949 3135 12962 3187
rect 13014 3135 13027 3187
rect 13079 3135 13092 3187
rect 13144 3135 13157 3187
rect 13209 3135 13222 3187
rect 13274 3135 13287 3187
rect 13339 3135 13352 3187
rect 13404 3135 13417 3187
rect 13469 3135 13482 3187
rect 13534 3135 13547 3187
rect 13599 3135 13612 3187
rect 13664 3135 13677 3187
rect 13729 3135 13742 3187
rect 13794 3135 13806 3187
rect 13858 3135 13870 3187
rect 13922 3135 13934 3187
rect 13986 3135 13998 3187
rect 14050 3135 14062 3187
rect 14114 3135 14126 3187
rect 14178 3135 14190 3187
rect 14242 3135 14254 3187
rect 14306 3135 14318 3187
rect 14370 3135 14382 3187
rect 14434 3135 14446 3187
rect 14498 3135 14510 3187
rect 14562 3135 14574 3187
rect 14626 3135 14638 3187
rect 14690 3135 14702 3187
rect 14754 3135 14766 3187
rect 14818 3135 14830 3187
rect 14882 3135 14894 3187
rect 14946 3135 14958 3187
rect 15010 3135 15022 3187
rect 15074 3135 15086 3187
rect 15138 3135 15150 3187
rect 15202 3135 15214 3187
rect 15266 3135 15278 3187
rect 15330 3135 15342 3187
rect 15394 3135 15406 3187
rect 15458 3135 15470 3187
rect 15522 3135 15534 3187
rect 15586 3135 15598 3187
rect 15650 3135 15662 3187
rect 15714 3135 15726 3187
rect 15778 3135 15790 3187
rect 15842 3135 15854 3187
rect 15906 3135 15918 3187
rect 15970 3135 15982 3187
rect 16034 3135 16046 3187
rect 16098 3135 16110 3187
rect 16162 3135 16174 3187
rect 16226 3135 16238 3187
rect 16290 3135 16302 3187
rect 16354 3135 16366 3187
rect 16418 3135 16430 3187
rect 16482 3135 16494 3187
rect 16546 3135 16558 3187
rect 16610 3135 16622 3187
rect 16674 3135 16686 3187
rect 16738 3135 16750 3187
rect 16802 3135 16814 3187
rect 16866 3135 16878 3187
rect 16930 3135 16942 3187
rect 16994 3135 17006 3187
rect 17058 3135 17070 3187
rect 17122 3135 17128 3187
rect 11916 3064 17128 3135
rect 11916 3030 11994 3064
rect 12028 3030 12066 3064
rect 12100 3030 12138 3064
rect 12172 3030 12210 3064
rect 12244 3030 12282 3064
rect 12316 3030 12354 3064
rect 12388 3030 12426 3064
rect 12460 3030 12498 3064
rect 12532 3030 12570 3064
rect 12604 3030 12642 3064
rect 12676 3030 12714 3064
rect 12748 3030 12786 3064
rect 12820 3030 12858 3064
rect 12892 3030 12930 3064
rect 12964 3030 13002 3064
rect 13036 3030 13074 3064
rect 13108 3030 13146 3064
rect 13180 3030 13218 3064
rect 13252 3030 13290 3064
rect 13324 3030 13362 3064
rect 13396 3030 13434 3064
rect 13468 3030 13506 3064
rect 13540 3030 13578 3064
rect 13612 3030 13650 3064
rect 13684 3030 13722 3064
rect 13756 3030 13794 3064
rect 13828 3030 13866 3064
rect 13900 3030 13938 3064
rect 13972 3030 14010 3064
rect 14044 3030 14082 3064
rect 14116 3030 14154 3064
rect 14188 3030 14226 3064
rect 14260 3030 14298 3064
rect 14332 3030 14370 3064
rect 14404 3030 14442 3064
rect 14476 3030 14514 3064
rect 14548 3030 14586 3064
rect 14620 3030 14658 3064
rect 14692 3030 14730 3064
rect 14764 3030 14802 3064
rect 14836 3030 14874 3064
rect 14908 3030 14946 3064
rect 14980 3030 15018 3064
rect 15052 3030 15090 3064
rect 15124 3030 15162 3064
rect 15196 3030 15234 3064
rect 15268 3030 15306 3064
rect 15340 3030 15378 3064
rect 15412 3030 15450 3064
rect 15484 3030 15522 3064
rect 15556 3030 15594 3064
rect 15628 3030 15666 3064
rect 15700 3030 15738 3064
rect 15772 3030 15810 3064
rect 15844 3030 15882 3064
rect 15916 3030 15954 3064
rect 15988 3030 16026 3064
rect 16060 3030 16098 3064
rect 16132 3030 16170 3064
rect 16204 3030 16243 3064
rect 16277 3030 16316 3064
rect 16350 3030 16389 3064
rect 16423 3030 16462 3064
rect 16496 3030 16572 3064
rect 16606 3030 16646 3064
rect 16680 3030 16720 3064
rect 16754 3030 16794 3064
rect 16828 3030 16868 3064
rect 16902 3030 16942 3064
rect 16976 3030 17016 3064
rect 17050 3030 17128 3064
rect 11916 3024 17128 3030
rect 11916 2992 11964 3024
tri 11964 2992 11996 3024 nw
tri 14495 2992 14527 3024 ne
rect 14527 2992 14577 3024
tri 14577 2992 14609 3024 nw
tri 17048 2992 17080 3024 ne
rect 17080 2992 17128 3024
rect 11916 2958 11922 2992
rect 11956 2958 11962 2992
tri 11962 2990 11964 2992 nw
tri 14527 2990 14529 2992 ne
rect 11916 2919 11962 2958
rect 11916 2885 11922 2919
rect 11956 2885 11962 2919
rect 11916 2846 11962 2885
rect 11916 2812 11922 2846
rect 11956 2812 11962 2846
rect 11916 2773 11962 2812
rect 14529 2961 14575 2992
tri 14575 2990 14577 2992 nw
tri 17080 2990 17082 2992 ne
rect 14529 2927 14535 2961
rect 14569 2927 14575 2961
rect 14529 2887 14575 2927
rect 16837 2982 16965 2988
rect 16889 2930 16913 2982
rect 14529 2853 14535 2887
rect 14569 2853 14575 2887
rect 14529 2813 14575 2853
rect 11916 2739 11922 2773
rect 11956 2739 11962 2773
rect 11916 2700 11962 2739
rect 11916 2666 11922 2700
rect 11956 2666 11962 2700
rect 11916 2627 11962 2666
rect 11916 2593 11922 2627
rect 11956 2593 11962 2627
rect 12196 2778 14222 2784
rect 12196 2744 12208 2778
rect 12242 2744 12281 2778
rect 12315 2744 12354 2778
rect 12388 2744 12427 2778
rect 12461 2744 12500 2778
rect 12534 2744 12573 2778
rect 12607 2744 12646 2778
rect 12680 2744 12719 2778
rect 12753 2744 12792 2778
rect 12826 2744 12865 2778
rect 12899 2744 12938 2778
rect 12972 2744 13011 2778
rect 13045 2744 13084 2778
rect 13118 2744 13157 2778
rect 13191 2744 13230 2778
rect 13264 2744 13303 2778
rect 13337 2744 13376 2778
rect 13410 2744 13449 2778
rect 13483 2744 13522 2778
rect 13556 2744 13595 2778
rect 13629 2744 13668 2778
rect 13702 2744 13741 2778
rect 13775 2744 13814 2778
rect 13848 2744 13887 2778
rect 13921 2744 13960 2778
rect 13994 2744 14032 2778
rect 14066 2744 14104 2778
rect 14138 2744 14176 2778
rect 14210 2744 14222 2778
rect 12196 2660 14222 2744
rect 12196 2626 12252 2660
rect 12286 2626 12326 2660
rect 12360 2626 12400 2660
rect 12434 2626 12474 2660
rect 12508 2626 12548 2660
rect 12582 2626 12622 2660
rect 12656 2626 12696 2660
rect 12730 2626 12770 2660
rect 12804 2626 12844 2660
rect 12878 2626 12918 2660
rect 12952 2626 12992 2660
rect 13026 2626 13066 2660
rect 13100 2626 13140 2660
rect 13174 2626 13214 2660
rect 13248 2626 13288 2660
rect 13322 2626 13362 2660
rect 13396 2626 13436 2660
rect 13470 2626 13510 2660
rect 13544 2626 13584 2660
rect 13618 2626 13658 2660
rect 13692 2626 13732 2660
rect 13766 2626 13806 2660
rect 13840 2626 13880 2660
rect 13914 2626 13954 2660
rect 13988 2626 14028 2660
rect 14062 2626 14102 2660
rect 14136 2626 14176 2660
rect 14210 2626 14222 2660
rect 12196 2620 14222 2626
tri 14000 2598 14022 2620 ne
rect 14022 2598 14222 2620
rect 14529 2779 14535 2813
rect 14569 2779 14575 2813
rect 14529 2739 14575 2779
rect 14529 2705 14535 2739
rect 14569 2705 14575 2739
rect 14529 2665 14575 2705
rect 14529 2631 14535 2665
rect 14569 2631 14575 2665
rect 11916 2554 11962 2593
tri 14022 2591 14029 2598 ne
rect 14029 2591 14222 2598
tri 14029 2588 14032 2591 ne
rect 14032 2588 14222 2591
tri 14032 2586 14034 2588 ne
rect 11916 2520 11922 2554
rect 11956 2520 11962 2554
rect 11916 2481 11962 2520
rect 11916 2447 11922 2481
rect 11956 2447 11962 2481
rect 11916 2408 11962 2447
rect 11916 2374 11922 2408
rect 11956 2374 11962 2408
rect 11916 2335 11962 2374
rect 11916 2301 11922 2335
rect 11956 2301 11962 2335
rect 11916 2262 11962 2301
rect 11916 2228 11922 2262
rect 11956 2228 11962 2262
rect 11916 2189 11962 2228
rect 11916 2155 11922 2189
rect 11956 2155 11962 2189
rect 11916 2116 11962 2155
rect 11916 2082 11922 2116
rect 11956 2082 11962 2116
rect 11916 2044 11962 2082
rect 11916 2010 11922 2044
rect 11956 2010 11962 2044
rect 11916 1972 11962 2010
rect 11916 1938 11922 1972
rect 11956 1938 11962 1972
rect 11916 1900 11962 1938
rect 12219 2378 12225 2430
rect 12277 2424 12301 2430
rect 12353 2424 13966 2430
rect 12286 2390 12301 2424
rect 12359 2390 12398 2424
rect 12432 2390 12471 2424
rect 12505 2390 12544 2424
rect 12578 2390 12617 2424
rect 12651 2390 12690 2424
rect 12724 2390 12763 2424
rect 12797 2390 12836 2424
rect 12870 2390 12909 2424
rect 12943 2390 12982 2424
rect 13016 2390 13055 2424
rect 13089 2390 13128 2424
rect 13162 2390 13200 2424
rect 13234 2390 13272 2424
rect 13306 2390 13344 2424
rect 13378 2390 13416 2424
rect 13450 2390 13488 2424
rect 13522 2390 13560 2424
rect 13594 2390 13632 2424
rect 13666 2390 13704 2424
rect 13738 2390 13776 2424
rect 13810 2390 13848 2424
rect 13882 2390 13920 2424
rect 13954 2390 13966 2424
rect 12277 2378 12301 2390
rect 12353 2384 13966 2390
rect 12353 2379 12388 2384
tri 12388 2379 12393 2384 nw
rect 12353 2378 12378 2379
rect 12219 2369 12378 2378
tri 12378 2369 12388 2379 nw
rect 12219 2356 12359 2369
rect 12219 2304 12225 2356
rect 12277 2304 12301 2356
rect 12353 2304 12359 2356
tri 12359 2350 12378 2369 nw
rect 12219 1988 12359 2304
rect 14034 2236 14222 2588
tri 14027 2221 14034 2228 se
rect 14034 2221 14040 2236
tri 14000 2194 14027 2221 se
rect 14027 2194 14040 2221
rect 12408 2188 14040 2194
rect 14092 2188 14164 2236
rect 12408 2154 12420 2188
rect 12454 2154 12494 2188
rect 12528 2154 12568 2188
rect 12602 2154 12642 2188
rect 12676 2154 12716 2188
rect 12750 2154 12789 2188
rect 12823 2154 12862 2188
rect 12896 2154 12935 2188
rect 12969 2154 13008 2188
rect 13042 2154 13081 2188
rect 13115 2154 13154 2188
rect 13188 2154 13227 2188
rect 13261 2154 13300 2188
rect 13334 2154 13373 2188
rect 13407 2154 13446 2188
rect 13480 2154 13519 2188
rect 13553 2154 13592 2188
rect 13626 2154 13665 2188
rect 13699 2154 13738 2188
rect 13772 2154 13811 2188
rect 13845 2154 13884 2188
rect 13918 2154 13957 2188
rect 13991 2154 14030 2188
rect 14092 2184 14103 2188
rect 14064 2160 14103 2184
rect 14092 2154 14103 2160
rect 14137 2184 14164 2188
rect 14216 2184 14222 2236
rect 14137 2160 14176 2184
rect 14210 2160 14222 2184
rect 14137 2154 14164 2160
rect 12408 2148 14040 2154
tri 14000 2147 14001 2148 ne
rect 14001 2147 14040 2148
tri 14001 2114 14034 2147 ne
rect 14034 2108 14040 2147
rect 14092 2108 14164 2154
rect 14216 2108 14222 2160
tri 12359 1988 12363 1992 sw
rect 12219 1964 12363 1988
tri 12363 1964 12387 1988 sw
rect 12219 1958 12387 1964
tri 12387 1958 12393 1964 sw
rect 12219 1952 13966 1958
rect 12219 1918 12252 1952
rect 12286 1918 12325 1952
rect 12359 1918 12398 1952
rect 12432 1918 12471 1952
rect 12505 1918 12544 1952
rect 12578 1918 12617 1952
rect 12651 1918 12690 1952
rect 12724 1918 12763 1952
rect 12797 1918 12836 1952
rect 12870 1918 12909 1952
rect 12943 1918 12982 1952
rect 13016 1918 13055 1952
rect 13089 1918 13128 1952
rect 13162 1918 13200 1952
rect 13234 1918 13272 1952
rect 13306 1918 13344 1952
rect 13378 1918 13416 1952
rect 13450 1918 13488 1952
rect 13522 1918 13560 1952
rect 13594 1918 13632 1952
rect 13666 1918 13704 1952
rect 13738 1918 13776 1952
rect 13810 1918 13848 1952
rect 13882 1918 13920 1952
rect 13954 1918 13966 1952
rect 14034 1921 14222 2108
rect 14260 2588 14313 2600
rect 14260 2554 14266 2588
rect 14300 2554 14313 2588
rect 14260 2508 14313 2554
rect 14260 2474 14266 2508
rect 14300 2474 14313 2508
rect 14260 2427 14313 2474
rect 14260 2393 14266 2427
rect 14300 2393 14313 2427
rect 14260 2346 14313 2393
rect 14312 2294 14313 2346
rect 14260 2282 14313 2294
rect 14312 2230 14313 2282
rect 14260 2184 14313 2230
rect 14260 2150 14266 2184
rect 14300 2150 14313 2184
rect 14260 2103 14313 2150
rect 14260 2069 14266 2103
rect 14300 2069 14313 2103
rect 14260 2022 14313 2069
rect 14260 1988 14266 2022
rect 14300 1988 14313 2022
rect 14260 1976 14313 1988
rect 14529 2591 14575 2631
rect 14884 2893 15024 2899
rect 14936 2841 14972 2893
rect 14884 2825 15024 2841
rect 14936 2778 14972 2825
rect 16837 2890 16965 2930
rect 16889 2838 16913 2890
tri 15024 2814 15028 2818 sw
rect 15024 2784 15028 2814
tri 15028 2784 15058 2814 sw
rect 15024 2778 16791 2784
rect 14936 2773 14970 2778
rect 15024 2773 15044 2778
rect 14884 2757 14896 2773
rect 14930 2757 14970 2773
rect 15004 2757 15044 2773
rect 14936 2744 14970 2757
rect 15024 2744 15044 2757
rect 15078 2744 15118 2778
rect 15152 2744 15192 2778
rect 15226 2744 15266 2778
rect 15300 2744 15340 2778
rect 15374 2744 15414 2778
rect 15448 2744 15488 2778
rect 15522 2744 15562 2778
rect 15596 2744 15636 2778
rect 15670 2744 15710 2778
rect 15744 2744 15784 2778
rect 15818 2744 15858 2778
rect 15892 2744 15932 2778
rect 15966 2744 16006 2778
rect 16040 2744 16080 2778
rect 16114 2744 16154 2778
rect 16188 2744 16228 2778
rect 16262 2744 16302 2778
rect 16336 2744 16376 2778
rect 16410 2744 16450 2778
rect 16484 2744 16524 2778
rect 16558 2744 16598 2778
rect 16632 2744 16672 2778
rect 16706 2744 16745 2778
rect 16779 2744 16791 2778
rect 14936 2705 14972 2744
rect 15024 2738 16791 2744
rect 14529 2557 14535 2591
rect 14569 2557 14575 2591
rect 14529 2517 14575 2557
rect 14529 2483 14535 2517
rect 14569 2483 14575 2517
rect 14529 2443 14575 2483
rect 14529 2409 14535 2443
rect 14569 2409 14575 2443
rect 14529 2369 14575 2409
rect 14529 2335 14535 2369
rect 14569 2335 14575 2369
rect 14529 2295 14575 2335
rect 14529 2261 14535 2295
rect 14569 2261 14575 2295
rect 14529 2221 14575 2261
rect 14529 2187 14535 2221
rect 14569 2187 14575 2221
rect 14529 2147 14575 2187
rect 14529 2113 14535 2147
rect 14569 2113 14575 2147
rect 14529 2073 14575 2113
rect 14529 2039 14535 2073
rect 14569 2039 14575 2073
rect 14529 1998 14575 2039
rect 14529 1964 14535 1998
rect 14569 1964 14575 1998
rect 14767 2588 14820 2600
rect 14767 2554 14780 2588
rect 14814 2554 14820 2588
rect 14767 2508 14820 2554
rect 14767 2474 14780 2508
rect 14814 2474 14820 2508
rect 14767 2427 14820 2474
rect 14767 2393 14780 2427
rect 14814 2393 14820 2427
rect 14767 2346 14820 2393
rect 14819 2294 14820 2346
rect 14767 2282 14820 2294
rect 14819 2230 14820 2282
rect 14767 2184 14820 2230
rect 14767 2150 14780 2184
rect 14814 2150 14820 2184
rect 14767 2103 14820 2150
rect 14767 2069 14780 2103
rect 14814 2069 14820 2103
rect 14767 2022 14820 2069
rect 14767 1988 14780 2022
rect 14814 1988 14820 2022
rect 14767 1976 14820 1988
rect 14884 2452 15024 2705
tri 15024 2704 15058 2738 nw
tri 16807 2670 16837 2700 se
rect 16837 2670 16965 2838
tri 16803 2666 16807 2670 se
rect 16807 2666 16965 2670
rect 15133 2660 16965 2666
rect 15133 2626 15145 2660
rect 15179 2626 15218 2660
rect 15252 2626 15291 2660
rect 15325 2626 15364 2660
rect 15398 2626 15437 2660
rect 15471 2626 15510 2660
rect 15544 2626 15583 2660
rect 15617 2626 15656 2660
rect 15690 2626 15729 2660
rect 15763 2626 15802 2660
rect 15836 2626 15875 2660
rect 15909 2626 15948 2660
rect 15982 2626 16021 2660
rect 16055 2626 16094 2660
rect 16128 2626 16167 2660
rect 16201 2626 16240 2660
rect 16274 2626 16313 2660
rect 16347 2626 16386 2660
rect 16420 2626 16459 2660
rect 16493 2626 16532 2660
rect 16566 2626 16604 2660
rect 16638 2626 16676 2660
rect 16710 2626 16748 2660
rect 16782 2626 16820 2660
rect 16854 2626 16965 2660
rect 15133 2620 16965 2626
tri 16803 2598 16825 2620 ne
rect 16825 2598 16965 2620
tri 16825 2586 16837 2598 ne
tri 15024 2452 15036 2464 sw
rect 14884 2430 15036 2452
tri 15036 2430 15058 2452 sw
rect 14884 2424 16650 2430
rect 14884 2390 14896 2424
rect 14930 2390 14971 2424
rect 15005 2390 15046 2424
rect 15080 2390 15121 2424
rect 15155 2390 15196 2424
rect 15230 2390 15271 2424
rect 15305 2390 15346 2424
rect 15380 2390 15420 2424
rect 15454 2390 15494 2424
rect 15528 2390 15568 2424
rect 15602 2390 15642 2424
rect 15676 2390 15716 2424
rect 15750 2390 15790 2424
rect 15824 2390 15864 2424
rect 15898 2390 15938 2424
rect 15972 2390 16012 2424
rect 16046 2390 16086 2424
rect 16120 2390 16160 2424
rect 16194 2390 16234 2424
rect 16268 2390 16308 2424
rect 16342 2390 16382 2424
rect 16416 2390 16456 2424
rect 16490 2390 16530 2424
rect 16564 2390 16604 2424
rect 16638 2390 16650 2424
rect 14884 2384 16650 2390
rect 14884 2379 15053 2384
tri 15053 2379 15058 2384 nw
rect 14529 1923 14575 1964
rect 12219 1912 13966 1918
rect 11916 1866 11922 1900
rect 11956 1866 11962 1900
rect 11916 1828 11962 1866
rect 11916 1794 11922 1828
rect 11956 1794 11962 1828
rect 11916 1756 11962 1794
rect 11916 1722 11922 1756
rect 11956 1722 11962 1756
rect 14529 1889 14535 1923
rect 14569 1889 14575 1923
rect 14884 1975 15024 2379
tri 15024 2350 15053 2379 nw
tri 16803 2194 16837 2228 se
rect 16837 2194 16965 2598
rect 15052 2188 16965 2194
rect 15052 2154 15064 2188
rect 15098 2154 15138 2188
rect 15172 2154 15212 2188
rect 15246 2154 15286 2188
rect 15320 2154 15360 2188
rect 15394 2154 15433 2188
rect 15467 2154 15506 2188
rect 15540 2154 15579 2188
rect 15613 2154 15652 2188
rect 15686 2154 15725 2188
rect 15759 2154 15798 2188
rect 15832 2154 15871 2188
rect 15905 2154 15944 2188
rect 15978 2154 16017 2188
rect 16051 2154 16090 2188
rect 16124 2154 16163 2188
rect 16197 2154 16236 2188
rect 16270 2154 16309 2188
rect 16343 2154 16382 2188
rect 16416 2154 16455 2188
rect 16489 2154 16528 2188
rect 16562 2154 16601 2188
rect 16635 2154 16674 2188
rect 16708 2154 16747 2188
rect 16781 2154 16820 2188
rect 16854 2154 16965 2188
rect 15052 2148 16965 2154
rect 17082 2958 17088 2992
rect 17122 2958 17128 2992
rect 17082 2920 17128 2958
rect 17082 2886 17088 2920
rect 17122 2886 17128 2920
rect 17082 2848 17128 2886
rect 17082 2814 17088 2848
rect 17122 2814 17128 2848
rect 17082 2776 17128 2814
rect 17082 2742 17088 2776
rect 17122 2742 17128 2776
rect 17082 2704 17128 2742
rect 17082 2670 17088 2704
rect 17122 2670 17128 2704
rect 17082 2632 17128 2670
rect 17082 2598 17088 2632
rect 17122 2598 17128 2632
rect 17082 2559 17128 2598
rect 17082 2525 17088 2559
rect 17122 2525 17128 2559
rect 17082 2486 17128 2525
rect 17082 2452 17088 2486
rect 17122 2452 17128 2486
rect 17082 2413 17128 2452
rect 17082 2379 17088 2413
rect 17122 2379 17128 2413
rect 17082 2340 17128 2379
rect 17082 2306 17088 2340
rect 17122 2306 17128 2340
rect 17082 2267 17128 2306
rect 17082 2233 17088 2267
rect 17122 2233 17128 2267
rect 17082 2194 17128 2233
rect 17082 2160 17088 2194
rect 17122 2160 17128 2194
rect 17082 2121 17128 2160
rect 17082 2087 17088 2121
rect 17122 2087 17128 2121
rect 17082 2048 17128 2087
rect 17082 2014 17088 2048
rect 17122 2014 17128 2048
tri 15024 1975 15041 1992 sw
rect 17082 1975 17128 2014
rect 14884 1958 15041 1975
tri 15041 1958 15058 1975 sw
rect 14884 1952 16866 1958
rect 14884 1918 14896 1952
rect 14930 1918 14971 1952
rect 15005 1918 15046 1952
rect 15080 1918 15121 1952
rect 15155 1918 15196 1952
rect 15230 1918 15271 1952
rect 15305 1918 15346 1952
rect 15380 1918 15420 1952
rect 15454 1918 15494 1952
rect 15528 1918 15568 1952
rect 15602 1918 15642 1952
rect 15676 1918 15716 1952
rect 15750 1918 15790 1952
rect 15824 1918 15864 1952
rect 15898 1918 15938 1952
rect 15972 1918 16012 1952
rect 16046 1918 16086 1952
rect 16120 1918 16160 1952
rect 16194 1918 16234 1952
rect 16268 1918 16308 1952
rect 16342 1918 16382 1952
rect 16416 1918 16456 1952
rect 16490 1918 16530 1952
rect 16564 1918 16604 1952
rect 16638 1918 16866 1952
rect 14884 1912 16866 1918
rect 17082 1941 17088 1975
rect 17122 1941 17128 1975
tri 15671 1902 15681 1912 ne
rect 15681 1902 15789 1912
tri 15789 1902 15799 1912 nw
rect 17082 1902 17128 1941
rect 14529 1848 14575 1889
tri 15681 1878 15705 1902 ne
rect 14529 1814 14535 1848
rect 14569 1814 14575 1848
rect 14529 1773 14575 1814
rect 14529 1739 14535 1773
rect 14569 1739 14575 1773
tri 11962 1722 11964 1724 sw
tri 14527 1722 14529 1724 se
rect 14529 1722 14575 1739
tri 14575 1722 14577 1724 sw
rect 11916 1690 11964 1722
tri 11964 1690 11996 1722 sw
tri 14495 1690 14527 1722 se
rect 14527 1690 14577 1722
tri 14577 1690 14609 1722 sw
rect 11916 1684 15661 1690
tri 9685 1644 9691 1650 se
rect 9691 1644 9751 1650
rect 11916 1650 11994 1684
rect 12028 1650 12068 1684
rect 12102 1650 12142 1684
rect 12176 1650 12216 1684
rect 12250 1650 12290 1684
rect 12324 1650 12364 1684
rect 12398 1650 12438 1684
rect 12472 1650 12512 1684
rect 12546 1650 12586 1684
rect 12620 1650 12660 1684
rect 12694 1650 12734 1684
rect 12768 1650 12808 1684
rect 12842 1650 12882 1684
rect 12916 1650 12956 1684
rect 12990 1650 13030 1684
rect 13064 1650 13104 1684
rect 13138 1650 13178 1684
rect 13212 1650 13252 1684
rect 13286 1650 13326 1684
rect 13360 1650 13399 1684
rect 13433 1650 13472 1684
rect 13506 1650 13545 1684
rect 13579 1650 13618 1684
rect 13652 1650 13691 1684
rect 13725 1650 13764 1684
rect 13798 1650 13837 1684
rect 13871 1650 13910 1684
rect 13944 1650 13983 1684
rect 14017 1650 14056 1684
rect 14090 1650 14129 1684
rect 14163 1650 14202 1684
rect 14236 1650 14275 1684
rect 14309 1650 14348 1684
rect 14382 1650 14421 1684
rect 14455 1650 14494 1684
rect 14528 1650 14567 1684
rect 14601 1650 14640 1684
rect 14674 1650 14713 1684
rect 14747 1650 14786 1684
rect 14820 1650 14859 1684
rect 14893 1650 14932 1684
rect 14966 1650 15005 1684
rect 15039 1650 15078 1684
rect 15112 1650 15151 1684
rect 15185 1650 15224 1684
rect 15258 1650 15297 1684
rect 15331 1650 15370 1684
rect 15404 1650 15443 1684
rect 15477 1650 15516 1684
rect 15550 1650 15589 1684
rect 15623 1650 15661 1684
rect 11916 1644 15661 1650
tri 9665 1624 9685 1644 se
rect 9685 1624 9751 1644
rect 8180 1002 8186 1054
rect 8238 1002 8264 1054
rect 8316 1002 8322 1054
rect 8180 978 8322 1002
rect 8180 926 8186 978
rect 8238 926 8264 978
rect 8316 926 8322 978
rect 8360 1094 9322 1146
rect 8360 1060 8366 1094
rect 8400 1074 9322 1094
tri 9355 1209 9376 1230 se
rect 9376 1209 9458 1230
rect 9355 1206 9458 1209
rect 9355 1196 9448 1206
tri 9448 1196 9458 1206 nw
rect 9592 1594 9751 1624
rect 8400 1060 8426 1074
tri 8426 1060 8440 1074 nw
rect 8360 1059 8425 1060
tri 8425 1059 8426 1060 nw
rect 8360 1019 8406 1059
tri 8406 1040 8425 1059 nw
rect 8360 985 8366 1019
rect 8400 985 8406 1019
rect 8360 944 8406 985
rect 7925 869 7977 910
rect 8360 910 8366 944
rect 8400 910 8406 944
rect 7925 835 7934 869
rect 7968 835 7977 869
rect 7925 794 7977 835
rect 7925 760 7934 794
rect 7968 760 7977 794
rect 7925 736 7977 760
rect 7925 672 7977 684
rect 7925 610 7934 620
rect 7968 610 7977 620
rect 7925 569 7977 610
rect 7925 535 7934 569
rect 7968 535 7977 569
rect 7925 494 7977 535
rect 7925 460 7934 494
rect 7968 460 7977 494
rect 7925 419 7977 460
rect 7925 385 7934 419
rect 7968 385 7977 419
rect 7925 344 7977 385
rect 7925 310 7934 344
rect 7968 310 7977 344
rect 7925 269 7977 310
rect 7925 235 7934 269
rect 7968 235 7977 269
rect 7925 194 7977 235
rect 7925 160 7934 194
rect 7968 160 7977 194
rect 7925 148 7977 160
rect 8141 892 8193 898
rect 8141 828 8193 840
rect 8141 733 8193 776
rect 8141 699 8150 733
rect 8184 699 8193 733
rect 8141 656 8193 699
rect 8141 622 8150 656
rect 8184 622 8193 656
rect 8141 579 8193 622
rect 8141 545 8150 579
rect 8184 545 8193 579
rect 8141 502 8193 545
rect 8141 468 8150 502
rect 8184 468 8193 502
rect 8141 425 8193 468
rect 8141 391 8150 425
rect 8184 391 8193 425
rect 8141 348 8193 391
rect 8141 314 8150 348
rect 8184 314 8193 348
rect 8141 271 8193 314
rect 8141 237 8150 271
rect 8184 237 8193 271
rect 8141 194 8193 237
rect 8141 160 8150 194
rect 8184 160 8193 194
rect 8141 148 8193 160
rect 8360 869 8406 910
rect 8360 835 8366 869
rect 8400 835 8406 869
rect 8360 794 8406 835
rect 8360 760 8366 794
rect 8400 760 8406 794
rect 8360 719 8406 760
rect 8360 685 8366 719
rect 8400 685 8406 719
rect 8360 644 8406 685
rect 8360 610 8366 644
rect 8400 610 8406 644
rect 8360 569 8406 610
rect 8360 535 8366 569
rect 8400 535 8406 569
rect 8360 494 8406 535
rect 8360 460 8366 494
rect 8400 460 8406 494
rect 8360 419 8406 460
rect 8360 385 8366 419
rect 8400 385 8406 419
rect 8360 344 8406 385
rect 8360 310 8366 344
rect 8400 310 8406 344
rect 8360 269 8406 310
rect 8360 235 8366 269
rect 8400 235 8406 269
rect 8360 194 8406 235
rect 8360 160 8366 194
rect 8400 160 8406 194
rect 8360 148 8406 160
rect 8573 1008 8625 1020
rect 8573 974 8582 1008
rect 8616 974 8625 1008
rect 8573 934 8625 974
rect 8573 900 8582 934
rect 8616 900 8625 934
rect 8573 892 8625 900
rect 8573 828 8582 840
rect 8616 828 8625 840
rect 8573 752 8582 776
rect 8616 752 8625 776
rect 8573 712 8625 752
rect 8573 678 8582 712
rect 8616 678 8625 712
rect 8573 638 8625 678
rect 8573 604 8582 638
rect 8616 604 8625 638
rect 8573 564 8625 604
rect 8573 530 8582 564
rect 8616 530 8625 564
rect 8573 490 8625 530
rect 8573 456 8582 490
rect 8616 456 8625 490
rect 8573 416 8625 456
rect 8573 382 8582 416
rect 8616 382 8625 416
rect 8573 342 8625 382
rect 8573 308 8582 342
rect 8616 308 8625 342
rect 8573 268 8625 308
rect 8573 234 8582 268
rect 8616 234 8625 268
rect 8573 194 8625 234
rect 8573 160 8582 194
rect 8616 160 8625 194
rect 8573 148 8625 160
rect 8789 1008 8841 1020
rect 8789 974 8798 1008
rect 8832 974 8841 1008
rect 8789 934 8841 974
rect 8789 900 8798 934
rect 8832 900 8841 934
rect 8789 860 8841 900
rect 8789 826 8798 860
rect 8832 826 8841 860
rect 8789 786 8841 826
rect 8789 752 8798 786
rect 8832 752 8841 786
rect 8789 712 8841 752
rect 8789 678 8798 712
rect 8832 678 8841 712
rect 8789 638 8841 678
rect 8789 604 8798 638
rect 8832 604 8841 638
rect 8789 564 8841 604
rect 8789 530 8798 564
rect 8832 530 8841 564
rect 8789 490 8841 530
rect 8789 456 8798 490
rect 8832 456 8841 490
rect 8789 416 8841 456
rect 8789 382 8798 416
rect 8832 382 8841 416
rect 8789 342 8841 382
rect 8789 308 8798 342
rect 8832 308 8841 342
rect 8789 268 8841 308
rect 8789 234 8798 268
rect 8832 234 8841 268
rect 8789 224 8841 234
rect 8789 160 8798 172
rect 8832 160 8841 172
rect 3504 121 3590 132
tri 3590 121 3601 132 sw
tri 3663 121 3674 132 ne
rect 3674 121 6629 132
tri 6629 121 6640 132 nw
rect 3504 120 3601 121
tri 3601 120 3602 121 sw
rect 3504 84 3602 120
tri 3602 84 3638 120 sw
tri 7193 84 7227 118 se
rect 7227 96 7279 108
rect 3504 80 3638 84
tri 3638 80 3642 84 sw
rect 3504 74 5680 80
rect 3504 40 3946 74
rect 3980 40 4020 74
rect 4054 40 4094 74
rect 4128 40 4168 74
rect 4202 40 4242 74
rect 4276 40 4316 74
rect 4350 40 4390 74
rect 4424 40 4464 74
rect 4498 40 4538 74
rect 4572 40 4612 74
rect 4646 40 4685 74
rect 4719 40 4758 74
rect 4792 40 4831 74
rect 4865 40 4904 74
rect 4938 40 4977 74
rect 5011 40 5050 74
rect 5084 40 5123 74
rect 5157 40 5196 74
rect 5230 40 5269 74
rect 5303 40 5342 74
rect 5376 40 5415 74
rect 5449 40 5488 74
rect 5522 40 5561 74
rect 5595 40 5634 74
rect 5668 40 5680 74
rect 3504 34 5680 40
rect 5877 78 7227 84
tri 7279 84 7313 118 sw
tri 8755 84 8789 118 se
rect 9005 1008 9057 1020
rect 9005 974 9014 1008
rect 9048 974 9057 1008
rect 9005 934 9057 974
rect 9005 900 9014 934
rect 9048 900 9057 934
rect 9005 892 9057 900
rect 9005 828 9014 840
rect 9048 828 9057 840
rect 9005 752 9014 776
rect 9048 752 9057 776
rect 9005 712 9057 752
rect 9005 678 9014 712
rect 9048 678 9057 712
rect 9005 638 9057 678
rect 9005 604 9014 638
rect 9048 604 9057 638
rect 9005 564 9057 604
rect 9005 530 9014 564
rect 9048 530 9057 564
rect 9005 490 9057 530
rect 9005 456 9014 490
rect 9048 456 9057 490
rect 9005 416 9057 456
rect 9005 382 9014 416
rect 9048 382 9057 416
rect 9005 342 9057 382
rect 9005 308 9014 342
rect 9048 308 9057 342
rect 9005 268 9057 308
rect 9005 234 9014 268
rect 9048 234 9057 268
rect 9005 194 9057 234
rect 9005 160 9014 194
rect 9048 160 9057 194
rect 9005 148 9057 160
rect 9221 1008 9273 1020
rect 9221 974 9230 1008
rect 9264 974 9273 1008
rect 9221 934 9273 974
rect 9221 900 9230 934
rect 9264 900 9273 934
rect 9221 860 9273 900
rect 9221 826 9230 860
rect 9264 826 9273 860
rect 9221 786 9273 826
rect 9221 752 9230 786
rect 9264 752 9273 786
rect 9221 712 9273 752
rect 9221 678 9230 712
rect 9264 678 9273 712
rect 9221 638 9273 678
rect 9221 604 9230 638
rect 9264 604 9273 638
rect 9355 736 9407 1196
tri 9407 1155 9448 1196 nw
rect 9355 672 9407 684
rect 9355 614 9407 620
rect 9437 1008 9489 1020
rect 9437 974 9446 1008
rect 9480 974 9489 1008
rect 9437 934 9489 974
rect 9437 900 9446 934
rect 9480 900 9489 934
rect 9437 892 9489 900
rect 9437 828 9446 840
rect 9480 828 9489 840
rect 9437 752 9446 776
rect 9480 752 9489 776
rect 9437 712 9489 752
rect 9437 678 9446 712
rect 9480 678 9489 712
rect 9437 638 9489 678
rect 9221 564 9273 604
rect 9221 530 9230 564
rect 9264 530 9273 564
rect 9221 490 9273 530
rect 9221 456 9230 490
rect 9264 456 9273 490
rect 9221 416 9273 456
rect 9221 382 9230 416
rect 9264 382 9273 416
rect 9221 342 9273 382
rect 9221 308 9230 342
rect 9264 308 9273 342
rect 9221 268 9273 308
rect 9221 234 9230 268
rect 9264 234 9273 268
rect 9221 224 9273 234
rect 9221 160 9230 172
rect 9264 160 9273 172
rect 8789 96 8841 108
rect 7279 78 8789 84
tri 8841 84 8875 118 sw
tri 9187 84 9221 118 se
rect 9437 604 9446 638
rect 9480 604 9489 638
rect 9437 564 9489 604
rect 9437 530 9446 564
rect 9480 530 9489 564
rect 9437 490 9489 530
rect 9437 456 9446 490
rect 9480 456 9489 490
rect 9437 416 9489 456
tri 9571 581 9592 602 se
rect 9592 581 9623 1594
tri 9623 1560 9657 1594 nw
rect 9693 1489 9699 1541
rect 9751 1489 9763 1541
rect 9815 1489 9821 1541
rect 9693 1236 9821 1489
rect 10514 1489 10520 1541
rect 10572 1489 10584 1541
rect 10636 1489 10642 1541
tri 9821 1236 9855 1270 sw
tri 10480 1236 10514 1270 se
rect 10514 1236 10642 1489
rect 12176 1409 12182 1461
rect 12234 1409 12246 1461
rect 12298 1409 12304 1461
tri 10642 1236 10676 1270 sw
tri 12142 1236 12176 1270 se
rect 12176 1236 12304 1409
rect 14456 1409 14462 1461
rect 14514 1409 14526 1461
rect 14578 1409 14584 1461
tri 12304 1236 12338 1270 sw
tri 14422 1236 14456 1270 se
rect 14456 1236 14584 1409
tri 14584 1236 14618 1270 sw
rect 9693 1230 11101 1236
rect 9693 1196 9705 1230
rect 9739 1196 9780 1230
rect 9814 1196 9855 1230
rect 9889 1196 9930 1230
rect 9964 1196 10005 1230
rect 10039 1196 10080 1230
rect 10114 1196 10155 1230
rect 10189 1196 10230 1230
rect 10264 1196 10305 1230
rect 10339 1196 10380 1230
rect 10414 1196 10455 1230
rect 10489 1196 10530 1230
rect 10564 1196 10605 1230
rect 10639 1196 10680 1230
rect 10714 1196 10755 1230
rect 10789 1196 10830 1230
rect 10864 1196 10905 1230
rect 10939 1196 10980 1230
rect 11014 1196 11055 1230
rect 11089 1196 11101 1230
rect 9693 1190 11101 1196
rect 11245 1230 15212 1236
rect 11245 1196 11257 1230
rect 11291 1196 11330 1230
rect 11364 1196 11403 1230
rect 11437 1196 11476 1230
rect 11510 1196 11549 1230
rect 11583 1196 11622 1230
rect 11656 1196 11695 1230
rect 11729 1196 11768 1230
rect 11802 1196 11841 1230
rect 11875 1196 11914 1230
rect 11948 1196 11987 1230
rect 12021 1196 12060 1230
rect 12094 1196 12133 1230
rect 12167 1196 12206 1230
rect 12240 1196 12279 1230
rect 12313 1196 12352 1230
rect 12386 1196 12425 1230
rect 12459 1196 12498 1230
rect 12532 1196 12571 1230
rect 12605 1196 12644 1230
rect 12678 1196 12717 1230
rect 12751 1196 12790 1230
rect 12824 1196 12863 1230
rect 12897 1196 12936 1230
rect 12970 1196 13009 1230
rect 13043 1196 13082 1230
rect 13116 1196 13155 1230
rect 13189 1196 13228 1230
rect 13262 1196 13301 1230
rect 13335 1196 13374 1230
rect 13408 1196 13447 1230
rect 13481 1196 13520 1230
rect 13554 1196 13593 1230
rect 13627 1196 13666 1230
rect 13700 1196 13739 1230
rect 13773 1196 13812 1230
rect 13846 1196 13885 1230
rect 13919 1196 13958 1230
rect 13992 1196 14031 1230
rect 14065 1196 14104 1230
rect 14138 1196 14177 1230
rect 14211 1196 14250 1230
rect 14284 1196 14323 1230
rect 14357 1196 14396 1230
rect 14430 1196 14469 1230
rect 14503 1196 14542 1230
rect 14576 1196 14615 1230
rect 14649 1196 14688 1230
rect 14722 1196 14761 1230
rect 14795 1196 14833 1230
rect 14867 1196 14905 1230
rect 14939 1196 14977 1230
rect 15011 1196 15212 1230
rect 11245 1190 15212 1196
rect 15240 1230 15415 1236
rect 15240 1196 15252 1230
rect 15286 1196 15369 1230
rect 15403 1196 15415 1230
rect 15240 1190 15415 1196
tri 15132 1156 15166 1190 ne
rect 9869 1094 9921 1106
rect 9869 1060 9878 1094
rect 9912 1060 9921 1094
rect 9571 575 9623 581
rect 9571 511 9623 523
rect 9571 453 9623 459
rect 9653 1008 9705 1020
rect 9653 974 9662 1008
rect 9696 974 9705 1008
rect 9653 934 9705 974
rect 9653 900 9662 934
rect 9696 900 9705 934
rect 9653 860 9705 900
rect 9653 826 9662 860
rect 9696 826 9705 860
rect 9653 786 9705 826
rect 9653 752 9662 786
rect 9696 752 9705 786
rect 9653 712 9705 752
rect 9653 678 9662 712
rect 9696 678 9705 712
rect 9653 638 9705 678
rect 9653 604 9662 638
rect 9696 604 9705 638
rect 9653 564 9705 604
rect 9653 530 9662 564
rect 9696 530 9705 564
rect 9653 490 9705 530
rect 9653 456 9662 490
rect 9696 456 9705 490
rect 9437 382 9446 416
rect 9480 382 9489 416
rect 9437 342 9489 382
rect 9437 308 9446 342
rect 9480 308 9489 342
rect 9437 268 9489 308
rect 9437 234 9446 268
rect 9480 234 9489 268
rect 9437 194 9489 234
rect 9437 160 9446 194
rect 9480 160 9489 194
rect 9437 148 9489 160
rect 9653 416 9705 456
rect 9653 382 9662 416
rect 9696 382 9705 416
rect 9653 342 9705 382
rect 9653 308 9662 342
rect 9696 308 9705 342
rect 9653 268 9705 308
rect 9653 234 9662 268
rect 9696 234 9705 268
rect 9653 224 9705 234
rect 9653 160 9662 172
rect 9696 160 9705 172
rect 9221 96 9273 108
rect 8841 78 9221 84
tri 9273 84 9307 118 sw
tri 9619 84 9653 118 se
rect 9869 1019 9921 1060
rect 9869 985 9878 1019
rect 9912 985 9921 1019
rect 9869 944 9921 985
rect 9869 910 9878 944
rect 9912 910 9921 944
rect 9869 892 9921 910
rect 9869 835 9878 840
rect 9912 835 9921 840
rect 9869 828 9921 835
rect 9869 760 9878 776
rect 9912 760 9921 776
rect 9869 719 9921 760
rect 9869 685 9878 719
rect 9912 685 9921 719
rect 9869 644 9921 685
rect 9869 610 9878 644
rect 9912 610 9921 644
rect 9869 569 9921 610
rect 9869 535 9878 569
rect 9912 535 9921 569
rect 9869 494 9921 535
rect 9869 460 9878 494
rect 9912 460 9921 494
rect 9869 419 9921 460
rect 9869 385 9878 419
rect 9912 385 9921 419
rect 9869 344 9921 385
rect 9869 310 9878 344
rect 9912 310 9921 344
rect 9869 269 9921 310
rect 9869 235 9878 269
rect 9912 235 9921 269
rect 9869 194 9921 235
rect 9869 160 9878 194
rect 9912 160 9921 194
rect 9869 148 9921 160
rect 10085 1094 10137 1106
rect 10085 1060 10094 1094
rect 10128 1060 10137 1094
rect 10085 1048 10137 1060
rect 10517 1094 10569 1106
rect 10517 1060 10526 1094
rect 10560 1060 10569 1094
rect 10517 1048 10569 1060
rect 10085 985 10094 996
rect 10128 985 10137 996
rect 10085 984 10137 985
rect 10085 910 10094 932
rect 10128 910 10137 932
rect 10085 869 10137 910
rect 10085 835 10094 869
rect 10128 835 10137 869
rect 10085 794 10137 835
rect 10085 760 10094 794
rect 10128 760 10137 794
rect 10085 719 10137 760
rect 10085 685 10094 719
rect 10128 685 10137 719
rect 10085 644 10137 685
rect 10085 610 10094 644
rect 10128 610 10137 644
rect 10085 569 10137 610
rect 10085 535 10094 569
rect 10128 535 10137 569
rect 10085 494 10137 535
rect 10085 460 10094 494
rect 10128 460 10137 494
rect 10085 419 10137 460
rect 10085 385 10094 419
rect 10128 385 10137 419
rect 10085 344 10137 385
rect 10085 310 10094 344
rect 10128 310 10137 344
rect 10085 269 10137 310
rect 10085 235 10094 269
rect 10128 235 10137 269
rect 10085 194 10137 235
rect 10085 160 10094 194
rect 10128 160 10137 194
rect 10085 148 10137 160
rect 10301 1008 10353 1020
rect 10301 974 10310 1008
rect 10344 974 10353 1008
rect 10301 934 10353 974
rect 10301 900 10310 934
rect 10344 900 10353 934
rect 10301 892 10353 900
rect 10301 828 10310 840
rect 10344 828 10353 840
rect 10301 752 10310 776
rect 10344 752 10353 776
rect 10301 712 10353 752
rect 10301 678 10310 712
rect 10344 678 10353 712
rect 10301 638 10353 678
rect 10301 604 10310 638
rect 10344 604 10353 638
rect 10301 564 10353 604
rect 10301 530 10310 564
rect 10344 530 10353 564
rect 10301 490 10353 530
rect 10301 456 10310 490
rect 10344 456 10353 490
rect 10301 416 10353 456
rect 10301 382 10310 416
rect 10344 382 10353 416
rect 10301 342 10353 382
rect 10301 308 10310 342
rect 10344 308 10353 342
rect 10301 268 10353 308
rect 10301 234 10310 268
rect 10344 234 10353 268
rect 10301 194 10353 234
rect 10301 160 10310 194
rect 10344 160 10353 194
rect 10301 148 10353 160
rect 10949 1094 11001 1106
rect 10949 1060 10958 1094
rect 10992 1060 11001 1094
rect 10949 1048 11001 1060
rect 10517 985 10526 996
rect 10560 985 10569 996
rect 10517 984 10569 985
rect 10517 910 10526 932
rect 10560 910 10569 932
rect 10517 869 10569 910
rect 10517 835 10526 869
rect 10560 835 10569 869
rect 10517 794 10569 835
rect 10517 760 10526 794
rect 10560 760 10569 794
rect 10517 719 10569 760
rect 10517 685 10526 719
rect 10560 685 10569 719
rect 10517 644 10569 685
rect 10517 610 10526 644
rect 10560 610 10569 644
rect 10517 569 10569 610
rect 10517 535 10526 569
rect 10560 535 10569 569
rect 10517 494 10569 535
rect 10517 460 10526 494
rect 10560 460 10569 494
rect 10517 419 10569 460
rect 10517 385 10526 419
rect 10560 385 10569 419
rect 10517 344 10569 385
rect 10517 310 10526 344
rect 10560 310 10569 344
rect 10517 269 10569 310
rect 10517 235 10526 269
rect 10560 235 10569 269
rect 10517 194 10569 235
rect 10517 160 10526 194
rect 10560 160 10569 194
rect 10517 148 10569 160
rect 10733 1008 10785 1020
rect 10733 974 10742 1008
rect 10776 974 10785 1008
rect 10733 934 10785 974
rect 10733 900 10742 934
rect 10776 900 10785 934
rect 10733 892 10785 900
rect 10733 828 10742 840
rect 10776 828 10785 840
rect 10733 752 10742 776
rect 10776 752 10785 776
rect 10733 712 10785 752
rect 10733 678 10742 712
rect 10776 678 10785 712
rect 10733 638 10785 678
rect 10733 604 10742 638
rect 10776 604 10785 638
rect 10733 564 10785 604
rect 10733 530 10742 564
rect 10776 530 10785 564
rect 10733 490 10785 530
rect 10733 456 10742 490
rect 10776 456 10785 490
rect 10733 416 10785 456
rect 10733 382 10742 416
rect 10776 382 10785 416
rect 10733 342 10785 382
rect 10733 308 10742 342
rect 10776 308 10785 342
rect 10733 268 10785 308
rect 10733 234 10742 268
rect 10776 234 10785 268
rect 10733 194 10785 234
rect 10733 160 10742 194
rect 10776 160 10785 194
rect 10733 148 10785 160
rect 11381 1094 11433 1106
rect 11381 1060 11390 1094
rect 11424 1060 11433 1094
rect 11381 1048 11433 1060
rect 10949 985 10958 996
rect 10992 985 11001 996
rect 10949 984 11001 985
rect 10949 910 10958 932
rect 10992 910 11001 932
rect 10949 869 11001 910
rect 10949 835 10958 869
rect 10992 835 11001 869
rect 10949 794 11001 835
rect 10949 760 10958 794
rect 10992 760 11001 794
rect 10949 719 11001 760
rect 10949 685 10958 719
rect 10992 685 11001 719
rect 10949 644 11001 685
rect 10949 610 10958 644
rect 10992 610 11001 644
rect 10949 569 11001 610
rect 10949 535 10958 569
rect 10992 535 11001 569
rect 10949 494 11001 535
rect 10949 460 10958 494
rect 10992 460 11001 494
rect 10949 419 11001 460
rect 10949 385 10958 419
rect 10992 385 11001 419
rect 10949 344 11001 385
rect 10949 310 10958 344
rect 10992 310 11001 344
rect 10949 269 11001 310
rect 10949 235 10958 269
rect 10992 235 11001 269
rect 10949 194 11001 235
rect 10949 160 10958 194
rect 10992 160 11001 194
rect 10949 148 11001 160
rect 11165 1008 11217 1020
rect 11165 974 11174 1008
rect 11208 974 11217 1008
rect 11165 934 11217 974
rect 11165 900 11174 934
rect 11208 900 11217 934
rect 11165 892 11217 900
rect 11165 828 11174 840
rect 11208 828 11217 840
rect 11165 752 11174 776
rect 11208 752 11217 776
rect 11165 712 11217 752
rect 11165 678 11174 712
rect 11208 678 11217 712
rect 11165 638 11217 678
rect 11165 604 11174 638
rect 11208 604 11217 638
rect 11165 564 11217 604
rect 11165 530 11174 564
rect 11208 530 11217 564
rect 11165 490 11217 530
rect 11165 456 11174 490
rect 11208 456 11217 490
rect 11165 416 11217 456
rect 11165 382 11174 416
rect 11208 382 11217 416
rect 11165 342 11217 382
rect 11165 308 11174 342
rect 11208 308 11217 342
rect 11165 268 11217 308
rect 11165 234 11174 268
rect 11208 234 11217 268
rect 11165 194 11217 234
rect 11165 160 11174 194
rect 11208 160 11217 194
rect 11165 148 11217 160
rect 11814 1094 11866 1106
rect 11814 1060 11823 1094
rect 11857 1060 11866 1094
rect 11814 1048 11866 1060
rect 11381 985 11390 996
rect 11424 985 11433 996
rect 11381 984 11433 985
rect 11381 910 11390 932
rect 11424 910 11433 932
rect 11381 869 11433 910
rect 11381 835 11390 869
rect 11424 835 11433 869
rect 11381 794 11433 835
rect 11381 760 11390 794
rect 11424 760 11433 794
rect 11381 719 11433 760
rect 11381 685 11390 719
rect 11424 685 11433 719
rect 11381 644 11433 685
rect 11381 610 11390 644
rect 11424 610 11433 644
rect 11381 569 11433 610
rect 11381 535 11390 569
rect 11424 535 11433 569
rect 11381 494 11433 535
rect 11381 460 11390 494
rect 11424 460 11433 494
rect 11381 419 11433 460
rect 11381 385 11390 419
rect 11424 385 11433 419
rect 11381 344 11433 385
rect 11381 310 11390 344
rect 11424 310 11433 344
rect 11381 269 11433 310
rect 11381 235 11390 269
rect 11424 235 11433 269
rect 11381 194 11433 235
rect 11381 160 11390 194
rect 11424 160 11433 194
rect 11381 148 11433 160
rect 11597 1008 11649 1020
rect 11597 974 11606 1008
rect 11640 974 11649 1008
rect 11597 934 11649 974
rect 11597 900 11606 934
rect 11640 900 11649 934
rect 11597 892 11649 900
rect 11597 828 11606 840
rect 11640 828 11649 840
rect 11597 752 11606 776
rect 11640 752 11649 776
rect 11597 712 11649 752
rect 11597 678 11606 712
rect 11640 678 11649 712
rect 11597 638 11649 678
rect 11597 604 11606 638
rect 11640 604 11649 638
rect 11597 564 11649 604
rect 11597 530 11606 564
rect 11640 530 11649 564
rect 11597 490 11649 530
rect 11597 456 11606 490
rect 11640 456 11649 490
rect 11597 416 11649 456
rect 11597 382 11606 416
rect 11640 382 11649 416
rect 11597 342 11649 382
rect 11597 308 11606 342
rect 11640 308 11649 342
rect 11597 268 11649 308
rect 11597 234 11606 268
rect 11640 234 11649 268
rect 11597 194 11649 234
rect 11597 160 11606 194
rect 11640 160 11649 194
rect 11597 148 11649 160
rect 12245 1094 12297 1106
rect 12245 1060 12254 1094
rect 12288 1060 12297 1094
rect 12245 1048 12297 1060
rect 11814 985 11823 996
rect 11857 985 11866 996
rect 11814 984 11866 985
rect 11814 910 11823 932
rect 11857 910 11866 932
rect 11814 869 11866 910
rect 11814 835 11823 869
rect 11857 835 11866 869
rect 11814 794 11866 835
rect 11814 760 11823 794
rect 11857 760 11866 794
rect 11814 719 11866 760
rect 11814 685 11823 719
rect 11857 685 11866 719
rect 11814 644 11866 685
rect 11814 610 11823 644
rect 11857 610 11866 644
rect 11814 569 11866 610
rect 11814 535 11823 569
rect 11857 535 11866 569
rect 11814 494 11866 535
rect 11814 460 11823 494
rect 11857 460 11866 494
rect 11814 419 11866 460
rect 11814 385 11823 419
rect 11857 385 11866 419
rect 11814 344 11866 385
rect 11814 310 11823 344
rect 11857 310 11866 344
rect 11814 269 11866 310
rect 11814 235 11823 269
rect 11857 235 11866 269
rect 11814 194 11866 235
rect 11814 160 11823 194
rect 11857 160 11866 194
rect 11814 148 11866 160
rect 12029 1008 12081 1020
rect 12029 974 12038 1008
rect 12072 974 12081 1008
rect 12029 934 12081 974
rect 12029 900 12038 934
rect 12072 900 12081 934
rect 12029 892 12081 900
rect 12029 828 12038 840
rect 12072 828 12081 840
rect 12029 752 12038 776
rect 12072 752 12081 776
rect 12029 712 12081 752
rect 12029 678 12038 712
rect 12072 678 12081 712
rect 12029 638 12081 678
rect 12029 604 12038 638
rect 12072 604 12081 638
rect 12029 564 12081 604
rect 12029 530 12038 564
rect 12072 530 12081 564
rect 12029 490 12081 530
rect 12029 456 12038 490
rect 12072 456 12081 490
rect 12029 416 12081 456
rect 12029 382 12038 416
rect 12072 382 12081 416
rect 12029 342 12081 382
rect 12029 308 12038 342
rect 12072 308 12081 342
rect 12029 268 12081 308
rect 12029 234 12038 268
rect 12072 234 12081 268
rect 12029 194 12081 234
rect 12029 160 12038 194
rect 12072 160 12081 194
rect 12029 148 12081 160
rect 15166 1093 15212 1190
rect 15705 1106 15765 1902
tri 15765 1878 15789 1902 nw
rect 17082 1868 17088 1902
rect 17122 1868 17128 1902
rect 17082 1829 17128 1868
rect 17082 1795 17088 1829
rect 17122 1795 17128 1829
rect 17082 1756 17128 1795
tri 17080 1722 17082 1724 se
rect 17082 1722 17088 1756
rect 17122 1722 17128 1756
tri 17048 1690 17080 1722 se
rect 17080 1690 17128 1722
rect 15817 1684 17128 1690
rect 15817 1650 15855 1684
rect 15889 1650 15929 1684
rect 15963 1650 16003 1684
rect 16037 1650 16077 1684
rect 16111 1650 16151 1684
rect 16185 1650 16225 1684
rect 16259 1650 16299 1684
rect 16333 1650 16373 1684
rect 16407 1650 16447 1684
rect 16481 1650 16521 1684
rect 16555 1650 16595 1684
rect 16629 1650 16668 1684
rect 16702 1650 16741 1684
rect 16775 1650 16814 1684
rect 16848 1650 16887 1684
rect 16921 1650 16960 1684
rect 16994 1650 17128 1684
rect 15817 1644 17128 1650
rect 15817 1230 16013 1236
rect 15817 1196 15829 1230
rect 15863 1196 15913 1230
rect 15947 1196 16013 1230
rect 15817 1190 16013 1196
tri 15927 1156 15961 1190 ne
tri 15765 1106 15794 1135 sw
rect 15166 1059 15172 1093
rect 15206 1059 15212 1093
rect 12245 985 12254 996
rect 12288 985 12297 996
rect 12245 984 12297 985
rect 12245 910 12254 932
rect 12288 910 12297 932
rect 12245 869 12297 910
rect 12245 835 12254 869
rect 12288 835 12297 869
rect 12245 794 12297 835
rect 12245 760 12254 794
rect 12288 760 12297 794
rect 12245 719 12297 760
rect 12245 685 12254 719
rect 12288 685 12297 719
rect 12245 644 12297 685
rect 12245 610 12254 644
rect 12288 610 12297 644
rect 12245 569 12297 610
rect 12245 535 12254 569
rect 12288 535 12297 569
rect 12245 494 12297 535
rect 12245 460 12254 494
rect 12288 460 12297 494
rect 12245 419 12297 460
rect 12245 385 12254 419
rect 12288 385 12297 419
rect 12245 344 12297 385
rect 12245 310 12254 344
rect 12288 310 12297 344
rect 12245 269 12297 310
rect 12245 235 12254 269
rect 12288 235 12297 269
rect 12245 194 12297 235
rect 12245 160 12254 194
rect 12288 160 12297 194
rect 12245 148 12297 160
rect 12461 1008 12513 1020
rect 12461 974 12470 1008
rect 12504 974 12513 1008
rect 12461 934 12513 974
rect 12461 900 12470 934
rect 12504 900 12513 934
rect 12461 892 12513 900
rect 12461 828 12470 840
rect 12504 828 12513 840
rect 12461 752 12470 776
rect 12504 752 12513 776
rect 12461 712 12513 752
rect 12461 678 12470 712
rect 12504 678 12513 712
rect 12461 638 12513 678
rect 12461 604 12470 638
rect 12504 604 12513 638
rect 12461 564 12513 604
rect 12461 530 12470 564
rect 12504 530 12513 564
rect 12461 490 12513 530
rect 12461 456 12470 490
rect 12504 456 12513 490
rect 12461 416 12513 456
rect 12461 382 12470 416
rect 12504 382 12513 416
rect 12461 342 12513 382
rect 12461 308 12470 342
rect 12504 308 12513 342
rect 12461 268 12513 308
rect 12461 234 12470 268
rect 12504 234 12513 268
rect 12461 194 12513 234
rect 12461 160 12470 194
rect 12504 160 12513 194
rect 12461 148 12513 160
rect 12677 1008 12729 1020
rect 12677 974 12686 1008
rect 12720 974 12729 1008
rect 12677 934 12729 974
rect 12677 900 12686 934
rect 12720 900 12729 934
rect 12677 860 12729 900
rect 12677 826 12686 860
rect 12720 826 12729 860
rect 12677 786 12729 826
rect 12677 752 12686 786
rect 12720 752 12729 786
rect 12677 712 12729 752
rect 12677 678 12686 712
rect 12720 678 12729 712
rect 12677 638 12729 678
rect 12677 604 12686 638
rect 12720 604 12729 638
rect 12677 564 12729 604
rect 12677 530 12686 564
rect 12720 530 12729 564
rect 12677 490 12729 530
rect 12677 456 12686 490
rect 12720 456 12729 490
rect 12677 416 12729 456
rect 12677 382 12686 416
rect 12720 382 12729 416
rect 12677 342 12729 382
rect 12677 308 12686 342
rect 12720 308 12729 342
rect 12677 268 12729 308
rect 12677 234 12686 268
rect 12720 234 12729 268
rect 12677 224 12729 234
rect 12677 160 12686 172
rect 12720 160 12729 172
rect 9653 96 9705 108
rect 9273 78 9653 84
tri 9705 84 9739 118 sw
tri 12643 84 12677 118 se
rect 12893 1008 12945 1020
rect 12893 974 12902 1008
rect 12936 974 12945 1008
rect 12893 934 12945 974
rect 12893 900 12902 934
rect 12936 900 12945 934
rect 12893 892 12945 900
rect 12893 828 12902 840
rect 12936 828 12945 840
rect 12893 752 12902 776
rect 12936 752 12945 776
rect 12893 712 12945 752
rect 12893 678 12902 712
rect 12936 678 12945 712
rect 12893 638 12945 678
rect 12893 604 12902 638
rect 12936 604 12945 638
rect 12893 564 12945 604
rect 12893 530 12902 564
rect 12936 530 12945 564
rect 12893 490 12945 530
rect 12893 456 12902 490
rect 12936 456 12945 490
rect 12893 416 12945 456
rect 12893 382 12902 416
rect 12936 382 12945 416
rect 12893 342 12945 382
rect 12893 308 12902 342
rect 12936 308 12945 342
rect 12893 268 12945 308
rect 12893 234 12902 268
rect 12936 234 12945 268
rect 12893 194 12945 234
rect 12893 160 12902 194
rect 12936 160 12945 194
rect 12893 148 12945 160
rect 13109 1008 13161 1020
rect 13109 974 13118 1008
rect 13152 974 13161 1008
rect 13109 934 13161 974
rect 13109 900 13118 934
rect 13152 900 13161 934
rect 13109 860 13161 900
rect 13109 826 13118 860
rect 13152 826 13161 860
rect 13109 786 13161 826
rect 13109 752 13118 786
rect 13152 752 13161 786
rect 13109 712 13161 752
rect 13109 678 13118 712
rect 13152 678 13161 712
rect 13109 638 13161 678
rect 13109 604 13118 638
rect 13152 604 13161 638
rect 13109 564 13161 604
rect 13109 530 13118 564
rect 13152 530 13161 564
rect 13109 490 13161 530
rect 13109 456 13118 490
rect 13152 456 13161 490
rect 13109 416 13161 456
rect 13109 382 13118 416
rect 13152 382 13161 416
rect 13109 342 13161 382
rect 13109 308 13118 342
rect 13152 308 13161 342
rect 13109 268 13161 308
rect 13109 234 13118 268
rect 13152 234 13161 268
rect 13109 224 13161 234
rect 13109 160 13118 172
rect 13152 160 13161 172
rect 12677 96 12729 108
rect 9705 78 12677 84
tri 12729 84 12763 118 sw
tri 13075 84 13109 118 se
rect 13325 1008 13377 1020
rect 13325 974 13334 1008
rect 13368 974 13377 1008
rect 13325 934 13377 974
rect 13325 900 13334 934
rect 13368 900 13377 934
rect 13325 892 13377 900
rect 13325 828 13334 840
rect 13368 828 13377 840
rect 13325 752 13334 776
rect 13368 752 13377 776
rect 13325 712 13377 752
rect 13325 678 13334 712
rect 13368 678 13377 712
rect 13325 638 13377 678
rect 13325 604 13334 638
rect 13368 604 13377 638
rect 13325 564 13377 604
rect 13325 530 13334 564
rect 13368 530 13377 564
rect 13325 490 13377 530
rect 13325 456 13334 490
rect 13368 456 13377 490
rect 13325 416 13377 456
rect 13325 382 13334 416
rect 13368 382 13377 416
rect 13325 342 13377 382
rect 13325 308 13334 342
rect 13368 308 13377 342
rect 13325 268 13377 308
rect 13325 234 13334 268
rect 13368 234 13377 268
rect 13325 194 13377 234
rect 13325 160 13334 194
rect 13368 160 13377 194
rect 13325 148 13377 160
rect 13541 1008 13593 1020
rect 13541 974 13550 1008
rect 13584 974 13593 1008
rect 13541 934 13593 974
rect 13541 900 13550 934
rect 13584 900 13593 934
rect 13541 860 13593 900
rect 13541 826 13550 860
rect 13584 826 13593 860
rect 13541 786 13593 826
rect 13541 752 13550 786
rect 13584 752 13593 786
rect 13541 712 13593 752
rect 13541 678 13550 712
rect 13584 678 13593 712
rect 13541 638 13593 678
rect 13541 604 13550 638
rect 13584 604 13593 638
rect 13541 564 13593 604
rect 13541 530 13550 564
rect 13584 530 13593 564
rect 13541 490 13593 530
rect 13541 456 13550 490
rect 13584 456 13593 490
rect 13541 416 13593 456
rect 13541 382 13550 416
rect 13584 382 13593 416
rect 13541 342 13593 382
rect 13541 308 13550 342
rect 13584 308 13593 342
rect 13541 268 13593 308
rect 13541 234 13550 268
rect 13584 234 13593 268
rect 13541 224 13593 234
rect 13541 160 13550 172
rect 13584 160 13593 172
rect 13109 96 13161 108
rect 12729 78 13109 84
tri 13161 84 13195 118 sw
tri 13507 84 13541 118 se
rect 13757 1008 13809 1020
rect 13757 974 13766 1008
rect 13800 974 13809 1008
rect 13757 934 13809 974
rect 13757 900 13766 934
rect 13800 900 13809 934
rect 13757 892 13809 900
rect 13757 828 13766 840
rect 13800 828 13809 840
rect 13757 752 13766 776
rect 13800 752 13809 776
rect 13757 712 13809 752
rect 13757 678 13766 712
rect 13800 678 13809 712
rect 13757 638 13809 678
rect 13757 604 13766 638
rect 13800 604 13809 638
rect 13757 564 13809 604
rect 13757 530 13766 564
rect 13800 530 13809 564
rect 13757 490 13809 530
rect 13757 456 13766 490
rect 13800 456 13809 490
rect 13757 416 13809 456
rect 13757 382 13766 416
rect 13800 382 13809 416
rect 13757 342 13809 382
rect 13757 308 13766 342
rect 13800 308 13809 342
rect 13757 268 13809 308
rect 13757 234 13766 268
rect 13800 234 13809 268
rect 13757 194 13809 234
rect 13757 160 13766 194
rect 13800 160 13809 194
rect 13757 148 13809 160
rect 13973 1008 14025 1020
rect 13973 974 13982 1008
rect 14016 974 14025 1008
rect 13973 934 14025 974
rect 13973 900 13982 934
rect 14016 900 14025 934
rect 13973 860 14025 900
rect 13973 826 13982 860
rect 14016 826 14025 860
rect 13973 786 14025 826
rect 13973 752 13982 786
rect 14016 752 14025 786
rect 13973 712 14025 752
rect 13973 678 13982 712
rect 14016 678 14025 712
rect 13973 638 14025 678
rect 13973 604 13982 638
rect 14016 604 14025 638
rect 13973 564 14025 604
rect 13973 530 13982 564
rect 14016 530 14025 564
rect 13973 490 14025 530
rect 13973 456 13982 490
rect 14016 456 14025 490
rect 13973 416 14025 456
rect 13973 382 13982 416
rect 14016 382 14025 416
rect 13973 342 14025 382
rect 13973 308 13982 342
rect 14016 308 14025 342
rect 13973 268 14025 308
rect 13973 234 13982 268
rect 14016 234 14025 268
rect 13973 224 14025 234
rect 13973 160 13982 172
rect 14016 160 14025 172
rect 13541 96 13593 108
rect 13161 78 13541 84
tri 13593 84 13627 118 sw
tri 13939 84 13973 118 se
rect 14189 1008 14241 1020
rect 14189 974 14198 1008
rect 14232 974 14241 1008
rect 14189 934 14241 974
rect 14189 900 14198 934
rect 14232 900 14241 934
rect 14189 892 14241 900
rect 14189 828 14198 840
rect 14232 828 14241 840
rect 14189 752 14198 776
rect 14232 752 14241 776
rect 14189 712 14241 752
rect 14189 678 14198 712
rect 14232 678 14241 712
rect 14189 638 14241 678
rect 14189 604 14198 638
rect 14232 604 14241 638
rect 14189 564 14241 604
rect 14189 530 14198 564
rect 14232 530 14241 564
rect 14189 490 14241 530
rect 14189 456 14198 490
rect 14232 456 14241 490
rect 14189 416 14241 456
rect 14189 382 14198 416
rect 14232 382 14241 416
rect 14189 342 14241 382
rect 14189 308 14198 342
rect 14232 308 14241 342
rect 14189 268 14241 308
rect 14189 234 14198 268
rect 14232 234 14241 268
rect 14189 194 14241 234
rect 14189 160 14198 194
rect 14232 160 14241 194
rect 14189 148 14241 160
rect 14405 1008 14457 1020
rect 14405 974 14414 1008
rect 14448 974 14457 1008
rect 14405 934 14457 974
rect 14405 900 14414 934
rect 14448 900 14457 934
rect 14405 860 14457 900
rect 14405 826 14414 860
rect 14448 826 14457 860
rect 14405 786 14457 826
rect 14405 752 14414 786
rect 14448 752 14457 786
rect 14405 712 14457 752
rect 14405 678 14414 712
rect 14448 678 14457 712
rect 14405 638 14457 678
rect 14405 604 14414 638
rect 14448 604 14457 638
rect 14405 564 14457 604
rect 14405 530 14414 564
rect 14448 530 14457 564
rect 14405 490 14457 530
rect 14405 456 14414 490
rect 14448 456 14457 490
rect 14405 416 14457 456
rect 14405 382 14414 416
rect 14448 382 14457 416
rect 14405 342 14457 382
rect 14405 308 14414 342
rect 14448 308 14457 342
rect 14405 268 14457 308
rect 14405 234 14414 268
rect 14448 234 14457 268
rect 14405 224 14457 234
rect 14405 160 14414 172
rect 14448 160 14457 172
rect 13973 96 14025 108
rect 13593 78 13973 84
tri 14025 84 14059 118 sw
tri 14371 84 14405 118 se
rect 14621 1008 14673 1020
rect 14621 974 14630 1008
rect 14664 974 14673 1008
rect 14621 934 14673 974
rect 14621 900 14630 934
rect 14664 900 14673 934
rect 14621 892 14673 900
rect 14621 828 14630 840
rect 14664 828 14673 840
rect 14621 752 14630 776
rect 14664 752 14673 776
rect 14621 712 14673 752
rect 14621 678 14630 712
rect 14664 678 14673 712
rect 14621 638 14673 678
rect 14621 604 14630 638
rect 14664 604 14673 638
rect 14621 564 14673 604
rect 14621 530 14630 564
rect 14664 530 14673 564
rect 14621 490 14673 530
rect 14621 456 14630 490
rect 14664 456 14673 490
rect 14621 416 14673 456
rect 14621 382 14630 416
rect 14664 382 14673 416
rect 14621 342 14673 382
rect 14621 308 14630 342
rect 14664 308 14673 342
rect 14621 268 14673 308
rect 14621 234 14630 268
rect 14664 234 14673 268
rect 14621 194 14673 234
rect 14621 160 14630 194
rect 14664 160 14673 194
rect 14621 148 14673 160
rect 14837 1008 14889 1020
rect 14837 974 14846 1008
rect 14880 974 14889 1008
rect 14837 934 14889 974
rect 14837 900 14846 934
rect 14880 900 14889 934
rect 14837 860 14889 900
rect 14837 826 14846 860
rect 14880 826 14889 860
rect 14837 786 14889 826
rect 14837 752 14846 786
rect 14880 752 14889 786
rect 14837 712 14889 752
rect 14837 678 14846 712
rect 14880 678 14889 712
rect 14837 638 14889 678
rect 14837 604 14846 638
rect 14880 604 14889 638
rect 14837 564 14889 604
rect 14837 530 14846 564
rect 14880 530 14889 564
rect 14837 490 14889 530
rect 14837 456 14846 490
rect 14880 456 14889 490
rect 14837 416 14889 456
rect 14837 382 14846 416
rect 14880 382 14889 416
rect 14837 342 14889 382
rect 14837 308 14846 342
rect 14880 308 14889 342
rect 14837 268 14889 308
rect 14837 234 14846 268
rect 14880 234 14889 268
rect 14837 224 14889 234
rect 14837 160 14846 172
rect 14880 160 14889 172
rect 14405 96 14457 108
rect 14025 78 14405 84
tri 14457 84 14491 118 sw
tri 14803 84 14837 118 se
rect 15053 1008 15105 1020
rect 15053 974 15062 1008
rect 15096 974 15105 1008
rect 15053 934 15105 974
rect 15053 900 15062 934
rect 15096 900 15105 934
rect 15053 892 15105 900
rect 15053 828 15062 840
rect 15096 828 15105 840
rect 15053 752 15062 776
rect 15096 752 15105 776
rect 15053 712 15105 752
rect 15053 678 15062 712
rect 15096 678 15105 712
rect 15053 638 15105 678
rect 15053 604 15062 638
rect 15096 604 15105 638
rect 15053 564 15105 604
rect 15053 530 15062 564
rect 15096 530 15105 564
rect 15166 1012 15212 1059
rect 15166 978 15172 1012
rect 15206 978 15212 1012
rect 15166 931 15212 978
rect 15166 897 15172 931
rect 15206 897 15212 931
rect 15166 850 15212 897
rect 15166 816 15172 850
rect 15206 816 15212 850
rect 15166 768 15212 816
rect 15166 734 15172 768
rect 15206 734 15212 768
rect 15166 686 15212 734
rect 15166 652 15172 686
rect 15206 652 15212 686
rect 15166 604 15212 652
rect 15166 570 15172 604
rect 15206 570 15212 604
rect 15166 558 15212 570
rect 15418 1093 15470 1105
rect 15418 1059 15428 1093
rect 15462 1059 15470 1093
rect 15418 1012 15470 1059
rect 15418 978 15428 1012
rect 15462 978 15470 1012
rect 15418 931 15470 978
rect 15418 897 15428 931
rect 15462 897 15470 931
rect 15418 850 15470 897
rect 15418 816 15428 850
rect 15462 816 15470 850
rect 15418 768 15470 816
rect 15418 734 15428 768
rect 15462 734 15470 768
rect 15418 686 15470 734
rect 15418 652 15428 686
rect 15462 652 15470 686
rect 15418 604 15470 652
rect 15418 570 15428 604
rect 15462 570 15470 604
rect 15053 490 15105 530
rect 15053 456 15062 490
rect 15096 456 15105 490
rect 15053 416 15105 456
rect 15053 382 15062 416
rect 15096 382 15105 416
rect 15053 342 15105 382
rect 15053 308 15062 342
rect 15096 308 15105 342
rect 15053 268 15105 308
rect 15053 234 15062 268
rect 15096 234 15105 268
rect 15053 194 15105 234
rect 15053 160 15062 194
rect 15096 160 15105 194
rect 15053 148 15105 160
rect 15418 224 15470 570
rect 15418 160 15470 172
rect 14837 96 14889 108
rect 14457 78 14837 84
tri 14889 84 14923 118 sw
tri 15384 84 15418 118 se
rect 15529 1094 15581 1106
rect 15529 1060 15538 1094
rect 15572 1060 15581 1094
rect 15529 1019 15581 1060
rect 15529 985 15538 1019
rect 15572 985 15581 1019
rect 15529 944 15581 985
rect 15529 910 15538 944
rect 15572 910 15581 944
rect 15529 869 15581 910
rect 15529 835 15538 869
rect 15572 835 15581 869
rect 15529 794 15581 835
rect 15529 760 15538 794
rect 15572 760 15581 794
rect 15529 719 15581 760
rect 15529 685 15538 719
rect 15572 685 15581 719
rect 15529 644 15581 685
rect 15529 610 15538 644
rect 15572 610 15581 644
rect 15529 569 15581 610
rect 15529 535 15538 569
rect 15572 535 15581 569
rect 15529 494 15581 535
rect 15529 460 15538 494
rect 15572 460 15581 494
rect 15529 419 15581 460
rect 15529 385 15538 419
rect 15572 385 15581 419
rect 15529 344 15581 385
rect 15529 332 15538 344
rect 15572 332 15581 344
rect 15529 269 15581 280
rect 15529 267 15538 269
rect 15572 267 15581 269
rect 15529 202 15581 215
rect 15529 144 15581 150
rect 15705 1094 15794 1106
rect 15705 1060 15754 1094
rect 15788 1060 15794 1094
rect 15705 1019 15794 1060
rect 15705 985 15754 1019
rect 15788 985 15794 1019
rect 15705 944 15794 985
rect 15705 910 15754 944
rect 15788 910 15794 944
rect 15705 869 15794 910
rect 15705 835 15754 869
rect 15788 835 15794 869
rect 15705 794 15794 835
rect 15705 760 15754 794
rect 15788 760 15794 794
rect 15705 719 15794 760
rect 15705 685 15754 719
rect 15788 685 15794 719
rect 15705 644 15794 685
rect 15705 610 15754 644
rect 15788 610 15794 644
rect 15705 569 15794 610
rect 15705 535 15754 569
rect 15788 535 15794 569
rect 15705 494 15794 535
rect 15705 460 15754 494
rect 15788 460 15794 494
rect 15705 419 15794 460
rect 15705 385 15754 419
rect 15788 385 15794 419
rect 15705 344 15794 385
rect 15705 310 15754 344
rect 15788 310 15794 344
rect 15705 269 15794 310
rect 15705 235 15754 269
rect 15788 235 15794 269
rect 15705 194 15794 235
rect 15705 160 15754 194
rect 15788 160 15794 194
rect 15705 148 15794 160
rect 15961 1094 16013 1190
rect 15961 1060 15970 1094
rect 16004 1060 16013 1094
rect 15961 1019 16013 1060
rect 15961 985 15970 1019
rect 16004 985 16013 1019
rect 15961 944 16013 985
rect 15961 910 15970 944
rect 16004 910 16013 944
rect 15961 869 16013 910
rect 15961 835 15970 869
rect 16004 835 16013 869
rect 15961 794 16013 835
rect 15961 760 15970 794
rect 16004 760 16013 794
rect 15961 719 16013 760
rect 15961 685 15970 719
rect 16004 685 16013 719
rect 15961 644 16013 685
rect 15961 610 15970 644
rect 16004 610 16013 644
rect 15961 569 16013 610
rect 15961 535 15970 569
rect 16004 535 16013 569
rect 15961 494 16013 535
rect 15961 460 15970 494
rect 16004 460 16013 494
rect 15961 419 16013 460
rect 15961 385 15970 419
rect 16004 385 16013 419
rect 15961 344 16013 385
rect 15961 332 15970 344
rect 16004 332 16013 344
rect 15961 269 16013 280
rect 15961 267 15970 269
rect 16004 267 16013 269
rect 15961 202 16013 215
rect 15961 144 16013 150
rect 15418 96 15470 108
rect 14889 78 15418 84
tri 15470 84 15504 118 sw
rect 15470 78 15997 84
rect 5877 44 5889 78
rect 5923 44 5962 78
rect 5996 44 6035 78
rect 6069 44 6108 78
rect 6142 44 6181 78
rect 6215 44 6254 78
rect 6288 44 6327 78
rect 6361 44 6400 78
rect 6434 44 6473 78
rect 6507 44 6546 78
rect 6580 44 6619 78
rect 6653 44 6692 78
rect 6726 44 6765 78
rect 6799 44 6838 78
rect 6872 44 6911 78
rect 6945 44 6984 78
rect 7018 44 7057 78
rect 7091 44 7130 78
rect 7164 44 7203 78
rect 7310 44 7349 78
rect 7383 44 7422 78
rect 7456 44 7495 78
rect 7529 44 7568 78
rect 7602 44 7641 78
rect 7675 44 7714 78
rect 7748 44 7787 78
rect 7821 44 7860 78
rect 7894 44 7933 78
rect 7967 44 8006 78
rect 8040 44 8079 78
rect 8113 44 8152 78
rect 8186 44 8225 78
rect 8259 44 8298 78
rect 8332 44 8371 78
rect 8405 44 8444 78
rect 8478 44 8517 78
rect 8551 44 8590 78
rect 8624 44 8663 78
rect 8697 44 8736 78
rect 8770 44 8789 78
rect 8843 44 8882 78
rect 8916 44 8955 78
rect 8989 44 9028 78
rect 9062 44 9101 78
rect 9135 44 9174 78
rect 9208 44 9221 78
rect 9281 44 9320 78
rect 9354 44 9393 78
rect 9427 44 9466 78
rect 9500 44 9539 78
rect 9573 44 9612 78
rect 9646 44 9653 78
rect 9719 44 9758 78
rect 9792 44 9831 78
rect 9865 44 9903 78
rect 9937 44 9975 78
rect 10009 44 10047 78
rect 10081 44 10119 78
rect 10153 44 10191 78
rect 10225 44 10263 78
rect 10297 44 10335 78
rect 10369 44 10407 78
rect 10441 44 10479 78
rect 10513 44 10551 78
rect 10585 44 10623 78
rect 10657 44 10695 78
rect 10729 44 10767 78
rect 10801 44 10839 78
rect 10873 44 10911 78
rect 10945 44 10983 78
rect 11017 44 11055 78
rect 11089 44 11127 78
rect 11161 44 11199 78
rect 11233 44 11271 78
rect 11305 44 11343 78
rect 11377 44 11415 78
rect 11449 44 11487 78
rect 11521 44 11559 78
rect 11593 44 11631 78
rect 11665 44 11703 78
rect 11737 44 11775 78
rect 11809 44 11847 78
rect 11881 44 11919 78
rect 11953 44 11991 78
rect 12025 44 12063 78
rect 12097 44 12135 78
rect 12169 44 12207 78
rect 12241 44 12279 78
rect 12313 44 12351 78
rect 12385 44 12423 78
rect 12457 44 12495 78
rect 12529 44 12567 78
rect 12601 44 12639 78
rect 12673 44 12677 78
rect 12745 44 12783 78
rect 12817 44 12855 78
rect 12889 44 12927 78
rect 12961 44 12999 78
rect 13033 44 13071 78
rect 13105 44 13109 78
rect 13177 44 13215 78
rect 13249 44 13287 78
rect 13321 44 13359 78
rect 13393 44 13431 78
rect 13465 44 13503 78
rect 13537 44 13541 78
rect 13609 44 13647 78
rect 13681 44 13719 78
rect 13753 44 13791 78
rect 13825 44 13863 78
rect 13897 44 13935 78
rect 13969 44 13973 78
rect 14041 44 14079 78
rect 14113 44 14151 78
rect 14185 44 14223 78
rect 14257 44 14295 78
rect 14329 44 14367 78
rect 14401 44 14405 78
rect 14473 44 14511 78
rect 14545 44 14583 78
rect 14617 44 14655 78
rect 14689 44 14727 78
rect 14761 44 14799 78
rect 14833 44 14837 78
rect 14905 44 14943 78
rect 14977 44 15015 78
rect 15049 44 15087 78
rect 15121 44 15159 78
rect 15193 44 15231 78
rect 15265 44 15303 78
rect 15337 44 15375 78
rect 15409 44 15418 78
rect 15481 44 15519 78
rect 15553 44 15591 78
rect 15625 44 15663 78
rect 15697 44 15735 78
rect 15769 44 15807 78
rect 15841 44 15879 78
rect 15913 44 15951 78
rect 15985 44 15997 78
rect 5877 38 15997 44
rect 3035 -885 3041 -833
rect 3093 -885 3131 -833
rect 3183 -867 15335 -833
rect 3183 -885 3189 -867
tri 3189 -885 3207 -867 nw
tri 15311 -885 15329 -867 ne
rect 15329 -885 15335 -867
rect 15387 -885 15399 -833
rect 15451 -885 15457 -833
<< via1 >>
rect -183 3030 -131 3082
rect -119 3030 -67 3082
rect 833 2891 885 2943
rect 897 2891 949 2943
rect 424 2198 433 2231
rect 433 2198 467 2231
rect 467 2198 476 2231
rect 424 2179 476 2198
rect 424 2158 476 2166
rect 424 2124 433 2158
rect 433 2124 467 2158
rect 467 2124 476 2158
rect 424 2114 476 2124
rect 711 2517 720 2544
rect 720 2517 754 2544
rect 754 2517 763 2544
rect 711 2492 763 2517
rect 711 2472 763 2480
rect 711 2438 720 2472
rect 720 2438 754 2472
rect 754 2438 763 2472
rect 711 2428 763 2438
rect 676 2028 728 2080
rect 740 2028 792 2080
rect 1023 2533 1032 2544
rect 1032 2533 1066 2544
rect 1066 2533 1075 2544
rect 1023 2492 1075 2533
rect 1023 2458 1032 2480
rect 1032 2458 1066 2480
rect 1066 2458 1075 2480
rect 1023 2428 1075 2458
rect 1133 2192 1185 2231
rect 1133 2179 1142 2192
rect 1142 2179 1176 2192
rect 1176 2179 1185 2192
rect 1133 2158 1142 2166
rect 1142 2158 1176 2166
rect 1176 2158 1185 2166
rect 1133 2117 1185 2158
rect 1133 2114 1142 2117
rect 1142 2114 1176 2117
rect 1176 2114 1185 2117
rect 1289 2833 1298 2843
rect 1298 2833 1332 2843
rect 1332 2833 1341 2843
rect 1289 2792 1341 2833
rect 1289 2791 1298 2792
rect 1298 2791 1332 2792
rect 1332 2791 1341 2792
rect 1289 2758 1298 2778
rect 1298 2758 1332 2778
rect 1332 2758 1341 2778
rect 1289 2726 1341 2758
rect 1289 2683 1298 2713
rect 1298 2683 1332 2713
rect 1332 2683 1341 2713
rect 1289 2661 1341 2683
rect 1289 2642 1341 2648
rect 1289 2608 1298 2642
rect 1298 2608 1332 2642
rect 1332 2608 1341 2642
rect 1289 2596 1341 2608
rect 1445 2200 1454 2231
rect 1454 2200 1488 2231
rect 1488 2200 1497 2231
rect 1445 2179 1497 2200
rect 1445 2154 1497 2166
rect 1445 2120 1454 2154
rect 1454 2120 1488 2154
rect 1488 2120 1497 2154
rect 1445 2114 1497 2120
rect 1601 2833 1610 2843
rect 1610 2833 1644 2843
rect 1644 2833 1653 2843
rect 1601 2792 1653 2833
rect 1601 2791 1610 2792
rect 1610 2791 1644 2792
rect 1644 2791 1653 2792
rect 1601 2758 1610 2778
rect 1610 2758 1644 2778
rect 1644 2758 1653 2778
rect 1601 2726 1653 2758
rect 1601 2683 1610 2713
rect 1610 2683 1644 2713
rect 1644 2683 1653 2713
rect 1601 2661 1653 2683
rect 1601 2642 1653 2648
rect 1601 2608 1610 2642
rect 1610 2608 1644 2642
rect 1644 2608 1653 2642
rect 1601 2596 1653 2608
rect 1757 2200 1766 2231
rect 1766 2200 1800 2231
rect 1800 2200 1809 2231
rect 1757 2179 1809 2200
rect 1757 2154 1809 2166
rect 1757 2120 1766 2154
rect 1766 2120 1800 2154
rect 1800 2120 1809 2154
rect 1757 2114 1809 2120
rect 1913 2833 1922 2843
rect 1922 2833 1956 2843
rect 1956 2833 1965 2843
rect 1913 2792 1965 2833
rect 1913 2791 1922 2792
rect 1922 2791 1956 2792
rect 1956 2791 1965 2792
rect 1913 2758 1922 2778
rect 1922 2758 1956 2778
rect 1956 2758 1965 2778
rect 1913 2726 1965 2758
rect 1913 2683 1922 2713
rect 1922 2683 1956 2713
rect 1956 2683 1965 2713
rect 1913 2661 1965 2683
rect 1913 2642 1965 2648
rect 1913 2608 1922 2642
rect 1922 2608 1956 2642
rect 1956 2608 1965 2642
rect 1913 2596 1965 2608
rect 1417 2028 1469 2080
rect 1481 2028 1533 2080
rect 2069 2192 2121 2231
rect 2069 2179 2078 2192
rect 2078 2179 2112 2192
rect 2112 2179 2121 2192
rect 2069 2158 2078 2166
rect 2078 2158 2112 2166
rect 2112 2158 2121 2166
rect 2069 2117 2121 2158
rect 2069 2114 2078 2117
rect 2078 2114 2112 2117
rect 2112 2114 2121 2117
rect 2225 2383 2234 2388
rect 2234 2383 2268 2388
rect 2268 2383 2277 2388
rect 2225 2342 2277 2383
rect 2225 2336 2234 2342
rect 2234 2336 2268 2342
rect 2268 2336 2277 2342
rect 2225 2308 2234 2324
rect 2234 2308 2268 2324
rect 2268 2308 2277 2324
rect 2225 2272 2277 2308
rect 2381 2192 2433 2231
rect 2381 2179 2390 2192
rect 2390 2179 2424 2192
rect 2424 2179 2433 2192
rect 2381 2158 2390 2166
rect 2390 2158 2424 2166
rect 2424 2158 2433 2166
rect 2381 2117 2433 2158
rect 2381 2114 2390 2117
rect 2390 2114 2424 2117
rect 2424 2114 2433 2117
rect 2537 2383 2546 2388
rect 2546 2383 2580 2388
rect 2580 2383 2589 2388
rect 2537 2342 2589 2383
rect 2537 2336 2546 2342
rect 2546 2336 2580 2342
rect 2580 2336 2589 2342
rect 2537 2308 2546 2324
rect 2546 2308 2580 2324
rect 2580 2308 2589 2324
rect 2537 2272 2589 2308
rect 2693 2192 2745 2231
rect 2693 2179 2702 2192
rect 2702 2179 2736 2192
rect 2736 2179 2745 2192
rect 2693 2158 2702 2166
rect 2702 2158 2736 2166
rect 2736 2158 2745 2166
rect 2693 2117 2745 2158
rect 2693 2114 2702 2117
rect 2702 2114 2736 2117
rect 2736 2114 2745 2117
rect 2849 2533 2858 2544
rect 2858 2533 2892 2544
rect 2892 2533 2901 2544
rect 2849 2492 2901 2533
rect 2849 2458 2858 2480
rect 2858 2458 2892 2480
rect 2892 2458 2901 2480
rect 2849 2428 2901 2458
rect 3005 2192 3057 2231
rect 3005 2179 3014 2192
rect 3014 2179 3048 2192
rect 3048 2179 3057 2192
rect 3005 2158 3014 2166
rect 3014 2158 3048 2166
rect 3048 2158 3057 2166
rect 3005 2117 3057 2158
rect 3005 2114 3014 2117
rect 3014 2114 3048 2117
rect 3048 2114 3057 2117
rect 3161 2533 3170 2544
rect 3170 2533 3204 2544
rect 3204 2533 3213 2544
rect 3161 2492 3213 2533
rect 3161 2458 3170 2480
rect 3170 2458 3204 2480
rect 3204 2458 3213 2480
rect 3161 2428 3213 2458
rect 3317 2192 3369 2231
rect 3317 2179 3326 2192
rect 3326 2179 3360 2192
rect 3360 2179 3369 2192
rect 3317 2158 3326 2166
rect 3326 2158 3360 2166
rect 3360 2158 3369 2166
rect 3317 2117 3369 2158
rect 3317 2114 3326 2117
rect 3326 2114 3360 2117
rect 3360 2114 3369 2117
rect 3629 2204 3638 2231
rect 3638 2204 3672 2231
rect 3672 2204 3681 2231
rect 3629 2179 3681 2204
rect 3629 2159 3681 2166
rect 3629 2125 3638 2159
rect 3638 2125 3672 2159
rect 3672 2125 3681 2159
rect 3629 2114 3681 2125
rect 3941 2210 3950 2231
rect 3950 2210 3984 2231
rect 3984 2210 3993 2231
rect 3941 2179 3993 2210
rect 3941 2132 3950 2166
rect 3950 2132 3984 2166
rect 3984 2132 3993 2166
rect 3941 2114 3993 2132
rect 4292 2805 4344 2857
rect 4292 2741 4344 2793
rect 4361 2213 4413 2231
rect 4361 2179 4372 2213
rect 4372 2179 4406 2213
rect 4406 2179 4413 2213
rect 4361 2131 4413 2166
rect 4361 2114 4372 2131
rect 4372 2114 4406 2131
rect 4406 2114 4413 2131
rect 2225 1873 2277 1882
rect 2225 1839 2239 1873
rect 2239 1839 2273 1873
rect 2273 1839 2277 1873
rect 2225 1830 2277 1839
rect 2289 1873 2341 1882
rect 2289 1839 2312 1873
rect 2312 1839 2341 1873
rect 2289 1830 2341 1839
rect 2756 1873 2808 1882
rect 2756 1839 2762 1873
rect 2762 1839 2796 1873
rect 2796 1839 2808 1873
rect 2756 1830 2808 1839
rect 2820 1873 2872 1882
rect 2820 1839 2845 1873
rect 2845 1839 2872 1873
rect 2820 1830 2872 1839
rect 827 1729 879 1781
rect 891 1729 943 1781
rect 4664 2201 4673 2231
rect 4673 2201 4707 2231
rect 4707 2201 4716 2231
rect 4664 2179 4716 2201
rect 4664 2161 4716 2166
rect 4664 2127 4673 2161
rect 4673 2127 4707 2161
rect 4707 2127 4716 2161
rect 4664 2114 4716 2127
rect 3978 1649 4030 1701
rect 4042 1649 4094 1701
rect 4787 1942 4839 1994
rect 4787 1878 4839 1930
rect 3556 1569 3608 1621
rect 3620 1569 3672 1621
rect 5221 2961 5273 3013
rect 5221 2897 5273 2949
rect 5221 2649 5273 2701
rect 5221 2585 5273 2637
rect 5626 2891 5678 2943
rect 5690 2891 5742 2943
rect 5348 2677 5400 2701
rect 5348 2649 5357 2677
rect 5357 2649 5391 2677
rect 5391 2649 5400 2677
rect 5348 2602 5400 2637
rect 5348 2585 5357 2602
rect 5357 2585 5391 2602
rect 5391 2585 5400 2602
rect 5493 2683 5502 2701
rect 5502 2683 5536 2701
rect 5536 2683 5545 2701
rect 5493 2649 5545 2683
rect 5493 2608 5502 2637
rect 5502 2608 5536 2637
rect 5536 2608 5545 2637
rect 5493 2585 5545 2608
rect 5803 2683 5812 2701
rect 5812 2683 5846 2701
rect 5846 2683 5855 2701
rect 5803 2649 5855 2683
rect 5803 2608 5812 2637
rect 5812 2608 5846 2637
rect 5846 2608 5855 2637
rect 5803 2585 5855 2608
rect 5619 2028 5671 2080
rect 5683 2028 5735 2080
rect 6021 2833 6030 2857
rect 6030 2833 6064 2857
rect 6064 2833 6073 2857
rect 6021 2805 6073 2833
rect 6021 2792 6073 2793
rect 6021 2758 6030 2792
rect 6030 2758 6064 2792
rect 6064 2758 6073 2792
rect 6021 2741 6073 2758
rect 6237 2683 6246 2701
rect 6246 2683 6280 2701
rect 6280 2683 6289 2701
rect 6237 2649 6289 2683
rect 6237 2608 6246 2637
rect 6246 2608 6280 2637
rect 6280 2608 6289 2637
rect 6237 2585 6289 2608
rect 6424 2805 6476 2857
rect 6424 2741 6476 2793
rect 5194 1841 5246 1893
rect 5258 1841 5310 1893
rect 6506 2675 6512 2701
rect 6512 2675 6546 2701
rect 6546 2675 6558 2701
rect 6506 2649 6558 2675
rect 6506 2629 6558 2637
rect 6506 2595 6512 2629
rect 6512 2595 6546 2629
rect 6546 2595 6558 2629
rect 6506 2585 6558 2595
rect 6648 2679 6700 2701
rect 6648 2649 6657 2679
rect 6657 2649 6691 2679
rect 6691 2649 6700 2679
rect 6648 2605 6700 2637
rect 6648 2585 6657 2605
rect 6657 2585 6691 2605
rect 6691 2585 6700 2605
rect 6274 1649 6326 1701
rect 6338 1649 6390 1701
rect 8137 2914 8189 2966
rect 8210 2914 8262 2966
rect 8283 2914 8335 2966
rect 8356 2914 8408 2966
rect 8429 2914 8481 2966
rect 8502 2914 8554 2966
rect 7216 2682 7268 2700
rect 7216 2648 7225 2682
rect 7225 2648 7259 2682
rect 7259 2648 7268 2682
rect 7216 2609 7268 2636
rect 7216 2584 7225 2609
rect 7225 2584 7259 2609
rect 7259 2584 7268 2609
rect 7361 2833 7370 2857
rect 7370 2833 7404 2857
rect 7404 2833 7413 2857
rect 7361 2805 7413 2833
rect 7361 2792 7413 2793
rect 7361 2758 7370 2792
rect 7370 2758 7404 2792
rect 7404 2758 7413 2792
rect 7361 2741 7413 2758
rect 7577 2683 7586 2700
rect 7586 2683 7620 2700
rect 7620 2683 7629 2700
rect 7577 2648 7629 2683
rect 7577 2608 7586 2630
rect 7586 2608 7620 2630
rect 7620 2608 7629 2630
rect 7577 2578 7629 2608
rect 7577 2533 7586 2560
rect 7586 2533 7620 2560
rect 7620 2533 7629 2560
rect 7577 2508 7629 2533
rect 7793 2833 7802 2857
rect 7802 2833 7836 2857
rect 7836 2833 7845 2857
rect 7793 2805 7845 2833
rect 7793 2792 7845 2793
rect 7793 2758 7802 2792
rect 7802 2758 7836 2792
rect 7836 2758 7845 2792
rect 7793 2741 7845 2758
rect 8009 2696 8061 2700
rect 8009 2662 8018 2696
rect 8018 2662 8052 2696
rect 8052 2662 8061 2696
rect 8009 2648 8061 2662
rect 8009 2624 8061 2630
rect 8009 2590 8018 2624
rect 8018 2590 8052 2624
rect 8052 2590 8061 2624
rect 8009 2578 8061 2590
rect 8009 2551 8061 2560
rect 8009 2517 8018 2551
rect 8018 2517 8052 2551
rect 8052 2517 8061 2551
rect 8009 2508 8061 2517
rect 8321 2683 8330 2700
rect 8330 2683 8364 2700
rect 8364 2683 8373 2700
rect 8321 2648 8373 2683
rect 8321 2608 8330 2630
rect 8330 2608 8364 2630
rect 8364 2608 8373 2630
rect 8321 2578 8373 2608
rect 8321 2533 8330 2560
rect 8330 2533 8364 2560
rect 8364 2533 8373 2560
rect 8321 2508 8373 2533
rect 8633 2683 8642 2700
rect 8642 2683 8676 2700
rect 8676 2683 8685 2700
rect 8633 2648 8685 2683
rect 8633 2608 8642 2630
rect 8642 2608 8676 2630
rect 8676 2608 8685 2630
rect 8633 2578 8685 2608
rect 8633 2533 8642 2560
rect 8642 2533 8676 2560
rect 8676 2533 8685 2560
rect 8633 2508 8685 2533
rect 8786 2679 8838 2700
rect 8786 2648 8795 2679
rect 8795 2648 8829 2679
rect 8829 2648 8838 2679
rect 8786 2605 8838 2630
rect 8786 2578 8795 2605
rect 8795 2578 8829 2605
rect 8829 2578 8838 2605
rect 8786 2531 8838 2560
rect 8786 2508 8795 2531
rect 8795 2508 8829 2531
rect 8829 2508 8838 2531
rect 8133 2028 8185 2080
rect 8197 2028 8249 2080
rect 8445 2028 8497 2080
rect 8509 2028 8561 2080
rect 5948 1489 6000 1541
rect 6012 1489 6064 1541
rect 7217 1649 7269 1701
rect 7281 1649 7333 1701
rect 3800 1104 3852 1156
rect 3864 1104 3916 1156
rect 1886 541 1938 593
rect 1886 474 1938 526
rect 3504 508 3556 560
rect 3248 458 3300 471
rect 3248 424 3257 458
rect 3257 424 3291 458
rect 3291 424 3300 458
rect 3248 419 3300 424
rect 3248 386 3300 407
rect 3248 355 3257 386
rect 3257 355 3291 386
rect 3291 355 3300 386
rect 3504 433 3556 485
rect 3504 358 3556 410
rect 3504 282 3556 334
rect 1586 178 1638 230
rect 1656 178 1708 230
rect 1726 178 1778 230
rect 1796 178 1848 230
rect 1866 178 1918 230
rect 1936 178 1988 230
rect 2006 178 2058 230
rect 2076 178 2128 230
rect 2146 178 2198 230
rect 2216 178 2268 230
rect 2285 178 2337 230
rect 1586 108 1638 160
rect 1656 108 1708 160
rect 1726 108 1778 160
rect 1796 108 1848 160
rect 1866 108 1918 160
rect 1936 108 1988 160
rect 2006 108 2058 160
rect 2076 108 2128 160
rect 2146 108 2198 160
rect 2216 108 2268 160
rect 2285 108 2337 160
rect 1586 82 1638 90
rect 1656 82 1708 90
rect 1726 82 1778 90
rect 1796 82 1848 90
rect 1866 82 1918 90
rect 1936 82 1988 90
rect 2006 82 2058 90
rect 2076 82 2128 90
rect 2146 82 2198 90
rect 2216 82 2268 90
rect 1586 48 1622 82
rect 1622 48 1638 82
rect 1656 48 1696 82
rect 1696 48 1708 82
rect 1726 48 1730 82
rect 1730 48 1770 82
rect 1770 48 1778 82
rect 1796 48 1804 82
rect 1804 48 1844 82
rect 1844 48 1848 82
rect 1866 48 1878 82
rect 1878 48 1918 82
rect 1936 48 1952 82
rect 1952 48 1988 82
rect 2006 48 2026 82
rect 2026 48 2058 82
rect 2076 48 2100 82
rect 2100 48 2128 82
rect 2146 48 2174 82
rect 2174 48 2198 82
rect 2216 48 2248 82
rect 2248 48 2268 82
rect 1586 38 1638 48
rect 1656 38 1708 48
rect 1726 38 1778 48
rect 1796 38 1848 48
rect 1866 38 1918 48
rect 1936 38 1988 48
rect 2006 38 2058 48
rect 2076 38 2128 48
rect 2146 38 2198 48
rect 2216 38 2268 48
rect 2285 82 2337 90
rect 2285 48 2287 82
rect 2287 48 2321 82
rect 2321 48 2337 82
rect 2285 38 2337 48
rect 2959 178 3011 230
rect 3029 178 3081 230
rect 3098 178 3150 230
rect 3167 178 3219 230
rect 3236 178 3288 230
rect 3305 178 3357 230
rect 3374 178 3426 230
rect 2959 108 3011 160
rect 3029 108 3081 160
rect 3098 108 3150 160
rect 3167 108 3219 160
rect 3236 108 3288 160
rect 3305 108 3357 160
rect 3374 108 3426 160
rect 2959 82 3011 90
rect 3029 82 3081 90
rect 3098 82 3150 90
rect 3167 82 3219 90
rect 3236 82 3288 90
rect 3305 82 3357 90
rect 3374 82 3426 90
rect 2959 48 2991 82
rect 2991 48 3011 82
rect 3029 48 3065 82
rect 3065 48 3081 82
rect 3098 48 3099 82
rect 3099 48 3139 82
rect 3139 48 3150 82
rect 3167 48 3173 82
rect 3173 48 3213 82
rect 3213 48 3219 82
rect 3236 48 3247 82
rect 3247 48 3288 82
rect 3305 48 3322 82
rect 3322 48 3357 82
rect 3374 48 3397 82
rect 3397 48 3426 82
rect 2959 38 3011 48
rect 3029 38 3081 48
rect 3098 38 3150 48
rect 3167 38 3219 48
rect 3236 38 3288 48
rect 3305 38 3357 48
rect 3374 38 3426 48
rect 3690 508 3742 560
rect 3754 508 3806 560
rect 3690 433 3742 485
rect 3754 433 3806 485
rect 3690 358 3742 410
rect 3754 358 3806 410
rect 3690 282 3742 334
rect 3754 282 3806 334
rect 3933 547 3942 560
rect 3942 547 3976 560
rect 3976 547 3985 560
rect 3933 508 3985 547
rect 3933 473 3942 484
rect 3942 473 3976 484
rect 3976 473 3985 484
rect 3933 433 3985 473
rect 3933 432 3942 433
rect 3942 432 3976 433
rect 3976 432 3985 433
rect 3933 399 3942 409
rect 3942 399 3976 409
rect 3976 399 3985 409
rect 3933 359 3985 399
rect 3933 357 3942 359
rect 3942 357 3976 359
rect 3976 357 3985 359
rect 3933 325 3942 334
rect 3942 325 3976 334
rect 3976 325 3985 334
rect 3933 285 3985 325
rect 3933 282 3942 285
rect 3942 282 3976 285
rect 3976 282 3985 285
rect 4039 938 4091 949
rect 4039 904 4048 938
rect 4048 904 4082 938
rect 4082 904 4091 938
rect 4039 897 4091 904
rect 4039 866 4091 873
rect 4039 832 4048 866
rect 4048 832 4082 866
rect 4082 832 4091 866
rect 4039 821 4091 832
rect 4039 794 4091 798
rect 4039 760 4048 794
rect 4048 760 4082 794
rect 4082 760 4091 794
rect 4039 746 4091 760
rect 4039 722 4091 723
rect 4039 688 4048 722
rect 4048 688 4082 722
rect 4082 688 4091 722
rect 4039 671 4091 688
rect 4145 543 4154 560
rect 4154 543 4188 560
rect 4188 543 4197 560
rect 4145 508 4197 543
rect 4145 470 4154 484
rect 4154 470 4188 484
rect 4188 470 4197 484
rect 4145 432 4197 470
rect 4145 397 4154 409
rect 4154 397 4188 409
rect 4188 397 4197 409
rect 4145 358 4197 397
rect 4145 357 4154 358
rect 4154 357 4188 358
rect 4188 357 4197 358
rect 4145 324 4154 334
rect 4154 324 4188 334
rect 4188 324 4197 334
rect 4145 285 4197 324
rect 4145 282 4154 285
rect 4154 282 4188 285
rect 4188 282 4197 285
rect 4251 938 4303 949
rect 4251 904 4260 938
rect 4260 904 4294 938
rect 4294 904 4303 938
rect 4251 897 4303 904
rect 4251 866 4303 873
rect 4251 832 4260 866
rect 4260 832 4294 866
rect 4294 832 4303 866
rect 4251 821 4303 832
rect 4251 794 4303 798
rect 4251 760 4260 794
rect 4260 760 4294 794
rect 4294 760 4303 794
rect 4251 746 4303 760
rect 4251 722 4303 723
rect 4251 688 4260 722
rect 4260 688 4294 722
rect 4294 688 4303 722
rect 4251 671 4303 688
rect 4357 543 4366 560
rect 4366 543 4400 560
rect 4400 543 4409 560
rect 4357 508 4409 543
rect 4357 470 4366 484
rect 4366 470 4400 484
rect 4400 470 4409 484
rect 4357 432 4409 470
rect 4357 397 4366 409
rect 4366 397 4400 409
rect 4400 397 4409 409
rect 4357 358 4409 397
rect 4357 357 4366 358
rect 4366 357 4400 358
rect 4400 357 4409 358
rect 4357 324 4366 334
rect 4366 324 4400 334
rect 4400 324 4409 334
rect 4357 285 4409 324
rect 4357 282 4366 285
rect 4366 282 4400 285
rect 4400 282 4409 285
rect 4463 938 4515 949
rect 4463 904 4472 938
rect 4472 904 4506 938
rect 4506 904 4515 938
rect 4463 897 4515 904
rect 4463 866 4515 873
rect 4463 832 4472 866
rect 4472 832 4506 866
rect 4506 832 4515 866
rect 4463 821 4515 832
rect 4463 794 4515 798
rect 4463 760 4472 794
rect 4472 760 4506 794
rect 4506 760 4515 794
rect 4463 746 4515 760
rect 4463 722 4515 723
rect 4463 688 4472 722
rect 4472 688 4506 722
rect 4506 688 4515 722
rect 4463 671 4515 688
rect 4569 543 4578 560
rect 4578 543 4612 560
rect 4612 543 4621 560
rect 4569 508 4621 543
rect 4569 470 4578 484
rect 4578 470 4612 484
rect 4612 470 4621 484
rect 4569 432 4621 470
rect 4569 397 4578 409
rect 4578 397 4612 409
rect 4612 397 4621 409
rect 4569 358 4621 397
rect 4569 357 4578 358
rect 4578 357 4612 358
rect 4612 357 4621 358
rect 4569 324 4578 334
rect 4578 324 4612 334
rect 4612 324 4621 334
rect 4569 285 4621 324
rect 4569 282 4578 285
rect 4578 282 4612 285
rect 4612 282 4621 285
rect 4675 938 4727 949
rect 4675 904 4684 938
rect 4684 904 4718 938
rect 4718 904 4727 938
rect 4675 897 4727 904
rect 4675 866 4727 873
rect 4675 832 4684 866
rect 4684 832 4718 866
rect 4718 832 4727 866
rect 4675 821 4727 832
rect 4675 794 4727 798
rect 4675 760 4684 794
rect 4684 760 4718 794
rect 4718 760 4727 794
rect 4675 746 4727 760
rect 4675 722 4727 723
rect 4675 688 4684 722
rect 4684 688 4718 722
rect 4718 688 4727 722
rect 4675 671 4727 688
rect 4781 543 4790 560
rect 4790 543 4824 560
rect 4824 543 4833 560
rect 4781 508 4833 543
rect 4781 470 4790 484
rect 4790 470 4824 484
rect 4824 470 4833 484
rect 4781 432 4833 470
rect 4781 397 4790 409
rect 4790 397 4824 409
rect 4824 397 4833 409
rect 4781 358 4833 397
rect 4781 357 4790 358
rect 4790 357 4824 358
rect 4824 357 4833 358
rect 4781 324 4790 334
rect 4790 324 4824 334
rect 4824 324 4833 334
rect 4781 285 4833 324
rect 4781 282 4790 285
rect 4790 282 4824 285
rect 4824 282 4833 285
rect 4887 938 4939 949
rect 4887 904 4896 938
rect 4896 904 4930 938
rect 4930 904 4939 938
rect 4887 897 4939 904
rect 4887 866 4939 873
rect 4887 832 4896 866
rect 4896 832 4930 866
rect 4930 832 4939 866
rect 4887 821 4939 832
rect 4887 794 4939 798
rect 4887 760 4896 794
rect 4896 760 4930 794
rect 4930 760 4939 794
rect 4887 746 4939 760
rect 4887 722 4939 723
rect 4887 688 4896 722
rect 4896 688 4930 722
rect 4930 688 4939 722
rect 4887 671 4939 688
rect 4993 543 5002 560
rect 5002 543 5036 560
rect 5036 543 5045 560
rect 4993 508 5045 543
rect 4993 470 5002 484
rect 5002 470 5036 484
rect 5036 470 5045 484
rect 4993 432 5045 470
rect 4993 397 5002 409
rect 5002 397 5036 409
rect 5036 397 5045 409
rect 4993 358 5045 397
rect 4993 357 5002 358
rect 5002 357 5036 358
rect 5036 357 5045 358
rect 4993 324 5002 334
rect 5002 324 5036 334
rect 5036 324 5045 334
rect 4993 285 5045 324
rect 4993 282 5002 285
rect 5002 282 5036 285
rect 5036 282 5045 285
rect 5099 938 5151 949
rect 5099 904 5108 938
rect 5108 904 5142 938
rect 5142 904 5151 938
rect 5099 897 5151 904
rect 5099 866 5151 873
rect 5099 832 5108 866
rect 5108 832 5142 866
rect 5142 832 5151 866
rect 5099 821 5151 832
rect 5099 794 5151 798
rect 5099 760 5108 794
rect 5108 760 5142 794
rect 5142 760 5151 794
rect 5099 746 5151 760
rect 5099 722 5151 723
rect 5099 688 5108 722
rect 5108 688 5142 722
rect 5142 688 5151 722
rect 5099 671 5151 688
rect 5205 543 5214 560
rect 5214 543 5248 560
rect 5248 543 5257 560
rect 5205 508 5257 543
rect 5205 470 5214 484
rect 5214 470 5248 484
rect 5248 470 5257 484
rect 5205 432 5257 470
rect 5205 397 5214 409
rect 5214 397 5248 409
rect 5248 397 5257 409
rect 5205 358 5257 397
rect 5205 357 5214 358
rect 5214 357 5248 358
rect 5248 357 5257 358
rect 5205 324 5214 334
rect 5214 324 5248 334
rect 5248 324 5257 334
rect 5205 285 5257 324
rect 5205 282 5214 285
rect 5214 282 5248 285
rect 5248 282 5257 285
rect 5311 938 5363 949
rect 5311 904 5320 938
rect 5320 904 5354 938
rect 5354 904 5363 938
rect 5311 897 5363 904
rect 5311 866 5363 873
rect 5311 832 5320 866
rect 5320 832 5354 866
rect 5354 832 5363 866
rect 5311 821 5363 832
rect 5311 794 5363 798
rect 5311 760 5320 794
rect 5320 760 5354 794
rect 5354 760 5363 794
rect 5311 746 5363 760
rect 5311 722 5363 723
rect 5311 688 5320 722
rect 5320 688 5354 722
rect 5354 688 5363 722
rect 5311 671 5363 688
rect 5417 543 5426 560
rect 5426 543 5460 560
rect 5460 543 5469 560
rect 5417 508 5469 543
rect 5417 470 5426 484
rect 5426 470 5460 484
rect 5460 470 5469 484
rect 5417 432 5469 470
rect 5417 397 5426 409
rect 5426 397 5460 409
rect 5460 397 5469 409
rect 5417 358 5469 397
rect 5417 357 5426 358
rect 5426 357 5460 358
rect 5460 357 5469 358
rect 5417 324 5426 334
rect 5426 324 5460 334
rect 5460 324 5469 334
rect 5417 285 5469 324
rect 5417 282 5426 285
rect 5426 282 5460 285
rect 5460 282 5469 285
rect 5523 938 5575 949
rect 5523 904 5532 938
rect 5532 904 5566 938
rect 5566 904 5575 938
rect 5523 897 5575 904
rect 5523 866 5575 873
rect 5523 832 5532 866
rect 5532 832 5566 866
rect 5566 832 5575 866
rect 5523 821 5575 832
rect 5523 794 5575 798
rect 5523 760 5532 794
rect 5532 760 5566 794
rect 5566 760 5575 794
rect 5523 746 5575 760
rect 5523 722 5575 723
rect 5523 688 5532 722
rect 5532 688 5566 722
rect 5566 688 5575 722
rect 5523 671 5575 688
rect 5629 543 5638 560
rect 5638 543 5672 560
rect 5672 543 5681 560
rect 5629 508 5681 543
rect 5629 470 5638 484
rect 5638 470 5672 484
rect 5672 470 5681 484
rect 5629 432 5681 470
rect 5629 397 5638 409
rect 5638 397 5672 409
rect 5672 397 5681 409
rect 5629 358 5681 397
rect 5629 357 5638 358
rect 5638 357 5672 358
rect 5672 357 5681 358
rect 5629 324 5638 334
rect 5638 324 5672 334
rect 5672 324 5681 334
rect 5629 285 5681 324
rect 5629 282 5638 285
rect 5638 282 5672 285
rect 5672 282 5681 285
rect 6726 996 6778 1048
rect 6726 932 6778 984
rect 7392 1569 7444 1621
rect 7456 1569 7508 1621
rect 9503 3245 9555 3297
rect 9639 3245 9691 3297
rect 9775 3245 9827 3297
rect 9911 3245 9963 3297
rect 10047 3245 10099 3297
rect 10183 3245 10235 3297
rect 10319 3245 10371 3297
rect 10455 3245 10507 3297
rect 10591 3245 10643 3297
rect 10727 3245 10779 3297
rect 10863 3245 10915 3297
rect 10999 3245 11051 3297
rect 11135 3245 11187 3297
rect 11271 3245 11323 3297
rect 11407 3245 11459 3297
rect 11542 3245 11594 3297
rect 11677 3245 11729 3297
rect 9503 3135 9555 3187
rect 9639 3135 9691 3187
rect 9775 3135 9827 3187
rect 9911 3135 9963 3187
rect 10047 3135 10099 3187
rect 10183 3135 10235 3187
rect 10319 3135 10371 3187
rect 10455 3135 10507 3187
rect 10591 3135 10643 3187
rect 10727 3135 10779 3187
rect 10863 3135 10915 3187
rect 10999 3135 11051 3187
rect 11135 3135 11187 3187
rect 11271 3135 11323 3187
rect 11407 3135 11459 3187
rect 11542 3135 11594 3187
rect 11677 3135 11729 3187
rect 7562 1489 7614 1541
rect 7626 1489 7678 1541
rect 9103 2811 9155 2863
rect 9181 2811 9233 2863
rect 9103 2735 9155 2787
rect 9181 2735 9233 2787
rect 9276 2422 9328 2474
rect 9340 2422 9392 2474
rect 5730 282 5782 334
rect 5730 218 5782 270
rect 6542 358 6594 364
rect 6542 324 6548 358
rect 6548 324 6582 358
rect 6582 324 6594 358
rect 6542 312 6594 324
rect 6542 286 6594 300
rect 6542 252 6548 286
rect 6548 252 6582 286
rect 6582 252 6594 286
rect 6791 283 6843 335
rect 6855 283 6907 335
rect 6542 248 6594 252
rect 7227 207 7236 224
rect 7236 207 7270 224
rect 7270 207 7279 224
rect 7227 172 7279 207
rect 7493 719 7545 736
rect 7493 685 7502 719
rect 7502 685 7536 719
rect 7536 685 7545 719
rect 7493 684 7545 685
rect 7493 644 7545 672
rect 7493 620 7502 644
rect 7502 620 7536 644
rect 7536 620 7545 644
rect 7227 132 7236 160
rect 7236 132 7270 160
rect 7270 132 7279 160
rect 7709 860 7761 892
rect 7709 840 7718 860
rect 7718 840 7752 860
rect 7752 840 7761 860
rect 7709 826 7718 828
rect 7718 826 7752 828
rect 7752 826 7761 828
rect 7709 786 7761 826
rect 7709 776 7718 786
rect 7718 776 7752 786
rect 7752 776 7761 786
rect 9402 2336 9454 2388
rect 9402 2272 9454 2324
rect 9795 2378 9803 2388
rect 9803 2378 9837 2388
rect 9837 2378 9847 2388
rect 9795 2338 9847 2378
rect 9795 2336 9803 2338
rect 9803 2336 9837 2338
rect 9837 2336 9847 2338
rect 9795 2304 9803 2324
rect 9803 2304 9837 2324
rect 9837 2304 9847 2324
rect 9795 2272 9847 2304
rect 10074 2440 10116 2474
rect 10116 2440 10126 2474
rect 10138 2440 10150 2474
rect 10150 2440 10190 2474
rect 10074 2422 10126 2440
rect 10138 2422 10190 2440
rect 10419 2209 10428 2231
rect 10428 2209 10462 2231
rect 10462 2209 10471 2231
rect 10419 2179 10471 2209
rect 10419 2132 10428 2166
rect 10428 2132 10462 2166
rect 10462 2132 10471 2166
rect 10419 2114 10471 2132
rect 10731 2697 10740 2700
rect 10740 2697 10774 2700
rect 10774 2697 10783 2700
rect 10731 2651 10783 2697
rect 10731 2648 10740 2651
rect 10740 2648 10774 2651
rect 10774 2648 10783 2651
rect 10731 2617 10740 2630
rect 10740 2617 10774 2630
rect 10774 2617 10783 2630
rect 10731 2578 10783 2617
rect 10731 2537 10740 2560
rect 10740 2537 10774 2560
rect 10774 2537 10783 2560
rect 10731 2508 10783 2537
rect 10698 1948 10750 2000
rect 10762 1948 10814 2000
rect 11043 2395 11052 2426
rect 11052 2395 11086 2426
rect 11086 2395 11095 2426
rect 11043 2374 11095 2395
rect 11043 2352 11095 2362
rect 11043 2318 11052 2352
rect 11052 2318 11086 2352
rect 11086 2318 11095 2352
rect 11043 2310 11095 2318
rect 11316 2782 11368 2794
rect 11380 2782 11432 2794
rect 11316 2748 11364 2782
rect 11364 2748 11368 2782
rect 11380 2748 11398 2782
rect 11398 2748 11432 2782
rect 11316 2742 11368 2748
rect 11380 2742 11432 2748
rect 10948 1873 11000 1882
rect 10948 1839 10954 1873
rect 10954 1839 10988 1873
rect 10988 1839 11000 1873
rect 10948 1830 11000 1839
rect 11012 1873 11064 1882
rect 11012 1839 11047 1873
rect 11047 1839 11064 1873
rect 11012 1830 11064 1839
rect 11922 3245 11974 3297
rect 11987 3245 12039 3297
rect 12052 3245 12104 3297
rect 12117 3245 12169 3297
rect 12182 3245 12234 3297
rect 12247 3245 12299 3297
rect 12312 3245 12364 3297
rect 12377 3245 12429 3297
rect 12442 3245 12494 3297
rect 12507 3245 12559 3297
rect 12572 3245 12624 3297
rect 12637 3245 12689 3297
rect 12702 3245 12754 3297
rect 12767 3245 12819 3297
rect 12832 3245 12884 3297
rect 12897 3245 12949 3297
rect 12962 3245 13014 3297
rect 13027 3245 13079 3297
rect 13092 3245 13144 3297
rect 13157 3245 13209 3297
rect 13222 3245 13274 3297
rect 13287 3245 13339 3297
rect 13352 3245 13404 3297
rect 13417 3245 13469 3297
rect 13482 3245 13534 3297
rect 13547 3245 13599 3297
rect 13612 3245 13664 3297
rect 13677 3245 13729 3297
rect 13742 3245 13794 3297
rect 13806 3245 13858 3297
rect 13870 3245 13922 3297
rect 13934 3245 13986 3297
rect 13998 3245 14050 3297
rect 14062 3245 14114 3297
rect 14126 3245 14178 3297
rect 14190 3245 14242 3297
rect 14254 3245 14306 3297
rect 14318 3245 14370 3297
rect 14382 3245 14434 3297
rect 14446 3245 14498 3297
rect 14510 3245 14562 3297
rect 14574 3245 14626 3297
rect 14638 3245 14690 3297
rect 14702 3245 14754 3297
rect 14766 3245 14818 3297
rect 14830 3245 14882 3297
rect 14894 3245 14946 3297
rect 14958 3245 15010 3297
rect 15022 3245 15074 3297
rect 15086 3245 15138 3297
rect 15150 3245 15202 3297
rect 15214 3245 15266 3297
rect 15278 3245 15330 3297
rect 15342 3245 15394 3297
rect 15406 3245 15458 3297
rect 15470 3245 15522 3297
rect 15534 3245 15586 3297
rect 15598 3245 15650 3297
rect 15662 3245 15714 3297
rect 15726 3245 15778 3297
rect 15790 3245 15842 3297
rect 15854 3245 15906 3297
rect 15918 3245 15970 3297
rect 15982 3245 16034 3297
rect 16046 3245 16098 3297
rect 16110 3245 16162 3297
rect 16174 3245 16226 3297
rect 16238 3245 16290 3297
rect 16302 3245 16354 3297
rect 16366 3245 16418 3297
rect 16430 3245 16482 3297
rect 16494 3245 16546 3297
rect 16558 3245 16610 3297
rect 16622 3245 16674 3297
rect 16686 3245 16738 3297
rect 16750 3245 16802 3297
rect 16814 3245 16866 3297
rect 16878 3245 16930 3297
rect 16942 3245 16994 3297
rect 17006 3245 17058 3297
rect 17070 3245 17122 3297
rect 11922 3135 11974 3187
rect 11987 3135 12039 3187
rect 12052 3135 12104 3187
rect 12117 3135 12169 3187
rect 12182 3135 12234 3187
rect 12247 3135 12299 3187
rect 12312 3135 12364 3187
rect 12377 3135 12429 3187
rect 12442 3135 12494 3187
rect 12507 3135 12559 3187
rect 12572 3135 12624 3187
rect 12637 3135 12689 3187
rect 12702 3135 12754 3187
rect 12767 3135 12819 3187
rect 12832 3135 12884 3187
rect 12897 3135 12949 3187
rect 12962 3135 13014 3187
rect 13027 3135 13079 3187
rect 13092 3135 13144 3187
rect 13157 3135 13209 3187
rect 13222 3135 13274 3187
rect 13287 3135 13339 3187
rect 13352 3135 13404 3187
rect 13417 3135 13469 3187
rect 13482 3135 13534 3187
rect 13547 3135 13599 3187
rect 13612 3135 13664 3187
rect 13677 3135 13729 3187
rect 13742 3135 13794 3187
rect 13806 3135 13858 3187
rect 13870 3135 13922 3187
rect 13934 3135 13986 3187
rect 13998 3135 14050 3187
rect 14062 3135 14114 3187
rect 14126 3135 14178 3187
rect 14190 3135 14242 3187
rect 14254 3135 14306 3187
rect 14318 3135 14370 3187
rect 14382 3135 14434 3187
rect 14446 3135 14498 3187
rect 14510 3135 14562 3187
rect 14574 3135 14626 3187
rect 14638 3135 14690 3187
rect 14702 3135 14754 3187
rect 14766 3135 14818 3187
rect 14830 3135 14882 3187
rect 14894 3135 14946 3187
rect 14958 3135 15010 3187
rect 15022 3135 15074 3187
rect 15086 3135 15138 3187
rect 15150 3135 15202 3187
rect 15214 3135 15266 3187
rect 15278 3135 15330 3187
rect 15342 3135 15394 3187
rect 15406 3135 15458 3187
rect 15470 3135 15522 3187
rect 15534 3135 15586 3187
rect 15598 3135 15650 3187
rect 15662 3135 15714 3187
rect 15726 3135 15778 3187
rect 15790 3135 15842 3187
rect 15854 3135 15906 3187
rect 15918 3135 15970 3187
rect 15982 3135 16034 3187
rect 16046 3135 16098 3187
rect 16110 3135 16162 3187
rect 16174 3135 16226 3187
rect 16238 3135 16290 3187
rect 16302 3135 16354 3187
rect 16366 3135 16418 3187
rect 16430 3135 16482 3187
rect 16494 3135 16546 3187
rect 16558 3135 16610 3187
rect 16622 3135 16674 3187
rect 16686 3135 16738 3187
rect 16750 3135 16802 3187
rect 16814 3135 16866 3187
rect 16878 3135 16930 3187
rect 16942 3135 16994 3187
rect 17006 3135 17058 3187
rect 17070 3135 17122 3187
rect 16837 2930 16889 2982
rect 16913 2930 16965 2982
rect 12225 2424 12277 2430
rect 12301 2424 12353 2430
rect 12225 2390 12252 2424
rect 12252 2390 12277 2424
rect 12301 2390 12325 2424
rect 12325 2390 12353 2424
rect 12225 2378 12277 2390
rect 12301 2378 12353 2390
rect 12225 2304 12277 2356
rect 12301 2304 12353 2356
rect 14040 2188 14092 2236
rect 14164 2188 14216 2236
rect 14040 2184 14064 2188
rect 14064 2184 14092 2188
rect 14040 2154 14064 2160
rect 14064 2154 14092 2160
rect 14164 2184 14176 2188
rect 14176 2184 14210 2188
rect 14210 2184 14216 2188
rect 14164 2154 14176 2160
rect 14176 2154 14210 2160
rect 14210 2154 14216 2160
rect 14040 2108 14092 2154
rect 14164 2108 14216 2154
rect 14260 2312 14266 2346
rect 14266 2312 14300 2346
rect 14300 2312 14312 2346
rect 14260 2294 14312 2312
rect 14260 2265 14312 2282
rect 14260 2231 14266 2265
rect 14266 2231 14300 2265
rect 14300 2231 14312 2265
rect 14260 2230 14312 2231
rect 14884 2841 14936 2893
rect 14972 2841 15024 2893
rect 14884 2778 14936 2825
rect 14972 2778 15024 2825
rect 16837 2838 16889 2890
rect 16913 2838 16965 2890
rect 14884 2773 14896 2778
rect 14896 2773 14930 2778
rect 14930 2773 14936 2778
rect 14972 2773 15004 2778
rect 15004 2773 15024 2778
rect 14884 2744 14896 2757
rect 14896 2744 14930 2757
rect 14930 2744 14936 2757
rect 14972 2744 15004 2757
rect 15004 2744 15024 2757
rect 14884 2705 14936 2744
rect 14972 2705 15024 2744
rect 14767 2312 14780 2346
rect 14780 2312 14814 2346
rect 14814 2312 14819 2346
rect 14767 2294 14819 2312
rect 14767 2265 14819 2282
rect 14767 2231 14780 2265
rect 14780 2231 14814 2265
rect 14814 2231 14819 2265
rect 14767 2230 14819 2231
rect 8186 1002 8238 1054
rect 8264 1002 8316 1054
rect 8186 926 8238 978
rect 8264 926 8316 978
rect 7925 719 7977 736
rect 7925 685 7934 719
rect 7934 685 7968 719
rect 7968 685 7977 719
rect 7925 684 7977 685
rect 7925 644 7977 672
rect 7925 620 7934 644
rect 7934 620 7968 644
rect 7968 620 7977 644
rect 8141 886 8193 892
rect 8141 852 8150 886
rect 8150 852 8184 886
rect 8184 852 8193 886
rect 8141 840 8193 852
rect 8141 810 8193 828
rect 8141 776 8150 810
rect 8150 776 8184 810
rect 8184 776 8193 810
rect 8573 860 8625 892
rect 8573 840 8582 860
rect 8582 840 8616 860
rect 8616 840 8625 860
rect 8573 826 8582 828
rect 8582 826 8616 828
rect 8616 826 8625 828
rect 8573 786 8625 826
rect 8573 776 8582 786
rect 8582 776 8616 786
rect 8616 776 8625 786
rect 8789 194 8841 224
rect 8789 172 8798 194
rect 8798 172 8832 194
rect 8832 172 8841 194
rect 7227 108 7279 132
rect 7227 78 7279 96
rect 8789 108 8841 160
rect 9005 860 9057 892
rect 9005 840 9014 860
rect 9014 840 9048 860
rect 9048 840 9057 860
rect 9005 826 9014 828
rect 9014 826 9048 828
rect 9048 826 9057 828
rect 9005 786 9057 826
rect 9005 776 9014 786
rect 9014 776 9048 786
rect 9048 776 9057 786
rect 9355 684 9407 736
rect 9355 620 9407 672
rect 9437 860 9489 892
rect 9437 840 9446 860
rect 9446 840 9480 860
rect 9480 840 9489 860
rect 9437 826 9446 828
rect 9446 826 9480 828
rect 9480 826 9489 828
rect 9437 786 9489 826
rect 9437 776 9446 786
rect 9446 776 9480 786
rect 9480 776 9489 786
rect 9221 194 9273 224
rect 9221 172 9230 194
rect 9230 172 9264 194
rect 9264 172 9273 194
rect 8789 78 8841 96
rect 9221 108 9273 160
rect 9699 1489 9751 1541
rect 9763 1489 9815 1541
rect 10520 1489 10572 1541
rect 10584 1489 10636 1541
rect 12182 1409 12234 1461
rect 12246 1409 12298 1461
rect 14462 1409 14514 1461
rect 14526 1409 14578 1461
rect 9571 523 9623 575
rect 9571 459 9623 511
rect 9653 194 9705 224
rect 9653 172 9662 194
rect 9662 172 9696 194
rect 9696 172 9705 194
rect 9221 78 9273 96
rect 9653 108 9705 160
rect 9869 869 9921 892
rect 9869 840 9878 869
rect 9878 840 9912 869
rect 9912 840 9921 869
rect 9869 794 9921 828
rect 9869 776 9878 794
rect 9878 776 9912 794
rect 9912 776 9921 794
rect 10085 1019 10137 1048
rect 10085 996 10094 1019
rect 10094 996 10128 1019
rect 10128 996 10137 1019
rect 10085 944 10137 984
rect 10085 932 10094 944
rect 10094 932 10128 944
rect 10128 932 10137 944
rect 10301 860 10353 892
rect 10301 840 10310 860
rect 10310 840 10344 860
rect 10344 840 10353 860
rect 10301 826 10310 828
rect 10310 826 10344 828
rect 10344 826 10353 828
rect 10301 786 10353 826
rect 10301 776 10310 786
rect 10310 776 10344 786
rect 10344 776 10353 786
rect 10517 1019 10569 1048
rect 10517 996 10526 1019
rect 10526 996 10560 1019
rect 10560 996 10569 1019
rect 10517 944 10569 984
rect 10517 932 10526 944
rect 10526 932 10560 944
rect 10560 932 10569 944
rect 10733 860 10785 892
rect 10733 840 10742 860
rect 10742 840 10776 860
rect 10776 840 10785 860
rect 10733 826 10742 828
rect 10742 826 10776 828
rect 10776 826 10785 828
rect 10733 786 10785 826
rect 10733 776 10742 786
rect 10742 776 10776 786
rect 10776 776 10785 786
rect 10949 1019 11001 1048
rect 10949 996 10958 1019
rect 10958 996 10992 1019
rect 10992 996 11001 1019
rect 10949 944 11001 984
rect 10949 932 10958 944
rect 10958 932 10992 944
rect 10992 932 11001 944
rect 11165 860 11217 892
rect 11165 840 11174 860
rect 11174 840 11208 860
rect 11208 840 11217 860
rect 11165 826 11174 828
rect 11174 826 11208 828
rect 11208 826 11217 828
rect 11165 786 11217 826
rect 11165 776 11174 786
rect 11174 776 11208 786
rect 11208 776 11217 786
rect 11381 1019 11433 1048
rect 11381 996 11390 1019
rect 11390 996 11424 1019
rect 11424 996 11433 1019
rect 11381 944 11433 984
rect 11381 932 11390 944
rect 11390 932 11424 944
rect 11424 932 11433 944
rect 11597 860 11649 892
rect 11597 840 11606 860
rect 11606 840 11640 860
rect 11640 840 11649 860
rect 11597 826 11606 828
rect 11606 826 11640 828
rect 11640 826 11649 828
rect 11597 786 11649 826
rect 11597 776 11606 786
rect 11606 776 11640 786
rect 11640 776 11649 786
rect 11814 1019 11866 1048
rect 11814 996 11823 1019
rect 11823 996 11857 1019
rect 11857 996 11866 1019
rect 11814 944 11866 984
rect 11814 932 11823 944
rect 11823 932 11857 944
rect 11857 932 11866 944
rect 12029 860 12081 892
rect 12029 840 12038 860
rect 12038 840 12072 860
rect 12072 840 12081 860
rect 12029 826 12038 828
rect 12038 826 12072 828
rect 12072 826 12081 828
rect 12029 786 12081 826
rect 12029 776 12038 786
rect 12038 776 12072 786
rect 12072 776 12081 786
rect 12245 1019 12297 1048
rect 12245 996 12254 1019
rect 12254 996 12288 1019
rect 12288 996 12297 1019
rect 12245 944 12297 984
rect 12245 932 12254 944
rect 12254 932 12288 944
rect 12288 932 12297 944
rect 12461 860 12513 892
rect 12461 840 12470 860
rect 12470 840 12504 860
rect 12504 840 12513 860
rect 12461 826 12470 828
rect 12470 826 12504 828
rect 12504 826 12513 828
rect 12461 786 12513 826
rect 12461 776 12470 786
rect 12470 776 12504 786
rect 12504 776 12513 786
rect 12677 194 12729 224
rect 12677 172 12686 194
rect 12686 172 12720 194
rect 12720 172 12729 194
rect 9653 78 9705 96
rect 12677 108 12729 160
rect 12893 860 12945 892
rect 12893 840 12902 860
rect 12902 840 12936 860
rect 12936 840 12945 860
rect 12893 826 12902 828
rect 12902 826 12936 828
rect 12936 826 12945 828
rect 12893 786 12945 826
rect 12893 776 12902 786
rect 12902 776 12936 786
rect 12936 776 12945 786
rect 13109 194 13161 224
rect 13109 172 13118 194
rect 13118 172 13152 194
rect 13152 172 13161 194
rect 12677 78 12729 96
rect 13109 108 13161 160
rect 13325 860 13377 892
rect 13325 840 13334 860
rect 13334 840 13368 860
rect 13368 840 13377 860
rect 13325 826 13334 828
rect 13334 826 13368 828
rect 13368 826 13377 828
rect 13325 786 13377 826
rect 13325 776 13334 786
rect 13334 776 13368 786
rect 13368 776 13377 786
rect 13541 194 13593 224
rect 13541 172 13550 194
rect 13550 172 13584 194
rect 13584 172 13593 194
rect 13109 78 13161 96
rect 13541 108 13593 160
rect 13757 860 13809 892
rect 13757 840 13766 860
rect 13766 840 13800 860
rect 13800 840 13809 860
rect 13757 826 13766 828
rect 13766 826 13800 828
rect 13800 826 13809 828
rect 13757 786 13809 826
rect 13757 776 13766 786
rect 13766 776 13800 786
rect 13800 776 13809 786
rect 13973 194 14025 224
rect 13973 172 13982 194
rect 13982 172 14016 194
rect 14016 172 14025 194
rect 13541 78 13593 96
rect 13973 108 14025 160
rect 14189 860 14241 892
rect 14189 840 14198 860
rect 14198 840 14232 860
rect 14232 840 14241 860
rect 14189 826 14198 828
rect 14198 826 14232 828
rect 14232 826 14241 828
rect 14189 786 14241 826
rect 14189 776 14198 786
rect 14198 776 14232 786
rect 14232 776 14241 786
rect 14405 194 14457 224
rect 14405 172 14414 194
rect 14414 172 14448 194
rect 14448 172 14457 194
rect 13973 78 14025 96
rect 14405 108 14457 160
rect 14621 860 14673 892
rect 14621 840 14630 860
rect 14630 840 14664 860
rect 14664 840 14673 860
rect 14621 826 14630 828
rect 14630 826 14664 828
rect 14664 826 14673 828
rect 14621 786 14673 826
rect 14621 776 14630 786
rect 14630 776 14664 786
rect 14664 776 14673 786
rect 14837 194 14889 224
rect 14837 172 14846 194
rect 14846 172 14880 194
rect 14880 172 14889 194
rect 14405 78 14457 96
rect 14837 108 14889 160
rect 15053 860 15105 892
rect 15053 840 15062 860
rect 15062 840 15096 860
rect 15096 840 15105 860
rect 15053 826 15062 828
rect 15062 826 15096 828
rect 15096 826 15105 828
rect 15053 786 15105 826
rect 15053 776 15062 786
rect 15062 776 15096 786
rect 15096 776 15105 786
rect 15418 172 15470 224
rect 14837 78 14889 96
rect 15418 108 15470 160
rect 15529 310 15538 332
rect 15538 310 15572 332
rect 15572 310 15581 332
rect 15529 280 15581 310
rect 15529 235 15538 267
rect 15538 235 15572 267
rect 15572 235 15581 267
rect 15529 215 15581 235
rect 15529 194 15581 202
rect 15529 160 15538 194
rect 15538 160 15572 194
rect 15572 160 15581 194
rect 15529 150 15581 160
rect 15961 310 15970 332
rect 15970 310 16004 332
rect 16004 310 16013 332
rect 15961 280 16013 310
rect 15961 235 15970 267
rect 15970 235 16004 267
rect 16004 235 16013 267
rect 15961 215 16013 235
rect 15961 194 16013 202
rect 15961 160 15970 194
rect 15970 160 16004 194
rect 16004 160 16013 194
rect 15961 150 16013 160
rect 15418 78 15470 96
rect 7227 44 7237 78
rect 7237 44 7276 78
rect 7276 44 7279 78
rect 8789 44 8809 78
rect 8809 44 8841 78
rect 9221 44 9247 78
rect 9247 44 9273 78
rect 9653 44 9685 78
rect 9685 44 9705 78
rect 12677 44 12711 78
rect 12711 44 12729 78
rect 13109 44 13143 78
rect 13143 44 13161 78
rect 13541 44 13575 78
rect 13575 44 13593 78
rect 13973 44 14007 78
rect 14007 44 14025 78
rect 14405 44 14439 78
rect 14439 44 14457 78
rect 14837 44 14871 78
rect 14871 44 14889 78
rect 15418 44 15447 78
rect 15447 44 15470 78
rect 3041 -885 3093 -833
rect 3131 -885 3183 -833
rect 15335 -885 15387 -833
rect 15399 -885 15451 -833
<< metal2 >>
rect 92 3297 17128 3318
rect 92 3245 9503 3297
rect 9555 3245 9639 3297
rect 9691 3245 9775 3297
rect 9827 3245 9911 3297
rect 9963 3245 10047 3297
rect 10099 3245 10183 3297
rect 10235 3245 10319 3297
rect 10371 3245 10455 3297
rect 10507 3245 10591 3297
rect 10643 3245 10727 3297
rect 10779 3245 10863 3297
rect 10915 3245 10999 3297
rect 11051 3245 11135 3297
rect 11187 3245 11271 3297
rect 11323 3245 11407 3297
rect 11459 3245 11542 3297
rect 11594 3245 11677 3297
rect 11729 3245 11922 3297
rect 11974 3245 11987 3297
rect 12039 3245 12052 3297
rect 12104 3245 12117 3297
rect 12169 3245 12182 3297
rect 12234 3245 12247 3297
rect 12299 3245 12312 3297
rect 12364 3245 12377 3297
rect 12429 3245 12442 3297
rect 12494 3245 12507 3297
rect 12559 3245 12572 3297
rect 12624 3245 12637 3297
rect 12689 3245 12702 3297
rect 12754 3245 12767 3297
rect 12819 3245 12832 3297
rect 12884 3245 12897 3297
rect 12949 3245 12962 3297
rect 13014 3245 13027 3297
rect 13079 3245 13092 3297
rect 13144 3245 13157 3297
rect 13209 3245 13222 3297
rect 13274 3245 13287 3297
rect 13339 3245 13352 3297
rect 13404 3245 13417 3297
rect 13469 3245 13482 3297
rect 13534 3245 13547 3297
rect 13599 3245 13612 3297
rect 13664 3245 13677 3297
rect 13729 3245 13742 3297
rect 13794 3245 13806 3297
rect 13858 3245 13870 3297
rect 13922 3245 13934 3297
rect 13986 3245 13998 3297
rect 14050 3245 14062 3297
rect 14114 3245 14126 3297
rect 14178 3245 14190 3297
rect 14242 3245 14254 3297
rect 14306 3245 14318 3297
rect 14370 3245 14382 3297
rect 14434 3245 14446 3297
rect 14498 3245 14510 3297
rect 14562 3245 14574 3297
rect 14626 3245 14638 3297
rect 14690 3245 14702 3297
rect 14754 3245 14766 3297
rect 14818 3245 14830 3297
rect 14882 3245 14894 3297
rect 14946 3245 14958 3297
rect 15010 3245 15022 3297
rect 15074 3245 15086 3297
rect 15138 3245 15150 3297
rect 15202 3245 15214 3297
rect 15266 3245 15278 3297
rect 15330 3245 15342 3297
rect 15394 3245 15406 3297
rect 15458 3245 15470 3297
rect 15522 3245 15534 3297
rect 15586 3245 15598 3297
rect 15650 3245 15662 3297
rect 15714 3245 15726 3297
rect 15778 3245 15790 3297
rect 15842 3245 15854 3297
rect 15906 3245 15918 3297
rect 15970 3245 15982 3297
rect 16034 3245 16046 3297
rect 16098 3245 16110 3297
rect 16162 3245 16174 3297
rect 16226 3245 16238 3297
rect 16290 3245 16302 3297
rect 16354 3245 16366 3297
rect 16418 3245 16430 3297
rect 16482 3245 16494 3297
rect 16546 3245 16558 3297
rect 16610 3245 16622 3297
rect 16674 3245 16686 3297
rect 16738 3245 16750 3297
rect 16802 3245 16814 3297
rect 16866 3245 16878 3297
rect 16930 3245 16942 3297
rect 16994 3245 17006 3297
rect 17058 3245 17070 3297
rect 17122 3245 17128 3297
rect 92 3187 17128 3245
rect 92 3171 9503 3187
rect 92 3135 3739 3171
tri 3739 3135 3775 3171 nw
tri 4146 3135 4182 3171 ne
rect 4182 3135 9503 3171
rect 9555 3135 9639 3187
rect 9691 3135 9775 3187
rect 9827 3135 9911 3187
rect 9963 3135 10047 3187
rect 10099 3135 10183 3187
rect 10235 3135 10319 3187
rect 10371 3135 10455 3187
rect 10507 3135 10591 3187
rect 10643 3135 10727 3187
rect 10779 3135 10863 3187
rect 10915 3135 10999 3187
rect 11051 3135 11135 3187
rect 11187 3135 11271 3187
rect 11323 3135 11407 3187
rect 11459 3135 11542 3187
rect 11594 3135 11677 3187
rect 11729 3135 11922 3187
rect 11974 3135 11987 3187
rect 12039 3135 12052 3187
rect 12104 3135 12117 3187
rect 12169 3135 12182 3187
rect 12234 3135 12247 3187
rect 12299 3135 12312 3187
rect 12364 3135 12377 3187
rect 12429 3135 12442 3187
rect 12494 3135 12507 3187
rect 12559 3135 12572 3187
rect 12624 3135 12637 3187
rect 12689 3135 12702 3187
rect 12754 3135 12767 3187
rect 12819 3135 12832 3187
rect 12884 3135 12897 3187
rect 12949 3135 12962 3187
rect 13014 3135 13027 3187
rect 13079 3135 13092 3187
rect 13144 3135 13157 3187
rect 13209 3135 13222 3187
rect 13274 3135 13287 3187
rect 13339 3135 13352 3187
rect 13404 3135 13417 3187
rect 13469 3135 13482 3187
rect 13534 3135 13547 3187
rect 13599 3135 13612 3187
rect 13664 3135 13677 3187
rect 13729 3135 13742 3187
rect 13794 3135 13806 3187
rect 13858 3135 13870 3187
rect 13922 3135 13934 3187
rect 13986 3135 13998 3187
rect 14050 3135 14062 3187
rect 14114 3135 14126 3187
rect 14178 3135 14190 3187
rect 14242 3135 14254 3187
rect 14306 3135 14318 3187
rect 14370 3135 14382 3187
rect 14434 3135 14446 3187
rect 14498 3135 14510 3187
rect 14562 3135 14574 3187
rect 14626 3135 14638 3187
rect 14690 3135 14702 3187
rect 14754 3135 14766 3187
rect 14818 3135 14830 3187
rect 14882 3135 14894 3187
rect 14946 3135 14958 3187
rect 15010 3135 15022 3187
rect 15074 3135 15086 3187
rect 15138 3135 15150 3187
rect 15202 3135 15214 3187
rect 15266 3135 15278 3187
rect 15330 3135 15342 3187
rect 15394 3135 15406 3187
rect 15458 3135 15470 3187
rect 15522 3135 15534 3187
rect 15586 3135 15598 3187
rect 15650 3135 15662 3187
rect 15714 3135 15726 3187
rect 15778 3135 15790 3187
rect 15842 3135 15854 3187
rect 15906 3135 15918 3187
rect 15970 3135 15982 3187
rect 16034 3135 16046 3187
rect 16098 3135 16110 3187
rect 16162 3135 16174 3187
rect 16226 3135 16238 3187
rect 16290 3135 16302 3187
rect 16354 3135 16366 3187
rect 16418 3135 16430 3187
rect 16482 3135 16494 3187
rect 16546 3135 16558 3187
rect 16610 3135 16622 3187
rect 16674 3135 16686 3187
rect 16738 3135 16750 3187
rect 16802 3135 16814 3187
rect 16866 3135 16878 3187
rect 16930 3135 16942 3187
rect 16994 3135 17006 3187
rect 17058 3135 17070 3187
rect 17122 3135 17128 3187
rect 92 3118 3722 3135
tri 3722 3118 3739 3135 nw
tri 4182 3118 4199 3135 ne
rect 4199 3118 17128 3135
rect -2286 3082 -61 3085
rect -2286 3030 -183 3082
rect -131 3030 -119 3082
rect -67 3030 -61 3082
rect -2286 3025 -61 3030
rect -2286 3019 -2118 3025
tri -2118 3019 -2112 3025 nw
rect -2286 3013 -2124 3019
tri -2124 3013 -2118 3019 nw
rect 806 3013 3713 3019
tri 3713 3013 3719 3019 sw
rect -2286 2944 -2170 3013
tri -2170 2967 -2124 3013 nw
rect 806 2978 3719 3013
tri 3719 2978 3754 3013 sw
rect 806 2943 3754 2978
rect 806 2891 833 2943
rect 885 2891 897 2943
rect 949 2891 3754 2943
rect 4178 2983 4578 3019
rect 4178 2927 4187 2983
rect 4243 2927 4268 2983
rect 4324 2927 4349 2983
rect 4405 2927 4431 2983
rect 4487 2927 4513 2983
rect 4569 2927 4578 2983
rect 4178 2891 4578 2927
rect 5196 3013 5748 3019
rect 5196 2961 5221 3013
rect 5273 2961 5748 3013
rect 5196 2949 5748 2961
rect 5196 2897 5221 2949
rect 5273 2943 5748 2949
rect 5273 2897 5626 2943
rect 5196 2891 5626 2897
rect 5678 2891 5690 2943
rect 5742 2891 5748 2943
rect 6780 3007 8571 3064
rect 6780 2951 6793 3007
rect 6849 2951 6888 3007
rect 6944 2951 6984 3007
rect 7040 2951 7080 3007
rect 7136 2966 8571 3007
rect 7136 2951 8137 2966
rect 6780 2914 8137 2951
rect 8189 2914 8210 2966
rect 8262 2914 8283 2966
rect 8335 2914 8356 2966
rect 8408 2914 8429 2966
rect 8481 2914 8502 2966
rect 8554 2914 8571 2966
rect 6780 2891 8571 2914
rect 11310 2982 16965 3086
rect 11310 2930 16837 2982
rect 16889 2930 16913 2982
rect 11310 2927 16965 2930
rect 11310 2899 11444 2927
tri 11444 2899 11472 2927 nw
tri 16803 2899 16831 2927 ne
rect 16831 2899 16965 2927
tri 3574 2863 3602 2891 ne
rect 3602 2863 3754 2891
tri 3602 2857 3608 2863 ne
rect 3608 2857 3754 2863
tri 3608 2855 3610 2857 ne
rect 1289 2843 3569 2849
rect 1341 2791 1601 2843
rect 1653 2791 1913 2843
rect 1965 2838 3569 2843
rect 1965 2791 3345 2838
rect 1289 2782 3345 2791
rect 3401 2782 3425 2838
rect 3481 2782 3505 2838
rect 3561 2782 3569 2838
rect 1289 2778 3569 2782
rect 1341 2726 1601 2778
rect 1653 2726 1913 2778
rect 1965 2747 3569 2778
rect 1965 2726 3345 2747
rect 1289 2713 3345 2726
rect 1341 2661 1601 2713
rect 1653 2661 1913 2713
rect 1965 2691 3345 2713
rect 3401 2691 3425 2747
rect 3481 2691 3505 2747
rect 3561 2691 3569 2747
rect 1965 2661 3569 2691
rect 1289 2655 3569 2661
rect 1289 2648 3345 2655
rect 1341 2596 1601 2648
rect 1653 2596 1913 2648
rect 1965 2599 3345 2648
rect 3401 2599 3425 2655
rect 3481 2599 3505 2655
rect 3561 2599 3569 2655
rect 3610 2741 3754 2857
rect 4292 2857 9103 2863
rect 4344 2805 6021 2857
rect 6073 2805 6424 2857
rect 6476 2805 7361 2857
rect 7413 2805 7793 2857
rect 7845 2811 9103 2857
rect 9155 2811 9181 2863
rect 9233 2811 9239 2863
rect 7845 2805 9239 2811
rect 4292 2793 9239 2805
tri 3754 2741 3760 2747 sw
rect 4344 2741 6021 2793
rect 6073 2741 6424 2793
rect 6476 2741 7361 2793
rect 7413 2741 7793 2793
rect 7845 2787 9239 2793
rect 7845 2741 9103 2787
rect 3610 2735 3760 2741
tri 3760 2735 3766 2741 sw
rect 4292 2735 9103 2741
rect 9155 2735 9181 2787
rect 9233 2735 9239 2787
rect 11310 2794 11438 2899
tri 11438 2893 11444 2899 nw
rect 11939 2893 15024 2899
tri 16831 2893 16837 2899 ne
rect 11310 2742 11316 2794
rect 11368 2742 11380 2794
rect 11432 2742 11438 2794
rect 11939 2841 14884 2893
rect 14936 2841 14972 2893
rect 11939 2825 15024 2841
rect 16837 2890 16965 2899
rect 16889 2838 16913 2890
rect 16837 2832 16965 2838
rect 11939 2773 14884 2825
rect 14936 2773 14972 2825
rect 11939 2757 15024 2773
tri 11934 2735 11939 2740 se
rect 11939 2735 14884 2757
rect 3610 2707 3766 2735
tri 3766 2707 3794 2735 sw
tri 11906 2707 11934 2735 se
rect 11934 2707 14884 2735
rect 3610 2701 5300 2707
rect 3610 2664 5221 2701
tri 3610 2649 3625 2664 ne
rect 3625 2649 5221 2664
rect 5273 2649 5300 2701
tri 3625 2648 3626 2649 ne
rect 3626 2648 5300 2649
tri 3626 2637 3637 2648 ne
rect 3637 2637 5300 2648
rect 1965 2596 3569 2599
rect 1289 2590 3569 2596
tri 3637 2590 3684 2637 ne
rect 3684 2590 5221 2637
tri 3684 2585 3689 2590 ne
rect 3689 2585 5221 2590
rect 5273 2585 5300 2637
tri 3689 2584 3690 2585 ne
rect 3690 2584 5300 2585
tri 3690 2579 3695 2584 ne
rect 3695 2579 5300 2584
rect 5348 2701 6700 2707
tri 11905 2706 11906 2707 se
rect 11906 2706 14884 2707
rect 5400 2649 5493 2701
rect 5545 2649 5803 2701
rect 5855 2649 6237 2701
rect 6289 2649 6506 2701
rect 6558 2649 6648 2701
rect 5348 2637 6700 2649
rect 5400 2585 5493 2637
rect 5545 2585 5803 2637
rect 5855 2585 6237 2637
rect 6289 2585 6506 2637
rect 6558 2585 6648 2637
rect 5348 2579 6700 2585
rect 7199 2705 14884 2706
rect 14936 2705 14972 2757
rect 7199 2700 15024 2705
rect 7199 2648 7216 2700
rect 7268 2648 7577 2700
rect 7629 2648 8009 2700
rect 8061 2648 8321 2700
rect 8373 2648 8633 2700
rect 8685 2648 8786 2700
rect 8838 2648 10731 2700
rect 10783 2699 15024 2700
rect 10783 2648 12140 2699
tri 12140 2665 12174 2699 nw
rect 7199 2636 12140 2648
rect 7199 2584 7216 2636
rect 7268 2630 12140 2636
rect 7268 2584 7577 2630
rect 7199 2578 7577 2584
rect 7629 2578 8009 2630
rect 8061 2578 8321 2630
rect 8373 2578 8633 2630
rect 8685 2578 8786 2630
rect 8838 2578 10731 2630
rect 10783 2578 12140 2630
rect 7199 2560 12140 2578
rect 408 2544 6718 2550
rect 408 2492 711 2544
rect 763 2492 1023 2544
rect 1075 2492 2849 2544
rect 2901 2492 3161 2544
rect 3213 2502 6718 2544
rect 7199 2508 7577 2560
rect 7629 2508 8009 2560
rect 8061 2508 8321 2560
rect 8373 2508 8633 2560
rect 8685 2508 8786 2560
rect 8838 2508 10731 2560
rect 10783 2508 12140 2560
tri 6718 2502 6724 2508 sw
rect 7199 2502 12140 2508
rect 3213 2492 6724 2502
rect 408 2480 6724 2492
rect 408 2428 711 2480
rect 763 2428 1023 2480
rect 1075 2428 2849 2480
rect 2901 2428 3161 2480
rect 3213 2474 6724 2480
tri 6724 2474 6752 2502 sw
rect 3213 2428 9276 2474
rect 408 2422 9276 2428
rect 9328 2422 9340 2474
rect 9392 2422 10074 2474
rect 10126 2422 10138 2474
rect 10190 2422 10196 2474
rect 11043 2430 12359 2432
rect 11043 2426 12225 2430
rect 2208 2388 9847 2394
rect 2208 2336 2225 2388
rect 2277 2336 2537 2388
rect 2589 2336 9402 2388
rect 9454 2336 9795 2388
rect 2208 2324 9847 2336
rect 2208 2272 2225 2324
rect 2277 2272 2537 2324
rect 2589 2272 9402 2324
rect 9454 2272 9795 2324
rect 11095 2378 12225 2426
rect 12277 2378 12301 2430
rect 12353 2378 12359 2430
rect 11095 2374 12359 2378
rect 11043 2362 12359 2374
rect 11095 2356 12359 2362
rect 11095 2310 12225 2356
rect 11043 2304 12225 2310
rect 12277 2304 12301 2356
rect 12353 2304 12359 2356
tri 14238 2346 14244 2352 se
rect 14244 2346 17247 2352
tri 14233 2341 14238 2346 se
rect 14238 2341 14260 2346
rect 13546 2294 14260 2341
rect 14312 2294 14767 2346
rect 14819 2294 17247 2346
rect 13546 2285 17247 2294
tri 14233 2282 14236 2285 ne
rect 14236 2282 17247 2285
rect 2208 2266 9847 2272
tri 14236 2266 14252 2282 ne
rect 14252 2266 14260 2282
tri 14252 2258 14260 2266 ne
rect 196 2236 14222 2237
rect 196 2231 14040 2236
rect 196 2179 424 2231
rect 476 2179 1133 2231
rect 1185 2179 1445 2231
rect 1497 2179 1757 2231
rect 1809 2179 2069 2231
rect 2121 2179 2381 2231
rect 2433 2179 2693 2231
rect 2745 2179 3005 2231
rect 3057 2179 3317 2231
rect 3369 2179 3629 2231
rect 3681 2179 3941 2231
rect 3993 2179 4361 2231
rect 4413 2179 4664 2231
rect 4716 2179 10419 2231
rect 10471 2184 14040 2231
rect 14092 2184 14164 2236
rect 14216 2184 14222 2236
rect 14312 2230 14767 2282
rect 14819 2230 17247 2282
rect 14260 2224 17247 2230
rect 10471 2179 14222 2184
rect 196 2166 14222 2179
rect 196 2114 424 2166
rect 476 2114 1133 2166
rect 1185 2114 1445 2166
rect 1497 2114 1757 2166
rect 1809 2114 2069 2166
rect 2121 2114 2381 2166
rect 2433 2114 2693 2166
rect 2745 2114 3005 2166
rect 3057 2114 3317 2166
rect 3369 2114 3629 2166
rect 3681 2114 3941 2166
rect 3993 2114 4361 2166
rect 4413 2114 4664 2166
rect 4716 2114 10419 2166
rect 10471 2160 14222 2166
rect 10471 2114 14040 2160
rect 196 2108 14040 2114
rect 14092 2108 14164 2160
rect 14216 2108 14222 2160
rect 75 2028 676 2080
rect 728 2028 740 2080
rect 792 2028 1417 2080
rect 1469 2028 1481 2080
rect 1533 2028 5619 2080
rect 5671 2028 5683 2080
rect 5735 2028 8133 2080
rect 8185 2028 8197 2080
rect 8249 2028 8445 2080
rect 8497 2028 8509 2080
rect 8561 2028 8567 2080
rect 75 1994 10698 2000
rect 75 1948 4787 1994
tri 4753 1942 4759 1948 ne
rect 4759 1942 4787 1948
rect 4839 1948 10698 1994
rect 10750 1948 10762 2000
rect 10814 1948 10878 2000
tri 4759 1930 4771 1942 ne
rect 4771 1930 4839 1942
tri 4771 1914 4787 1930 ne
rect 75 1830 2225 1882
rect 2277 1830 2289 1882
rect 2341 1830 2347 1882
rect 2750 1830 2756 1882
rect 2808 1830 2820 1882
rect 2872 1830 2878 1882
tri 4839 1914 4873 1948 nw
rect 4787 1872 4839 1878
rect 5188 1893 7142 1914
tri 2716 1781 2750 1815 se
rect 2750 1810 2878 1830
rect 5188 1841 5194 1893
rect 5246 1841 5258 1893
rect 5310 1890 7142 1893
rect 5310 1841 6795 1890
rect 5188 1834 6795 1841
rect 6851 1834 6936 1890
rect 6992 1834 7077 1890
rect 7133 1834 7142 1890
tri 2878 1810 2883 1815 sw
rect 5188 1810 7142 1834
rect 10942 1830 10948 1882
rect 11000 1830 11012 1882
rect 11064 1830 11070 1882
tri 10937 1810 10942 1815 se
rect 10942 1810 11070 1830
rect 2750 1781 2883 1810
tri 2883 1781 2912 1810 sw
tri 10908 1781 10937 1810 se
rect 10937 1781 11070 1810
rect 75 1729 827 1781
rect 879 1729 891 1781
rect 943 1729 11070 1781
rect 3972 1649 3978 1701
rect 4030 1649 4042 1701
rect 4094 1649 6274 1701
rect 6326 1649 6338 1701
rect 6390 1649 7217 1701
rect 7269 1649 7281 1701
rect 7333 1649 11070 1701
rect 75 1569 3556 1621
rect 3608 1569 3620 1621
rect 3672 1569 7392 1621
rect 7444 1569 7456 1621
rect 7508 1569 11070 1621
rect 14 1489 5948 1541
rect 6000 1489 6012 1541
rect 6064 1489 7562 1541
rect 7614 1489 7626 1541
rect 7678 1489 9699 1541
rect 9751 1489 9763 1541
rect 9815 1489 10520 1541
rect 10572 1489 10584 1541
rect 10636 1489 10642 1541
rect 14 1409 12182 1461
rect 12234 1409 12246 1461
rect 12298 1409 14462 1461
rect 14514 1409 14526 1461
rect 14578 1409 15032 1461
rect 2202 1104 3800 1156
rect 3852 1104 3864 1156
rect 3916 1104 3922 1156
tri 2172 762 2202 792 se
rect 2202 762 2244 1104
tri 2244 1071 2277 1104 nw
rect 6708 1048 8186 1054
rect 6708 996 6726 1048
rect 6778 1002 8186 1048
rect 8238 1002 8264 1054
rect 8316 1048 12299 1054
rect 8316 1002 10085 1048
rect 6778 996 10085 1002
rect 10137 996 10517 1048
rect 10569 996 10949 1048
rect 11001 996 11381 1048
rect 11433 996 11814 1048
rect 11866 996 12245 1048
rect 12297 996 12299 1048
rect 6708 984 12299 996
rect 1886 710 2244 762
rect 3329 949 4731 955
rect 3329 946 4039 949
rect 3329 890 3345 946
rect 3401 890 3425 946
rect 3481 890 3505 946
rect 3561 897 4039 946
rect 4091 897 4251 949
rect 4303 897 4463 949
rect 4515 897 4675 949
rect 4727 897 4731 949
rect 3561 890 4731 897
rect 3329 873 4731 890
rect 3329 838 4039 873
rect 3329 782 3345 838
rect 3401 782 3425 838
rect 3481 782 3505 838
rect 3561 821 4039 838
rect 4091 821 4251 873
rect 4303 821 4463 873
rect 4515 821 4675 873
rect 4727 821 4731 873
rect 3561 798 4731 821
rect 3561 782 4039 798
rect 3329 746 4039 782
rect 4091 746 4251 798
rect 4303 746 4463 798
rect 4515 746 4675 798
rect 4727 746 4731 798
rect 3329 730 4731 746
rect 1886 593 1938 710
tri 1938 682 1966 710 nw
rect 3329 674 3345 730
rect 3401 674 3425 730
rect 3481 674 3505 730
rect 3561 723 4731 730
rect 3561 674 4039 723
rect 3329 671 4039 674
rect 4091 671 4251 723
rect 4303 671 4463 723
rect 4515 671 4675 723
rect 4727 671 4731 723
rect 3329 665 4731 671
rect 4883 949 5937 955
rect 4883 897 4887 949
rect 4939 897 5099 949
rect 5151 897 5311 949
rect 5363 897 5523 949
rect 5575 932 5937 949
tri 5937 932 5960 955 sw
rect 6708 932 6726 984
rect 6778 978 10085 984
rect 6778 932 8186 978
rect 5575 926 5960 932
tri 5960 926 5966 932 sw
rect 6708 926 8186 932
rect 8238 926 8264 978
rect 8316 932 10085 978
rect 10137 932 10517 984
rect 10569 932 10949 984
rect 11001 932 11381 984
rect 11433 932 11814 984
rect 11866 932 12245 984
rect 12297 932 12299 984
rect 8316 926 12299 932
rect 5575 898 5966 926
tri 5966 898 5994 926 sw
rect 5575 897 5994 898
rect 4883 892 5994 897
tri 5994 892 6000 898 sw
rect 7709 892 15105 898
rect 4883 878 6000 892
tri 6000 878 6014 892 sw
rect 4883 873 7146 878
rect 4883 821 4887 873
rect 4939 821 5099 873
rect 5151 821 5311 873
rect 5363 821 5523 873
rect 5575 856 7146 873
rect 5575 821 6793 856
rect 4883 800 6793 821
rect 6849 800 6888 856
rect 6944 800 6984 856
rect 7040 800 7080 856
rect 7136 800 7146 856
rect 4883 798 7146 800
rect 4883 746 4887 798
rect 4939 746 5099 798
rect 5151 746 5311 798
rect 5363 746 5523 798
rect 5575 776 7146 798
rect 5575 746 6793 776
rect 4883 723 6793 746
rect 4883 671 4887 723
rect 4939 671 5099 723
rect 5151 671 5311 723
rect 5363 671 5523 723
rect 5575 720 6793 723
rect 6849 720 6888 776
rect 6944 720 6984 776
rect 7040 720 7080 776
rect 7136 720 7146 776
rect 7761 840 8141 892
rect 8193 840 8573 892
rect 8625 840 9005 892
rect 9057 840 9437 892
rect 9489 840 9869 892
rect 9921 840 10301 892
rect 10353 840 10733 892
rect 10785 840 11165 892
rect 11217 840 11597 892
rect 11649 840 12029 892
rect 12081 840 12461 892
rect 12513 840 12893 892
rect 12945 840 13325 892
rect 13377 840 13757 892
rect 13809 840 14189 892
rect 14241 840 14621 892
rect 14673 840 15053 892
rect 7709 828 15105 840
rect 7761 776 8141 828
rect 8193 776 8573 828
rect 8625 776 9005 828
rect 9057 776 9437 828
rect 9489 776 9869 828
rect 9921 776 10301 828
rect 10353 776 10733 828
rect 10785 776 11165 828
rect 11217 776 11597 828
rect 11649 776 12029 828
rect 12081 776 12461 828
rect 12513 776 12893 828
rect 12945 776 13325 828
rect 13377 776 13757 828
rect 13809 776 14189 828
rect 14241 776 14621 828
rect 14673 776 15053 828
rect 7709 770 15105 776
rect 5575 696 7146 720
rect 5575 671 6793 696
rect 4883 665 6793 671
tri 5654 640 5679 665 ne
rect 5679 640 6793 665
rect 6849 640 6888 696
rect 6944 640 6984 696
rect 7040 640 7080 696
rect 7136 640 7146 696
tri 5679 625 5694 640 ne
rect 5694 625 7146 640
rect 7493 736 9407 742
rect 7545 684 7925 736
rect 7977 684 9355 736
rect 7493 672 9407 684
rect 7545 620 7925 672
rect 7977 620 9355 672
rect 7493 614 9407 620
tri 6886 575 6895 584 se
rect 6895 575 9623 584
tri 6877 566 6886 575 se
rect 6886 566 9571 575
rect 1886 526 1938 541
rect 3504 560 5684 566
rect 3556 508 3690 560
rect 3742 508 3754 560
rect 3806 508 3933 560
rect 3985 508 4145 560
rect 4197 557 4357 560
rect 4409 557 4569 560
rect 3504 501 4190 508
rect 4246 501 4270 557
rect 4326 501 4350 557
rect 4409 508 4430 557
rect 4406 501 4430 508
rect 4486 501 4510 557
rect 4566 508 4569 557
rect 4621 508 4781 560
rect 4833 508 4993 560
rect 5045 508 5205 560
rect 5257 508 5417 560
rect 5469 508 5629 560
rect 5681 508 5684 560
tri 6834 523 6877 566 se
rect 6877 523 9571 566
tri 6822 511 6834 523 se
rect 6834 511 6908 523
tri 6908 511 6920 523 nw
tri 9537 511 9549 523 ne
rect 9549 511 9623 523
rect 4566 501 5684 508
rect 3504 485 5684 501
tri 6809 498 6822 511 se
rect 6822 498 6895 511
tri 6895 498 6908 511 nw
tri 9549 498 9562 511 ne
rect 9562 498 9571 511
rect 1886 468 1938 474
rect 3246 472 3302 481
rect 3246 407 3302 416
rect 3246 392 3248 407
rect 3300 392 3302 407
rect 3246 327 3302 336
rect 3556 433 3690 485
rect 3742 433 3754 485
rect 3806 484 5684 485
rect 3806 433 3933 484
rect 3504 432 3933 433
rect 3985 432 4145 484
rect 4197 449 4357 484
rect 4409 449 4569 484
rect 3504 410 4190 432
rect 3556 358 3690 410
rect 3742 358 3754 410
rect 3806 409 4190 410
rect 3806 358 3933 409
rect 3504 357 3933 358
rect 3985 357 4145 409
rect 4246 393 4270 449
rect 4326 393 4350 449
rect 4409 432 4430 449
rect 4406 409 4430 432
rect 4409 393 4430 409
rect 4486 393 4510 449
rect 4566 432 4569 449
rect 4621 432 4781 484
rect 4833 432 4993 484
rect 5045 432 5205 484
rect 5257 432 5417 484
rect 5469 432 5629 484
rect 5681 432 5684 484
rect 4566 409 5684 432
rect 4566 393 4569 409
rect 4197 357 4357 393
rect 4409 357 4569 393
rect 4621 357 4781 409
rect 4833 357 4993 409
rect 5045 357 5205 409
rect 5257 357 5417 409
rect 5469 357 5629 409
rect 5681 357 5684 409
tri 6785 474 6809 498 se
rect 6809 474 6871 498
tri 6871 474 6895 498 nw
tri 9562 489 9571 498 ne
rect 6785 459 6856 474
tri 6856 459 6871 474 nw
rect 6785 453 6850 459
tri 6850 453 6856 459 nw
rect 9571 453 9623 459
rect 3504 341 5684 357
rect 3504 334 4190 341
rect 3556 282 3690 334
rect 3742 282 3754 334
rect 3806 282 3933 334
rect 3985 282 4145 334
rect 4246 285 4270 341
rect 4326 285 4350 341
rect 4406 334 4430 341
rect 4409 285 4430 334
rect 4486 285 4510 341
rect 4566 334 5684 341
rect 6542 364 6594 370
rect 4566 285 4569 334
rect 4197 282 4357 285
rect 4409 282 4569 285
rect 4621 282 4781 334
rect 4833 282 4993 334
rect 5045 282 5205 334
rect 5257 282 5417 334
rect 5469 282 5629 334
rect 5681 282 5684 334
rect 3504 276 5684 282
rect 5730 334 5782 340
rect 5730 270 5782 282
tri 5708 230 5730 252 se
rect 1580 178 1586 230
rect 1638 178 1656 230
rect 1708 178 1726 230
rect 1778 178 1796 230
rect 1848 178 1866 230
rect 1918 178 1936 230
rect 1988 178 2006 230
rect 2058 178 2076 230
rect 2128 178 2146 230
rect 2198 178 2216 230
rect 2268 178 2285 230
rect 2337 178 2959 230
rect 3011 178 3029 230
rect 3081 178 3098 230
rect 3150 178 3167 230
rect 3219 178 3236 230
rect 3288 178 3305 230
rect 3357 178 3374 230
rect 3426 218 5026 230
tri 5026 218 5038 230 sw
tri 5696 218 5708 230 se
rect 5708 218 5730 230
rect 6542 300 6594 312
tri 5782 248 5795 261 sw
tri 6529 248 6542 261 se
rect 6785 338 6845 453
tri 6845 448 6850 453 nw
tri 6845 338 6876 369 sw
rect 6785 335 6876 338
tri 6876 335 6879 338 sw
rect 6785 283 6791 335
rect 6843 283 6855 335
rect 6907 283 6913 335
rect 15529 332 15581 338
rect 15529 267 15581 280
tri 15526 261 15529 264 se
rect 5782 230 5795 248
tri 5795 230 5813 248 sw
tri 6511 230 6529 248 se
rect 6529 230 6594 248
tri 6594 230 6625 261 sw
tri 15495 230 15526 261 se
rect 15526 230 15529 261
rect 5782 224 5813 230
tri 5813 224 5819 230 sw
tri 6108 224 6114 230 se
rect 6114 224 15529 230
rect 5782 218 5819 224
rect 3426 212 5038 218
tri 5038 212 5044 218 sw
tri 5690 212 5696 218 se
rect 5696 212 5819 218
tri 5819 212 5831 224 sw
tri 6096 212 6108 224 se
rect 6108 212 7227 224
rect 3426 178 7227 212
rect 1580 172 7227 178
rect 7279 172 8789 224
rect 8841 172 9221 224
rect 9273 172 9653 224
rect 9705 172 12677 224
rect 12729 172 13109 224
rect 13161 172 13541 224
rect 13593 172 13973 224
rect 14025 172 14405 224
rect 14457 172 14837 224
rect 14889 172 15418 224
rect 15470 215 15529 224
rect 15961 332 16013 338
rect 15961 267 16013 280
tri 15581 230 15615 264 sw
tri 15927 230 15961 264 se
rect 15581 215 15961 230
rect 15470 202 16013 215
rect 15470 172 15529 202
rect 1580 160 15529 172
rect 1580 108 1586 160
rect 1638 108 1656 160
rect 1708 108 1726 160
rect 1778 108 1796 160
rect 1848 108 1866 160
rect 1918 108 1936 160
rect 1988 108 2006 160
rect 2058 108 2076 160
rect 2128 108 2146 160
rect 2198 108 2216 160
rect 2268 108 2285 160
rect 2337 108 2959 160
rect 3011 108 3029 160
rect 3081 108 3098 160
rect 3150 108 3167 160
rect 3219 108 3236 160
rect 3288 108 3305 160
rect 3357 108 3374 160
rect 3426 108 7227 160
rect 7279 108 8789 160
rect 8841 108 9221 160
rect 9273 108 9653 160
rect 9705 108 12677 160
rect 12729 108 13109 160
rect 13161 108 13541 160
rect 13593 108 13973 160
rect 14025 108 14405 160
rect 14457 108 14837 160
rect 14889 108 15418 160
rect 15470 150 15529 160
rect 15581 150 15961 202
rect 15470 108 16013 150
rect 1580 96 16013 108
rect 1580 90 7227 96
rect 1580 38 1586 90
rect 1638 38 1656 90
rect 1708 38 1726 90
rect 1778 38 1796 90
rect 1848 38 1866 90
rect 1918 38 1936 90
rect 1988 38 2006 90
rect 2058 38 2076 90
rect 2128 38 2146 90
rect 2198 38 2216 90
rect 2268 38 2285 90
rect 2337 38 2959 90
rect 3011 38 3029 90
rect 3081 38 3098 90
rect 3150 38 3167 90
rect 3219 38 3236 90
rect 3288 38 3305 90
rect 3357 38 3374 90
rect 3426 44 7227 90
rect 7279 44 8789 96
rect 8841 44 9221 96
rect 9273 44 9653 96
rect 9705 44 12677 96
rect 12729 44 13109 96
rect 13161 44 13541 96
rect 13593 44 13973 96
rect 14025 44 14405 96
rect 14457 44 14837 96
rect 14889 44 15418 96
rect 15470 44 16013 96
rect 3426 38 16013 44
rect 1580 34 16013 38
tri 3510 -79 3623 34 ne
rect 15303 -196 15312 -140
rect 15368 -196 15392 -140
rect 15448 -158 15462 -140
tri 15462 -158 15480 -140 sw
rect 15448 -196 16294 -158
rect 3035 -885 3041 -833
rect 3035 -889 3044 -885
rect 3100 -889 3124 -833
rect 3183 -885 3189 -833
rect 3180 -889 3189 -885
rect 15303 -889 15312 -833
rect 15387 -885 15392 -833
rect 15451 -885 15457 -833
rect 15368 -889 15392 -885
rect 15448 -889 15457 -885
<< via2 >>
rect 4187 2927 4243 2983
rect 4268 2927 4324 2983
rect 4349 2927 4405 2983
rect 4431 2927 4487 2983
rect 4513 2927 4569 2983
rect 6793 2951 6849 3007
rect 6888 2951 6944 3007
rect 6984 2951 7040 3007
rect 7080 2951 7136 3007
rect 3345 2782 3401 2838
rect 3425 2782 3481 2838
rect 3505 2782 3561 2838
rect 3345 2691 3401 2747
rect 3425 2691 3481 2747
rect 3505 2691 3561 2747
rect 3345 2599 3401 2655
rect 3425 2599 3481 2655
rect 3505 2599 3561 2655
rect 6795 1834 6851 1890
rect 6936 1834 6992 1890
rect 7077 1834 7133 1890
rect 3345 890 3401 946
rect 3425 890 3481 946
rect 3505 890 3561 946
rect 3345 782 3401 838
rect 3425 782 3481 838
rect 3505 782 3561 838
rect 3345 674 3401 730
rect 3425 674 3481 730
rect 3505 674 3561 730
rect 6793 800 6849 856
rect 6888 800 6944 856
rect 6984 800 7040 856
rect 7080 800 7136 856
rect 6793 720 6849 776
rect 6888 720 6944 776
rect 6984 720 7040 776
rect 7080 720 7136 776
rect 6793 640 6849 696
rect 6888 640 6944 696
rect 6984 640 7040 696
rect 7080 640 7136 696
rect 4190 508 4197 557
rect 4197 508 4246 557
rect 4190 501 4246 508
rect 4270 501 4326 557
rect 4350 508 4357 557
rect 4357 508 4406 557
rect 4350 501 4406 508
rect 4430 501 4486 557
rect 4510 501 4566 557
rect 3246 471 3302 472
rect 3246 419 3248 471
rect 3248 419 3300 471
rect 3300 419 3302 471
rect 3246 416 3302 419
rect 3246 355 3248 392
rect 3248 355 3300 392
rect 3300 355 3302 392
rect 3246 336 3302 355
rect 4190 432 4197 449
rect 4197 432 4246 449
rect 4190 409 4246 432
rect 4190 393 4197 409
rect 4197 393 4246 409
rect 4270 393 4326 449
rect 4350 432 4357 449
rect 4357 432 4406 449
rect 4350 409 4406 432
rect 4350 393 4357 409
rect 4357 393 4406 409
rect 4430 393 4486 449
rect 4510 393 4566 449
rect 4190 334 4246 341
rect 4190 285 4197 334
rect 4197 285 4246 334
rect 4270 285 4326 341
rect 4350 334 4406 341
rect 4350 285 4357 334
rect 4357 285 4406 334
rect 4430 285 4486 341
rect 4510 285 4566 341
rect 15312 -196 15368 -140
rect 15392 -196 15448 -140
rect 3044 -885 3093 -833
rect 3093 -885 3100 -833
rect 3044 -889 3100 -885
rect 3124 -885 3131 -833
rect 3131 -885 3180 -833
rect 3124 -889 3180 -885
rect 15312 -885 15335 -833
rect 15335 -885 15368 -833
rect 15392 -885 15399 -833
rect 15399 -885 15448 -833
rect 15312 -889 15368 -885
rect 15392 -889 15448 -885
<< metal3 >>
rect 3110 501 3184 3318
rect 4178 2983 4578 3024
rect 4178 2927 4187 2983
rect 4243 2927 4268 2983
rect 4324 2927 4349 2983
rect 4405 2927 4431 2983
rect 4487 2927 4513 2983
rect 4569 2927 4578 2983
rect 3329 2838 3570 2847
rect 3329 2782 3345 2838
rect 3401 2782 3425 2838
rect 3481 2782 3505 2838
rect 3561 2782 3570 2838
rect 3329 2747 3570 2782
rect 3329 2691 3345 2747
rect 3401 2691 3425 2747
rect 3481 2691 3505 2747
rect 3561 2691 3570 2747
rect 3329 2655 3570 2691
rect 3329 2599 3345 2655
rect 3401 2599 3425 2655
rect 3481 2599 3505 2655
rect 3561 2599 3570 2655
rect 3329 946 3570 2599
rect 3329 890 3345 946
rect 3401 890 3425 946
rect 3481 890 3505 946
rect 3561 890 3570 946
rect 3329 838 3570 890
rect 3329 782 3345 838
rect 3401 782 3425 838
rect 3481 782 3505 838
rect 3561 782 3570 838
rect 3329 730 3570 782
rect 3329 674 3345 730
rect 3401 674 3425 730
rect 3481 674 3505 730
rect 3561 674 3570 730
rect 3329 665 3570 674
rect 4178 557 4578 2927
rect 6786 3007 7142 3064
rect 6786 2951 6793 3007
rect 6849 2951 6888 3007
rect 6944 2951 6984 3007
rect 7040 2951 7080 3007
rect 7136 2951 7142 3007
rect 6786 1890 7142 2951
rect 6786 1834 6795 1890
rect 6851 1834 6936 1890
rect 6992 1834 7077 1890
rect 7133 1834 7142 1890
rect 6786 856 7142 1834
rect 6786 800 6793 856
rect 6849 800 6888 856
rect 6944 800 6984 856
rect 7040 800 7080 856
rect 7136 800 7142 856
rect 6786 776 7142 800
rect 6786 720 6793 776
rect 6849 720 6888 776
rect 6944 720 6984 776
rect 7040 720 7080 776
rect 7136 720 7142 776
rect 6786 696 7142 720
rect 6786 640 6793 696
rect 6849 640 6888 696
rect 6944 640 6984 696
rect 7040 640 7080 696
rect 7136 640 7142 696
rect 6786 629 7142 640
tri 3184 501 3226 543 sw
rect 4178 501 4190 557
rect 4246 501 4270 557
rect 4326 501 4350 557
rect 4406 501 4430 557
rect 4486 501 4510 557
rect 4566 501 4578 557
rect 3110 477 3226 501
tri 3226 477 3250 501 sw
rect 3110 472 3307 477
rect 3110 416 3246 472
rect 3302 416 3307 472
rect 3110 392 3307 416
rect 3110 336 3246 392
rect 3302 336 3307 392
rect 3110 331 3307 336
rect 4178 449 4578 501
rect 4178 393 4190 449
rect 4246 393 4270 449
rect 4326 393 4350 449
rect 4406 393 4430 449
rect 4486 393 4510 449
rect 4566 393 4578 449
rect 4178 341 4578 393
rect 3110 285 3197 331
tri 3197 285 3243 331 nw
rect 4178 285 4190 341
rect 4246 285 4270 341
rect 4326 285 4350 341
rect 4406 285 4430 341
rect 4486 285 4510 341
rect 4566 285 4578 341
tri 3039 -828 3110 -757 se
rect 3110 -828 3185 285
tri 3185 273 3197 285 nw
rect 4178 276 4578 285
rect 3039 -833 3185 -828
rect 3039 -889 3044 -833
rect 3100 -889 3124 -833
rect 3180 -889 3185 -833
rect 3039 -894 3185 -889
rect 15307 -140 15453 -135
rect 15307 -196 15312 -140
rect 15368 -196 15392 -140
rect 15448 -196 15453 -140
rect 15307 -833 15453 -196
rect 15307 -889 15312 -833
rect 15368 -889 15392 -833
rect 15448 -889 15453 -833
rect 15307 -894 15453 -889
use sky130_fd_pr__pfet_01v8__example_55959141808540  sky130_fd_pr__pfet_01v8__example_55959141808540_0
timestamp 1619862920
transform -1 0 6235 0 1 1921
box -28 0 404 471
use sky130_fd_pr__nfet_01v8__example_55959141808535  sky130_fd_pr__nfet_01v8__example_55959141808535_1
timestamp 1619862920
transform 1 0 15583 0 1 148
box -28 0 404 471
use sky130_fd_pr__nfet_01v8__example_55959141808535  sky130_fd_pr__nfet_01v8__example_55959141808535_0
timestamp 1619862920
transform -1 0 8571 0 1 148
box -28 0 404 471
use sky130_fd_pr__nfet_01v8__example_55959141808527  sky130_fd_pr__nfet_01v8__example_55959141808527_2
timestamp 1619862920
transform 1 0 5945 0 1 948
box -28 0 620 97
use sky130_fd_pr__nfet_01v8__example_55959141808527  sky130_fd_pr__nfet_01v8__example_55959141808527_1
timestamp 1619862920
transform 1 0 5945 0 1 618
box -28 0 620 97
use sky130_fd_pr__nfet_01v8__example_55959141808527  sky130_fd_pr__nfet_01v8__example_55959141808527_0
timestamp 1619862920
transform 1 0 5945 0 -1 446
box -28 0 620 97
use sky130_fd_pr__nfet_01v8__example_55959141808528  sky130_fd_pr__nfet_01v8__example_55959141808528_1
timestamp 1619862920
transform 1 0 7015 0 1 548
box -28 0 128 267
use sky130_fd_pr__nfet_01v8__example_55959141808528  sky130_fd_pr__nfet_01v8__example_55959141808528_0
timestamp 1619862920
transform 1 0 -56 0 1 2238
box -28 0 128 267
use sky130_fd_pr__pfet_01v8__example_55959141808537  sky130_fd_pr__pfet_01v8__example_55959141808537_0
timestamp 1619862920
transform 1 0 3371 0 1 1921
box -28 0 752 471
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_7
timestamp 1619862920
transform -1 0 10885 0 1 1921
box -28 0 284 471
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_6
timestamp 1619862920
transform -1 0 10261 0 1 1921
box -28 0 284 471
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_5
timestamp 1619862920
transform -1 0 9949 0 1 1921
box -28 0 284 471
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_4
timestamp 1619862920
transform -1 0 11197 0 1 1921
box -28 0 284 471
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_3
timestamp 1619862920
transform -1 0 11509 0 1 1921
box -28 0 284 471
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_2
timestamp 1619862920
transform -1 0 10573 0 1 1921
box -28 0 284 471
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_1
timestamp 1619862920
transform 1 0 765 0 1 1921
box -28 0 284 471
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_0
timestamp 1619862920
transform -1 0 5803 0 1 1921
box -28 0 284 471
use sky130_fd_pr__pfet_01v8__example_55959141808542  sky130_fd_pr__pfet_01v8__example_55959141808542_2
timestamp 1619862920
transform 1 0 8063 0 1 1921
box -28 0 596 471
use sky130_fd_pr__pfet_01v8__example_55959141808542  sky130_fd_pr__pfet_01v8__example_55959141808542_1
timestamp 1619862920
transform 1 0 2123 0 1 1921
box -28 0 596 471
use sky130_fd_pr__pfet_01v8__example_55959141808542  sky130_fd_pr__pfet_01v8__example_55959141808542_0
timestamp 1619862920
transform 1 0 2747 0 1 1921
box -28 0 596 471
use sky130_fd_pr__pfet_01v8__example_55959141808541  sky130_fd_pr__pfet_01v8__example_55959141808541_0
timestamp 1619862920
transform 1 0 7415 0 1 1921
box -28 0 620 471
use sky130_fd_pr__pfet_01v8__example_55959141808539  sky130_fd_pr__pfet_01v8__example_55959141808539_0
timestamp 1619862920
transform 1 0 1187 0 1 1921
box -28 0 908 471
use sky130_fd_pr__pfet_01v8__example_55959141808538  sky130_fd_pr__pfet_01v8__example_55959141808538_1
timestamp 1619862920
transform 1 0 4835 0 1 148
box -28 0 820 471
use sky130_fd_pr__pfet_01v8__example_55959141808538  sky130_fd_pr__pfet_01v8__example_55959141808538_0
timestamp 1619862920
transform 1 0 3987 0 1 148
box -28 0 820 471
use sky130_fd_pr__nfet_01v8__example_55959141808534  sky130_fd_pr__nfet_01v8__example_55959141808534_0
timestamp 1619862920
transform -1 0 8139 0 1 148
box -28 0 620 471
use sky130_fd_pr__nfet_01v8__example_55959141808531  sky130_fd_pr__nfet_01v8__example_55959141808531_2
timestamp 1619862920
transform 1 0 8627 0 1 148
box -28 0 1268 471
use sky130_fd_pr__nfet_01v8__example_55959141808531  sky130_fd_pr__nfet_01v8__example_55959141808531_1
timestamp 1619862920
transform 1 0 9923 0 1 148
box -28 0 1268 471
use sky130_fd_pr__nfet_01v8__example_55959141808531  sky130_fd_pr__nfet_01v8__example_55959141808531_0
timestamp 1619862920
transform 1 0 11219 0 1 148
box -28 0 1268 471
use sky130_fd_pr__nfet_01v8__example_55959141808530  sky130_fd_pr__nfet_01v8__example_55959141808530_0
timestamp 1619862920
transform 1 0 12515 0 1 148
box -28 0 2564 471
use sky130_fd_pr__nfet_01v8__example_55959141808529  sky130_fd_pr__nfet_01v8__example_55959141808529_0
timestamp 1619862920
transform -1 0 15417 0 1 548
box -28 0 228 267
use sky130_fd_pr__nfet_01v8__example_55959141808230  sky130_fd_pr__nfet_01v8__example_55959141808230_0
timestamp 1619862920
transform 1 0 6703 0 1 548
box -28 0 284 267
use sky130_fd_pr__nfet_01v8__example_55959141808533  sky130_fd_pr__nfet_01v8__example_55959141808533_0
timestamp 1619862920
transform 1 0 7281 0 1 148
box -28 0 128 471
use sky130_fd_pr__pfet_01v8__example_5595914180837  sky130_fd_pr__pfet_01v8__example_5595914180837_0
timestamp 1619862920
transform 1 0 4261 0 1 1921
box -28 0 284 267
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1619862920
transform 1 0 2004 0 1 14
box -46 24 399 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1619862920
transform -1 0 3456 0 1 17
box -42 24 569 1116
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1619862920
transform 1 0 1539 0 1 14
box 0 24 534 1116
use sky130_fd_pr__pfet_01v8__example_55959141808536  sky130_fd_pr__pfet_01v8__example_55959141808536_0
timestamp 1619862920
transform 1 0 6401 0 1 2321
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808532  sky130_fd_pr__nfet_01v8__example_55959141808532_0
timestamp 1619862920
transform 0 -1 16862 1 0 1963
box -28 0 680 981
use sky130_fd_pr__nfet_01v8__example_55959141808532  sky130_fd_pr__nfet_01v8__example_55959141808532_1
timestamp 1619862920
transform 0 -1 14218 1 0 1963
box -28 0 680 981
<< labels >>
flabel metal2 s 152 3162 402 3292 3 FreeSans 200 0 0 0 VDDIO_Q
port 1 nsew
flabel metal2 s 4338 2922 4472 3010 3 FreeSans 200 0 0 0 VCCHIB
port 2 nsew
flabel metal2 s 136 1493 256 1533 3 FreeSans 200 0 0 0 IN_H
port 3 nsew
flabel metal2 s 132 1413 224 1455 3 FreeSans 200 0 0 0 IN_VT
port 4 nsew
flabel metal2 s 131 1741 213 1779 3 FreeSans 200 0 0 0 MODE_REF_N
port 5 nsew
flabel metal2 s 17149 2235 17217 2342 3 FreeSans 200 0 0 0 VREFIN
port 6 nsew
flabel metal2 s 93 2032 163 2076 3 FreeSans 200 0 0 0 MODE_VCCD_N
port 7 nsew
flabel metal2 s 89 1953 180 1995 3 FreeSans 200 0 0 0 MODE_NORMAL_N
port 8 nsew
flabel metal2 s 94 1840 193 1878 3 FreeSans 200 0 0 0 MODE_REF_3V_N
port 9 nsew
flabel metal2 s 3973 1654 4053 1697 3 FreeSans 200 0 0 0 OUT
port 10 nsew
flabel metal2 s 128 1581 215 1617 3 FreeSans 200 0 0 0 OUT_N
port 11 nsew
flabel metal2 s 1617 53 1912 215 3 FreeSans 200 0 0 0 VSSD
port 12 nsew
flabel metal1 s 1689 350 1715 444 3 FreeSans 200 0 0 0 VTRIP_SEL_H
port 13 nsew
flabel metal1 s 7030 1199 7127 1232 3 FreeSans 200 0 0 0 EN_H_N
port 14 nsew
flabel metal1 s 15261 1201 15381 1230 3 FreeSans 200 0 0 0 VTRIP_SEL_H_N
port 15 nsew
flabel metal1 s 1812 908 1946 1038 3 FreeSans 200 0 0 0 VDDIO_Q
port 1 nsew
flabel metal1 s 5106 3168 5106 3168 3 FreeSans 200 0 0 0 VSSD
port 12 nsew
flabel comment s 13210 2838 13210 2838 0 FreeSans 200 0 0 0 CONDIODE
flabel comment s 16110 2838 16110 2838 0 FreeSans 200 0 0 0 CONDIODE
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 36158954
string GDS_START 35731676
<< end >>
