magic
tech sky130A
magscale 1 2
timestamp 1619862920
<< checkpaint >>
rect -25770 -4648 3730 18180
<< dnwell >>
rect -23658 7540 -22197 14448
<< nwell >>
rect -22303 14544 -21999 16920
rect -23743 14242 -21999 14544
rect -23743 7746 -23441 14242
rect -22303 7746 -21999 14242
rect -23743 7444 -21999 7746
rect -22303 7082 -21999 7444
rect -23283 2932 -22789 3664
rect -1000 0 1132 1118
<< pwell >>
rect -23381 14028 -22603 14182
rect -23381 9446 -23227 14028
rect -22757 9446 -22603 14028
rect -23381 8794 -22603 9446
rect -23381 7981 -23227 8794
rect -22757 7981 -22603 8794
rect -23381 7827 -22603 7981
<< mvnmos >>
rect -23120 8820 -23020 9420
rect -22964 8820 -22864 9420
<< mvpmos >>
rect -23164 2998 -23064 3598
rect -23008 2998 -22908 3598
rect -934 899 1066 999
rect -934 743 1066 843
rect -934 587 1066 687
rect -934 431 1066 531
rect -934 275 1066 375
rect -934 119 1066 219
<< mvndiff >>
rect -23173 9342 -23120 9420
rect -23173 9308 -23165 9342
rect -23131 9308 -23120 9342
rect -23173 9274 -23120 9308
rect -23173 9240 -23165 9274
rect -23131 9240 -23120 9274
rect -23173 9206 -23120 9240
rect -23173 9172 -23165 9206
rect -23131 9172 -23120 9206
rect -23173 9138 -23120 9172
rect -23173 9104 -23165 9138
rect -23131 9104 -23120 9138
rect -23173 9070 -23120 9104
rect -23173 9036 -23165 9070
rect -23131 9036 -23120 9070
rect -23173 9002 -23120 9036
rect -23173 8968 -23165 9002
rect -23131 8968 -23120 9002
rect -23173 8934 -23120 8968
rect -23173 8900 -23165 8934
rect -23131 8900 -23120 8934
rect -23173 8866 -23120 8900
rect -23173 8832 -23165 8866
rect -23131 8832 -23120 8866
rect -23173 8820 -23120 8832
rect -23020 9342 -22964 9420
rect -23020 9308 -23009 9342
rect -22975 9308 -22964 9342
rect -23020 9274 -22964 9308
rect -23020 9240 -23009 9274
rect -22975 9240 -22964 9274
rect -23020 9206 -22964 9240
rect -23020 9172 -23009 9206
rect -22975 9172 -22964 9206
rect -23020 9138 -22964 9172
rect -23020 9104 -23009 9138
rect -22975 9104 -22964 9138
rect -23020 9070 -22964 9104
rect -23020 9036 -23009 9070
rect -22975 9036 -22964 9070
rect -23020 9002 -22964 9036
rect -23020 8968 -23009 9002
rect -22975 8968 -22964 9002
rect -23020 8934 -22964 8968
rect -23020 8900 -23009 8934
rect -22975 8900 -22964 8934
rect -23020 8866 -22964 8900
rect -23020 8832 -23009 8866
rect -22975 8832 -22964 8866
rect -23020 8820 -22964 8832
rect -22864 9342 -22811 9420
rect -22864 9308 -22853 9342
rect -22819 9308 -22811 9342
rect -22864 9274 -22811 9308
rect -22864 9240 -22853 9274
rect -22819 9240 -22811 9274
rect -22864 9206 -22811 9240
rect -22864 9172 -22853 9206
rect -22819 9172 -22811 9206
rect -22864 9138 -22811 9172
rect -22864 9104 -22853 9138
rect -22819 9104 -22811 9138
rect -22864 9070 -22811 9104
rect -22864 9036 -22853 9070
rect -22819 9036 -22811 9070
rect -22864 9002 -22811 9036
rect -22864 8968 -22853 9002
rect -22819 8968 -22811 9002
rect -22864 8934 -22811 8968
rect -22864 8900 -22853 8934
rect -22819 8900 -22811 8934
rect -22864 8866 -22811 8900
rect -22864 8832 -22853 8866
rect -22819 8832 -22811 8866
rect -22864 8820 -22811 8832
<< mvpdiff >>
rect -23217 3586 -23164 3598
rect -23217 3552 -23209 3586
rect -23175 3552 -23164 3586
rect -23217 3518 -23164 3552
rect -23217 3484 -23209 3518
rect -23175 3484 -23164 3518
rect -23217 3450 -23164 3484
rect -23217 3416 -23209 3450
rect -23175 3416 -23164 3450
rect -23217 3382 -23164 3416
rect -23217 3348 -23209 3382
rect -23175 3348 -23164 3382
rect -23217 3314 -23164 3348
rect -23217 3280 -23209 3314
rect -23175 3280 -23164 3314
rect -23217 3246 -23164 3280
rect -23217 3212 -23209 3246
rect -23175 3212 -23164 3246
rect -23217 3178 -23164 3212
rect -23217 3144 -23209 3178
rect -23175 3144 -23164 3178
rect -23217 3110 -23164 3144
rect -23217 3076 -23209 3110
rect -23175 3076 -23164 3110
rect -23217 2998 -23164 3076
rect -23064 3586 -23008 3598
rect -23064 3552 -23053 3586
rect -23019 3552 -23008 3586
rect -23064 3518 -23008 3552
rect -23064 3484 -23053 3518
rect -23019 3484 -23008 3518
rect -23064 3450 -23008 3484
rect -23064 3416 -23053 3450
rect -23019 3416 -23008 3450
rect -23064 3382 -23008 3416
rect -23064 3348 -23053 3382
rect -23019 3348 -23008 3382
rect -23064 3314 -23008 3348
rect -23064 3280 -23053 3314
rect -23019 3280 -23008 3314
rect -23064 3246 -23008 3280
rect -23064 3212 -23053 3246
rect -23019 3212 -23008 3246
rect -23064 3178 -23008 3212
rect -23064 3144 -23053 3178
rect -23019 3144 -23008 3178
rect -23064 3110 -23008 3144
rect -23064 3076 -23053 3110
rect -23019 3076 -23008 3110
rect -23064 2998 -23008 3076
rect -22908 3586 -22855 3598
rect -22908 3552 -22897 3586
rect -22863 3552 -22855 3586
rect -22908 3518 -22855 3552
rect -22908 3484 -22897 3518
rect -22863 3484 -22855 3518
rect -22908 3450 -22855 3484
rect -22908 3416 -22897 3450
rect -22863 3416 -22855 3450
rect -22908 3382 -22855 3416
rect -22908 3348 -22897 3382
rect -22863 3348 -22855 3382
rect -22908 3314 -22855 3348
rect -22908 3280 -22897 3314
rect -22863 3280 -22855 3314
rect -22908 3246 -22855 3280
rect -22908 3212 -22897 3246
rect -22863 3212 -22855 3246
rect -22908 3178 -22855 3212
rect -22908 3144 -22897 3178
rect -22863 3144 -22855 3178
rect -22908 3110 -22855 3144
rect -22908 3076 -22897 3110
rect -22863 3076 -22855 3110
rect -22908 2998 -22855 3076
rect -934 1044 1066 1052
rect -934 1010 -884 1044
rect -850 1010 -816 1044
rect -782 1010 -748 1044
rect -714 1010 -680 1044
rect -646 1010 -612 1044
rect -578 1010 -544 1044
rect -510 1010 -476 1044
rect -442 1010 -408 1044
rect -374 1010 -340 1044
rect -306 1010 -272 1044
rect -238 1010 -204 1044
rect -170 1010 -136 1044
rect -102 1010 -68 1044
rect -34 1010 0 1044
rect 34 1010 68 1044
rect 102 1010 136 1044
rect 170 1010 204 1044
rect 238 1010 272 1044
rect 306 1010 340 1044
rect 374 1010 408 1044
rect 442 1010 476 1044
rect 510 1010 544 1044
rect 578 1010 612 1044
rect 646 1010 680 1044
rect 714 1010 748 1044
rect 782 1010 816 1044
rect 850 1010 884 1044
rect 918 1010 952 1044
rect 986 1010 1020 1044
rect 1054 1010 1066 1044
rect -934 999 1066 1010
rect -934 888 1066 899
rect -934 854 -884 888
rect -850 854 -816 888
rect -782 854 -748 888
rect -714 854 -680 888
rect -646 854 -612 888
rect -578 854 -544 888
rect -510 854 -476 888
rect -442 854 -408 888
rect -374 854 -340 888
rect -306 854 -272 888
rect -238 854 -204 888
rect -170 854 -136 888
rect -102 854 -68 888
rect -34 854 0 888
rect 34 854 68 888
rect 102 854 136 888
rect 170 854 204 888
rect 238 854 272 888
rect 306 854 340 888
rect 374 854 408 888
rect 442 854 476 888
rect 510 854 544 888
rect 578 854 612 888
rect 646 854 680 888
rect 714 854 748 888
rect 782 854 816 888
rect 850 854 884 888
rect 918 854 952 888
rect 986 854 1020 888
rect 1054 854 1066 888
rect -934 843 1066 854
rect -934 732 1066 743
rect -934 698 -884 732
rect -850 698 -816 732
rect -782 698 -748 732
rect -714 698 -680 732
rect -646 698 -612 732
rect -578 698 -544 732
rect -510 698 -476 732
rect -442 698 -408 732
rect -374 698 -340 732
rect -306 698 -272 732
rect -238 698 -204 732
rect -170 698 -136 732
rect -102 698 -68 732
rect -34 698 0 732
rect 34 698 68 732
rect 102 698 136 732
rect 170 698 204 732
rect 238 698 272 732
rect 306 698 340 732
rect 374 698 408 732
rect 442 698 476 732
rect 510 698 544 732
rect 578 698 612 732
rect 646 698 680 732
rect 714 698 748 732
rect 782 698 816 732
rect 850 698 884 732
rect 918 698 952 732
rect 986 698 1020 732
rect 1054 698 1066 732
rect -934 687 1066 698
rect -934 576 1066 587
rect -934 542 -884 576
rect -850 542 -816 576
rect -782 542 -748 576
rect -714 542 -680 576
rect -646 542 -612 576
rect -578 542 -544 576
rect -510 542 -476 576
rect -442 542 -408 576
rect -374 542 -340 576
rect -306 542 -272 576
rect -238 542 -204 576
rect -170 542 -136 576
rect -102 542 -68 576
rect -34 542 0 576
rect 34 542 68 576
rect 102 542 136 576
rect 170 542 204 576
rect 238 542 272 576
rect 306 542 340 576
rect 374 542 408 576
rect 442 542 476 576
rect 510 542 544 576
rect 578 542 612 576
rect 646 542 680 576
rect 714 542 748 576
rect 782 542 816 576
rect 850 542 884 576
rect 918 542 952 576
rect 986 542 1020 576
rect 1054 542 1066 576
rect -934 531 1066 542
rect -934 420 1066 431
rect -934 386 -884 420
rect -850 386 -816 420
rect -782 386 -748 420
rect -714 386 -680 420
rect -646 386 -612 420
rect -578 386 -544 420
rect -510 386 -476 420
rect -442 386 -408 420
rect -374 386 -340 420
rect -306 386 -272 420
rect -238 386 -204 420
rect -170 386 -136 420
rect -102 386 -68 420
rect -34 386 0 420
rect 34 386 68 420
rect 102 386 136 420
rect 170 386 204 420
rect 238 386 272 420
rect 306 386 340 420
rect 374 386 408 420
rect 442 386 476 420
rect 510 386 544 420
rect 578 386 612 420
rect 646 386 680 420
rect 714 386 748 420
rect 782 386 816 420
rect 850 386 884 420
rect 918 386 952 420
rect 986 386 1020 420
rect 1054 386 1066 420
rect -934 375 1066 386
rect -934 264 1066 275
rect -934 230 -884 264
rect -850 230 -816 264
rect -782 230 -748 264
rect -714 230 -680 264
rect -646 230 -612 264
rect -578 230 -544 264
rect -510 230 -476 264
rect -442 230 -408 264
rect -374 230 -340 264
rect -306 230 -272 264
rect -238 230 -204 264
rect -170 230 -136 264
rect -102 230 -68 264
rect -34 230 0 264
rect 34 230 68 264
rect 102 230 136 264
rect 170 230 204 264
rect 238 230 272 264
rect 306 230 340 264
rect 374 230 408 264
rect 442 230 476 264
rect 510 230 544 264
rect 578 230 612 264
rect 646 230 680 264
rect 714 230 748 264
rect 782 230 816 264
rect 850 230 884 264
rect 918 230 952 264
rect 986 230 1020 264
rect 1054 230 1066 264
rect -934 219 1066 230
rect -934 108 1066 119
rect -934 74 -884 108
rect -850 74 -816 108
rect -782 74 -748 108
rect -714 74 -680 108
rect -646 74 -612 108
rect -578 74 -544 108
rect -510 74 -476 108
rect -442 74 -408 108
rect -374 74 -340 108
rect -306 74 -272 108
rect -238 74 -204 108
rect -170 74 -136 108
rect -102 74 -68 108
rect -34 74 0 108
rect 34 74 68 108
rect 102 74 136 108
rect 170 74 204 108
rect 238 74 272 108
rect 306 74 340 108
rect 374 74 408 108
rect 442 74 476 108
rect 510 74 544 108
rect 578 74 612 108
rect 646 74 680 108
rect 714 74 748 108
rect 782 74 816 108
rect 850 74 884 108
rect 918 74 952 108
rect 986 74 1020 108
rect 1054 74 1066 108
rect -934 66 1066 74
<< mvndiffc >>
rect -23165 9308 -23131 9342
rect -23165 9240 -23131 9274
rect -23165 9172 -23131 9206
rect -23165 9104 -23131 9138
rect -23165 9036 -23131 9070
rect -23165 8968 -23131 9002
rect -23165 8900 -23131 8934
rect -23165 8832 -23131 8866
rect -23009 9308 -22975 9342
rect -23009 9240 -22975 9274
rect -23009 9172 -22975 9206
rect -23009 9104 -22975 9138
rect -23009 9036 -22975 9070
rect -23009 8968 -22975 9002
rect -23009 8900 -22975 8934
rect -23009 8832 -22975 8866
rect -22853 9308 -22819 9342
rect -22853 9240 -22819 9274
rect -22853 9172 -22819 9206
rect -22853 9104 -22819 9138
rect -22853 9036 -22819 9070
rect -22853 8968 -22819 9002
rect -22853 8900 -22819 8934
rect -22853 8832 -22819 8866
<< mvpdiffc >>
rect -23209 3552 -23175 3586
rect -23209 3484 -23175 3518
rect -23209 3416 -23175 3450
rect -23209 3348 -23175 3382
rect -23209 3280 -23175 3314
rect -23209 3212 -23175 3246
rect -23209 3144 -23175 3178
rect -23209 3076 -23175 3110
rect -23053 3552 -23019 3586
rect -23053 3484 -23019 3518
rect -23053 3416 -23019 3450
rect -23053 3348 -23019 3382
rect -23053 3280 -23019 3314
rect -23053 3212 -23019 3246
rect -23053 3144 -23019 3178
rect -23053 3076 -23019 3110
rect -22897 3552 -22863 3586
rect -22897 3484 -22863 3518
rect -22897 3416 -22863 3450
rect -22897 3348 -22863 3382
rect -22897 3280 -22863 3314
rect -22897 3212 -22863 3246
rect -22897 3144 -22863 3178
rect -22897 3076 -22863 3110
rect -884 1010 -850 1044
rect -816 1010 -782 1044
rect -748 1010 -714 1044
rect -680 1010 -646 1044
rect -612 1010 -578 1044
rect -544 1010 -510 1044
rect -476 1010 -442 1044
rect -408 1010 -374 1044
rect -340 1010 -306 1044
rect -272 1010 -238 1044
rect -204 1010 -170 1044
rect -136 1010 -102 1044
rect -68 1010 -34 1044
rect 0 1010 34 1044
rect 68 1010 102 1044
rect 136 1010 170 1044
rect 204 1010 238 1044
rect 272 1010 306 1044
rect 340 1010 374 1044
rect 408 1010 442 1044
rect 476 1010 510 1044
rect 544 1010 578 1044
rect 612 1010 646 1044
rect 680 1010 714 1044
rect 748 1010 782 1044
rect 816 1010 850 1044
rect 884 1010 918 1044
rect 952 1010 986 1044
rect 1020 1010 1054 1044
rect -884 854 -850 888
rect -816 854 -782 888
rect -748 854 -714 888
rect -680 854 -646 888
rect -612 854 -578 888
rect -544 854 -510 888
rect -476 854 -442 888
rect -408 854 -374 888
rect -340 854 -306 888
rect -272 854 -238 888
rect -204 854 -170 888
rect -136 854 -102 888
rect -68 854 -34 888
rect 0 854 34 888
rect 68 854 102 888
rect 136 854 170 888
rect 204 854 238 888
rect 272 854 306 888
rect 340 854 374 888
rect 408 854 442 888
rect 476 854 510 888
rect 544 854 578 888
rect 612 854 646 888
rect 680 854 714 888
rect 748 854 782 888
rect 816 854 850 888
rect 884 854 918 888
rect 952 854 986 888
rect 1020 854 1054 888
rect -884 698 -850 732
rect -816 698 -782 732
rect -748 698 -714 732
rect -680 698 -646 732
rect -612 698 -578 732
rect -544 698 -510 732
rect -476 698 -442 732
rect -408 698 -374 732
rect -340 698 -306 732
rect -272 698 -238 732
rect -204 698 -170 732
rect -136 698 -102 732
rect -68 698 -34 732
rect 0 698 34 732
rect 68 698 102 732
rect 136 698 170 732
rect 204 698 238 732
rect 272 698 306 732
rect 340 698 374 732
rect 408 698 442 732
rect 476 698 510 732
rect 544 698 578 732
rect 612 698 646 732
rect 680 698 714 732
rect 748 698 782 732
rect 816 698 850 732
rect 884 698 918 732
rect 952 698 986 732
rect 1020 698 1054 732
rect -884 542 -850 576
rect -816 542 -782 576
rect -748 542 -714 576
rect -680 542 -646 576
rect -612 542 -578 576
rect -544 542 -510 576
rect -476 542 -442 576
rect -408 542 -374 576
rect -340 542 -306 576
rect -272 542 -238 576
rect -204 542 -170 576
rect -136 542 -102 576
rect -68 542 -34 576
rect 0 542 34 576
rect 68 542 102 576
rect 136 542 170 576
rect 204 542 238 576
rect 272 542 306 576
rect 340 542 374 576
rect 408 542 442 576
rect 476 542 510 576
rect 544 542 578 576
rect 612 542 646 576
rect 680 542 714 576
rect 748 542 782 576
rect 816 542 850 576
rect 884 542 918 576
rect 952 542 986 576
rect 1020 542 1054 576
rect -884 386 -850 420
rect -816 386 -782 420
rect -748 386 -714 420
rect -680 386 -646 420
rect -612 386 -578 420
rect -544 386 -510 420
rect -476 386 -442 420
rect -408 386 -374 420
rect -340 386 -306 420
rect -272 386 -238 420
rect -204 386 -170 420
rect -136 386 -102 420
rect -68 386 -34 420
rect 0 386 34 420
rect 68 386 102 420
rect 136 386 170 420
rect 204 386 238 420
rect 272 386 306 420
rect 340 386 374 420
rect 408 386 442 420
rect 476 386 510 420
rect 544 386 578 420
rect 612 386 646 420
rect 680 386 714 420
rect 748 386 782 420
rect 816 386 850 420
rect 884 386 918 420
rect 952 386 986 420
rect 1020 386 1054 420
rect -884 230 -850 264
rect -816 230 -782 264
rect -748 230 -714 264
rect -680 230 -646 264
rect -612 230 -578 264
rect -544 230 -510 264
rect -476 230 -442 264
rect -408 230 -374 264
rect -340 230 -306 264
rect -272 230 -238 264
rect -204 230 -170 264
rect -136 230 -102 264
rect -68 230 -34 264
rect 0 230 34 264
rect 68 230 102 264
rect 136 230 170 264
rect 204 230 238 264
rect 272 230 306 264
rect 340 230 374 264
rect 408 230 442 264
rect 476 230 510 264
rect 544 230 578 264
rect 612 230 646 264
rect 680 230 714 264
rect 748 230 782 264
rect 816 230 850 264
rect 884 230 918 264
rect 952 230 986 264
rect 1020 230 1054 264
rect -884 74 -850 108
rect -816 74 -782 108
rect -748 74 -714 108
rect -680 74 -646 108
rect -612 74 -578 108
rect -544 74 -510 108
rect -476 74 -442 108
rect -408 74 -374 108
rect -340 74 -306 108
rect -272 74 -238 108
rect -204 74 -170 108
rect -136 74 -102 108
rect -68 74 -34 108
rect 0 74 34 108
rect 68 74 102 108
rect 136 74 170 108
rect 204 74 238 108
rect 272 74 306 108
rect 340 74 374 108
rect 408 74 442 108
rect 476 74 510 108
rect 544 74 578 108
rect 612 74 646 108
rect 680 74 714 108
rect 748 74 782 108
rect 816 74 850 108
rect 884 74 918 108
rect 952 74 986 108
rect 1020 74 1054 108
<< psubdiff >>
rect -23355 14122 -23279 14156
rect -23245 14122 -23139 14156
rect -23355 14088 -23139 14122
rect -23253 14054 -23139 14088
rect -22697 14075 -22629 14156
rect -22697 14054 -22663 14075
rect -22731 14041 -22663 14054
rect -22731 14007 -22629 14041
rect -23355 7968 -23253 8002
rect -23321 7955 -23253 7968
rect -23321 7934 -23287 7955
rect -23355 7853 -23287 7934
rect -22777 7921 -22731 7955
rect -22777 7887 -22629 7921
rect -22777 7853 -22743 7887
rect -22709 7853 -22629 7887
<< mvnsubdiff >>
rect -22236 16886 -22066 16920
rect -23677 14410 -23609 14478
rect -23643 14376 -23609 14410
rect -23167 14444 -23132 14478
rect -23098 14444 -23063 14478
rect -23029 14444 -22994 14478
rect -22960 14444 -22925 14478
rect -22891 14444 -22856 14478
rect -22822 14444 -22787 14478
rect -22753 14444 -22718 14478
rect -22684 14444 -22649 14478
rect -22615 14444 -22580 14478
rect -22546 14444 -22511 14478
rect -22477 14444 -22442 14478
rect -22408 14444 -22373 14478
rect -22339 14444 -22304 14478
rect -23167 14410 -22304 14444
rect -23167 14376 -23132 14410
rect -23098 14376 -23063 14410
rect -23029 14376 -22994 14410
rect -22960 14376 -22925 14410
rect -22891 14376 -22856 14410
rect -22822 14376 -22787 14410
rect -22753 14376 -22718 14410
rect -22684 14376 -22649 14410
rect -22615 14376 -22580 14410
rect -22546 14376 -22511 14410
rect -22477 14376 -22442 14410
rect -22408 14376 -22373 14410
rect -22339 14376 -22304 14410
rect -23677 14341 -23541 14376
rect -23643 14307 -23609 14341
rect -23575 14308 -23541 14341
rect -23167 14342 -22304 14376
rect -23167 14308 -23132 14342
rect -23098 14308 -23063 14342
rect -23029 14308 -22994 14342
rect -22960 14308 -22925 14342
rect -22891 14308 -22856 14342
rect -22822 14308 -22787 14342
rect -22753 14308 -22718 14342
rect -22684 14308 -22649 14342
rect -22615 14308 -22580 14342
rect -22546 14308 -22511 14342
rect -22477 14308 -22442 14342
rect -22408 14308 -22373 14342
rect -22339 14308 -22304 14342
rect -23575 14307 -23507 14308
rect -23677 14273 -23507 14307
rect -23677 14272 -23541 14273
rect -23643 14238 -23609 14272
rect -23575 14239 -23541 14272
rect -23575 14238 -23507 14239
rect -23677 14204 -23507 14238
rect -23677 14203 -23541 14204
rect -23643 14169 -23609 14203
rect -23575 14170 -23541 14203
rect -23575 14169 -23507 14170
rect -23677 14135 -23507 14169
rect -23677 14134 -23541 14135
rect -23643 14100 -23609 14134
rect -23575 14101 -23541 14134
rect -23575 14100 -23507 14101
rect -23677 14066 -23507 14100
rect -23677 14065 -23541 14066
rect -23643 14031 -23609 14065
rect -23575 14032 -23541 14065
rect -23575 14031 -23507 14032
rect -23677 13997 -23507 14031
rect -23677 13996 -23541 13997
rect -23643 13962 -23609 13996
rect -23575 13963 -23541 13996
rect -23575 13962 -23507 13963
rect -23677 13928 -23507 13962
rect -23677 13927 -23541 13928
rect -23643 13893 -23609 13927
rect -23575 13894 -23541 13927
rect -23575 13893 -23507 13894
rect -23677 13859 -23507 13893
rect -23677 13858 -23541 13859
rect -23643 13824 -23609 13858
rect -23575 13825 -23541 13858
rect -23575 13824 -23507 13825
rect -23677 13790 -23507 13824
rect -23677 13789 -23541 13790
rect -23643 13755 -23609 13789
rect -23575 13756 -23541 13789
rect -23575 13755 -23507 13756
rect -23677 13721 -23507 13755
rect -23677 13720 -23541 13721
rect -23643 13686 -23609 13720
rect -23575 13687 -23541 13720
rect -23575 13686 -23507 13687
rect -23677 13652 -23507 13686
rect -23677 13651 -23541 13652
rect -23643 13617 -23609 13651
rect -23575 13618 -23541 13651
rect -23575 13617 -23507 13618
rect -23677 13583 -23507 13617
rect -23677 13582 -23541 13583
rect -23643 13548 -23609 13582
rect -23575 13549 -23541 13582
rect -23575 13548 -23507 13549
rect -23677 13514 -23507 13548
rect -23677 13513 -23541 13514
rect -23643 13479 -23609 13513
rect -23575 13480 -23541 13513
rect -23575 13479 -23507 13480
rect -23677 13445 -23507 13479
rect -23677 13444 -23541 13445
rect -23643 13410 -23609 13444
rect -23575 13411 -23541 13444
rect -23575 13410 -23507 13411
rect -23677 13376 -23507 13410
rect -23677 13375 -23541 13376
rect -23643 13341 -23609 13375
rect -23575 13342 -23541 13375
rect -23575 13341 -23507 13342
rect -23677 13307 -23507 13341
rect -23677 13306 -23541 13307
rect -23643 13272 -23609 13306
rect -23575 13273 -23541 13306
rect -23575 13272 -23507 13273
rect -23677 13238 -23507 13272
rect -23677 13237 -23541 13238
rect -23643 13203 -23609 13237
rect -23575 13204 -23541 13237
rect -23575 13203 -23507 13204
rect -23677 13169 -23507 13203
rect -23677 13168 -23541 13169
rect -23643 13134 -23609 13168
rect -23575 13135 -23541 13168
rect -23575 13134 -23507 13135
rect -23677 13100 -23507 13134
rect -23677 13099 -23541 13100
rect -23643 13065 -23609 13099
rect -23575 13066 -23541 13099
rect -23575 13065 -23507 13066
rect -23677 13031 -23507 13065
rect -23677 13030 -23541 13031
rect -23643 12996 -23609 13030
rect -23575 12997 -23541 13030
rect -23575 12996 -23507 12997
rect -23677 12962 -23507 12996
rect -23677 12961 -23541 12962
rect -23643 12927 -23609 12961
rect -23575 12928 -23541 12961
rect -23575 12927 -23507 12928
rect -23677 12893 -23507 12927
rect -23677 12892 -23541 12893
rect -23643 12858 -23609 12892
rect -23575 12859 -23541 12892
rect -23575 12858 -23507 12859
rect -23677 12824 -23507 12858
rect -23677 12823 -23541 12824
rect -23643 12789 -23609 12823
rect -23575 12790 -23541 12823
rect -23575 12789 -23507 12790
rect -23677 12755 -23507 12789
rect -23677 12754 -23541 12755
rect -23643 12720 -23609 12754
rect -23575 12721 -23541 12754
rect -23575 12720 -23507 12721
rect -23677 12686 -23507 12720
rect -23677 12685 -23541 12686
rect -23643 12651 -23609 12685
rect -23575 12652 -23541 12685
rect -23575 12651 -23507 12652
rect -23677 12617 -23507 12651
rect -23677 12616 -23541 12617
rect -23643 12582 -23609 12616
rect -23575 12583 -23541 12616
rect -23575 12582 -23507 12583
rect -23677 12548 -23507 12582
rect -23677 12547 -23541 12548
rect -23643 12513 -23609 12547
rect -23575 12514 -23541 12547
rect -23575 12513 -23507 12514
rect -23677 12479 -23507 12513
rect -23677 12478 -23541 12479
rect -23643 12444 -23609 12478
rect -23575 12445 -23541 12478
rect -23575 12444 -23507 12445
rect -23677 12410 -23507 12444
rect -23677 12409 -23541 12410
rect -23643 12375 -23609 12409
rect -23575 12376 -23541 12409
rect -23575 12375 -23507 12376
rect -23677 12341 -23507 12375
rect -23677 12340 -23541 12341
rect -23643 12306 -23609 12340
rect -23575 12307 -23541 12340
rect -23575 12306 -23507 12307
rect -23677 12272 -23507 12306
rect -23677 12271 -23541 12272
rect -23643 12237 -23609 12271
rect -23575 12238 -23541 12271
rect -23575 12237 -23507 12238
rect -23677 12203 -23507 12237
rect -23677 12202 -23541 12203
rect -23643 12168 -23609 12202
rect -23575 12169 -23541 12202
rect -23575 12168 -23507 12169
rect -23677 12134 -23507 12168
rect -23677 12133 -23541 12134
rect -23643 12099 -23609 12133
rect -23575 12100 -23541 12133
rect -23575 12099 -23507 12100
rect -23677 12065 -23507 12099
rect -23677 12064 -23541 12065
rect -23643 12030 -23609 12064
rect -23575 12031 -23541 12064
rect -23575 12030 -23507 12031
rect -23677 11996 -23507 12030
rect -23677 11995 -23541 11996
rect -23643 11961 -23609 11995
rect -23575 11962 -23541 11995
rect -23575 11961 -23507 11962
rect -23677 11927 -23507 11961
rect -23677 11926 -23541 11927
rect -23643 11892 -23609 11926
rect -23575 11893 -23541 11926
rect -23575 11892 -23507 11893
rect -23677 11858 -23507 11892
rect -23677 11857 -23541 11858
rect -23643 11823 -23609 11857
rect -23575 11824 -23541 11857
rect -23575 11823 -23507 11824
rect -23677 11789 -23507 11823
rect -23677 11788 -23541 11789
rect -23643 11754 -23609 11788
rect -23575 11755 -23541 11788
rect -23575 11754 -23507 11755
rect -23677 11720 -23507 11754
rect -23677 11719 -23541 11720
rect -23643 11685 -23609 11719
rect -23575 11686 -23541 11719
rect -23575 11685 -23507 11686
rect -23677 11651 -23507 11685
rect -23677 11650 -23541 11651
rect -23643 11616 -23609 11650
rect -23575 11617 -23541 11650
rect -23575 11616 -23507 11617
rect -23677 11582 -23507 11616
rect -23677 11581 -23541 11582
rect -23643 11547 -23609 11581
rect -23575 11548 -23541 11581
rect -23575 11547 -23507 11548
rect -23677 11513 -23507 11547
rect -23677 11512 -23541 11513
rect -23643 11478 -23609 11512
rect -23575 11479 -23541 11512
rect -23575 11478 -23507 11479
rect -23677 11444 -23507 11478
rect -23677 11443 -23541 11444
rect -23643 11409 -23609 11443
rect -23575 11410 -23541 11443
rect -23575 11409 -23507 11410
rect -23677 11375 -23507 11409
rect -23677 11374 -23541 11375
rect -23643 11340 -23609 11374
rect -23575 11341 -23541 11374
rect -23575 11340 -23507 11341
rect -23677 11306 -23507 11340
rect -23677 11305 -23541 11306
rect -23643 11271 -23609 11305
rect -23575 11272 -23541 11305
rect -23575 11271 -23507 11272
rect -23677 11237 -23507 11271
rect -23677 11236 -23541 11237
rect -23643 11202 -23609 11236
rect -23575 11203 -23541 11236
rect -23575 11202 -23507 11203
rect -23677 11168 -23507 11202
rect -23677 11167 -23541 11168
rect -23643 11133 -23609 11167
rect -23575 11134 -23541 11167
rect -23575 11133 -23507 11134
rect -23677 11099 -23507 11133
rect -23677 11098 -23541 11099
rect -23643 11064 -23609 11098
rect -23575 11065 -23541 11098
rect -23575 11064 -23507 11065
rect -23677 11030 -23507 11064
rect -23677 11029 -23541 11030
rect -23643 10995 -23609 11029
rect -23575 10996 -23541 11029
rect -23575 10995 -23507 10996
rect -23677 10961 -23507 10995
rect -23677 10960 -23541 10961
rect -23643 10926 -23609 10960
rect -23575 10927 -23541 10960
rect -23575 10926 -23507 10927
rect -23677 10892 -23507 10926
rect -23677 10891 -23541 10892
rect -23643 10857 -23609 10891
rect -23575 10858 -23541 10891
rect -23575 10857 -23507 10858
rect -23677 10823 -23507 10857
rect -23677 10822 -23541 10823
rect -23643 10788 -23609 10822
rect -23575 10789 -23541 10822
rect -23575 10788 -23507 10789
rect -23677 10754 -23507 10788
rect -23677 10753 -23541 10754
rect -23643 10719 -23609 10753
rect -23575 10720 -23541 10753
rect -23575 10719 -23507 10720
rect -23677 10685 -23507 10719
rect -23677 10684 -23541 10685
rect -23643 10650 -23609 10684
rect -23575 10651 -23541 10684
rect -23575 10650 -23507 10651
rect -23677 10616 -23507 10650
rect -23677 10615 -23541 10616
rect -23643 10581 -23609 10615
rect -23575 10582 -23541 10615
rect -23575 10581 -23507 10582
rect -23677 10547 -23507 10581
rect -23677 10546 -23541 10547
rect -23643 10512 -23609 10546
rect -23575 10513 -23541 10546
rect -23575 10512 -23507 10513
rect -23677 10478 -23507 10512
rect -23677 10477 -23541 10478
rect -23643 10443 -23609 10477
rect -23575 10444 -23541 10477
rect -23575 10443 -23507 10444
rect -23677 10409 -23507 10443
rect -23677 10408 -23541 10409
rect -23643 10374 -23609 10408
rect -23575 10375 -23541 10408
rect -23575 10374 -23507 10375
rect -23677 10340 -23507 10374
rect -23677 10339 -23541 10340
rect -23643 10305 -23609 10339
rect -23575 10306 -23541 10339
rect -23575 10305 -23507 10306
rect -23677 10271 -23507 10305
rect -23677 10270 -23541 10271
rect -23643 10236 -23609 10270
rect -23575 10237 -23541 10270
rect -23575 10236 -23507 10237
rect -23677 10202 -23507 10236
rect -23677 10201 -23541 10202
rect -23643 10167 -23609 10201
rect -23575 10168 -23541 10201
rect -23575 10167 -23507 10168
rect -23677 10133 -23507 10167
rect -23677 10132 -23541 10133
rect -23643 10098 -23609 10132
rect -23575 10099 -23541 10132
rect -23575 10098 -23507 10099
rect -23677 10064 -23507 10098
rect -23677 10063 -23541 10064
rect -23643 10029 -23609 10063
rect -23575 10030 -23541 10063
rect -23575 10029 -23507 10030
rect -23677 9995 -23507 10029
rect -23677 9994 -23541 9995
rect -23643 9960 -23609 9994
rect -23575 9961 -23541 9994
rect -23575 9960 -23507 9961
rect -23677 9926 -23507 9960
rect -23677 9925 -23541 9926
rect -23643 9891 -23609 9925
rect -23575 9892 -23541 9925
rect -23575 9891 -23507 9892
rect -23677 9857 -23507 9891
rect -23677 9856 -23541 9857
rect -23575 9823 -23541 9856
rect -23575 9788 -23507 9823
rect -22236 7909 -22066 7944
rect -22202 7875 -22168 7909
rect -22134 7875 -22100 7909
rect -22236 7840 -22066 7875
rect -22202 7806 -22168 7840
rect -22134 7806 -22100 7840
rect -22236 7771 -22066 7806
rect -22202 7737 -22168 7771
rect -22134 7737 -22100 7771
rect -22236 7702 -22066 7737
rect -23507 7646 -23472 7680
rect -23438 7646 -23403 7680
rect -23369 7646 -23334 7680
rect -23300 7646 -23265 7680
rect -23231 7646 -23196 7680
rect -23162 7646 -23127 7680
rect -23093 7646 -23058 7680
rect -23024 7646 -22989 7680
rect -22955 7646 -22920 7680
rect -22886 7646 -22851 7680
rect -22817 7646 -22782 7680
rect -22748 7646 -22713 7680
rect -22679 7646 -22644 7680
rect -23575 7612 -22644 7646
rect -22270 7668 -22236 7680
rect -22202 7668 -22168 7702
rect -22134 7668 -22100 7702
rect -22270 7633 -22066 7668
rect -23575 7578 -23540 7612
rect -23506 7578 -23471 7612
rect -23437 7578 -23402 7612
rect -23368 7578 -23333 7612
rect -23299 7578 -23264 7612
rect -23230 7578 -23195 7612
rect -23161 7578 -23126 7612
rect -23092 7578 -23057 7612
rect -23023 7578 -22988 7612
rect -22954 7578 -22919 7612
rect -22885 7578 -22850 7612
rect -22816 7578 -22781 7612
rect -22747 7578 -22712 7612
rect -23677 7544 -22712 7578
rect -23677 7510 -23609 7544
rect -23575 7510 -23540 7544
rect -23506 7510 -23471 7544
rect -23437 7510 -23402 7544
rect -23368 7510 -23333 7544
rect -23299 7510 -23264 7544
rect -23230 7510 -23195 7544
rect -23161 7510 -23126 7544
rect -23092 7510 -23057 7544
rect -23023 7510 -22988 7544
rect -22954 7510 -22919 7544
rect -22885 7510 -22850 7544
rect -22816 7510 -22781 7544
rect -22747 7510 -22712 7544
rect -22270 7599 -22236 7633
rect -22202 7599 -22168 7633
rect -22134 7599 -22100 7633
rect -22270 7564 -22066 7599
rect -22270 7530 -22236 7564
rect -22202 7530 -22168 7564
rect -22134 7530 -22100 7564
rect -22270 7510 -22066 7530
rect -22236 7495 -22066 7510
rect -22202 7461 -22168 7495
rect -22134 7461 -22100 7495
rect -22236 7426 -22066 7461
rect -22202 7392 -22168 7426
rect -22134 7392 -22100 7426
rect -22236 7357 -22066 7392
rect -22202 7323 -22168 7357
rect -22134 7323 -22100 7357
rect -22236 7288 -22066 7323
rect -22202 7254 -22168 7288
rect -22134 7254 -22100 7288
rect -22236 7219 -22066 7254
rect -22202 7185 -22168 7219
rect -22134 7185 -22100 7219
rect -22236 7150 -22066 7185
rect -22202 7116 -22168 7150
rect -22134 7116 -22100 7150
rect -22236 7082 -22066 7116
<< psubdiffcont >>
rect -23279 14122 -23245 14156
rect -23355 8002 -23253 14088
rect -23139 14054 -22697 14156
rect -22663 14041 -22629 14075
rect -23355 7934 -23321 7968
rect -23287 7853 -22777 7955
rect -22731 7921 -22629 14007
rect -22743 7853 -22709 7887
<< mvnsubdiffcont >>
rect -22236 14478 -22066 16886
rect -23677 14376 -23643 14410
rect -23609 14376 -23167 14478
rect -23132 14444 -23098 14478
rect -23063 14444 -23029 14478
rect -22994 14444 -22960 14478
rect -22925 14444 -22891 14478
rect -22856 14444 -22822 14478
rect -22787 14444 -22753 14478
rect -22718 14444 -22684 14478
rect -22649 14444 -22615 14478
rect -22580 14444 -22546 14478
rect -22511 14444 -22477 14478
rect -22442 14444 -22408 14478
rect -22373 14444 -22339 14478
rect -23132 14376 -23098 14410
rect -23063 14376 -23029 14410
rect -22994 14376 -22960 14410
rect -22925 14376 -22891 14410
rect -22856 14376 -22822 14410
rect -22787 14376 -22753 14410
rect -22718 14376 -22684 14410
rect -22649 14376 -22615 14410
rect -22580 14376 -22546 14410
rect -22511 14376 -22477 14410
rect -22442 14376 -22408 14410
rect -22373 14376 -22339 14410
rect -23677 14307 -23643 14341
rect -23609 14307 -23575 14341
rect -23541 14308 -23167 14376
rect -23132 14308 -23098 14342
rect -23063 14308 -23029 14342
rect -22994 14308 -22960 14342
rect -22925 14308 -22891 14342
rect -22856 14308 -22822 14342
rect -22787 14308 -22753 14342
rect -22718 14308 -22684 14342
rect -22649 14308 -22615 14342
rect -22580 14308 -22546 14342
rect -22511 14308 -22477 14342
rect -22442 14308 -22408 14342
rect -22373 14308 -22339 14342
rect -22304 14308 -22066 14478
rect -23677 14238 -23643 14272
rect -23609 14238 -23575 14272
rect -23541 14239 -23507 14273
rect -23677 14169 -23643 14203
rect -23609 14169 -23575 14203
rect -23541 14170 -23507 14204
rect -23677 14100 -23643 14134
rect -23609 14100 -23575 14134
rect -23541 14101 -23507 14135
rect -23677 14031 -23643 14065
rect -23609 14031 -23575 14065
rect -23541 14032 -23507 14066
rect -23677 13962 -23643 13996
rect -23609 13962 -23575 13996
rect -23541 13963 -23507 13997
rect -23677 13893 -23643 13927
rect -23609 13893 -23575 13927
rect -23541 13894 -23507 13928
rect -23677 13824 -23643 13858
rect -23609 13824 -23575 13858
rect -23541 13825 -23507 13859
rect -23677 13755 -23643 13789
rect -23609 13755 -23575 13789
rect -23541 13756 -23507 13790
rect -23677 13686 -23643 13720
rect -23609 13686 -23575 13720
rect -23541 13687 -23507 13721
rect -23677 13617 -23643 13651
rect -23609 13617 -23575 13651
rect -23541 13618 -23507 13652
rect -23677 13548 -23643 13582
rect -23609 13548 -23575 13582
rect -23541 13549 -23507 13583
rect -23677 13479 -23643 13513
rect -23609 13479 -23575 13513
rect -23541 13480 -23507 13514
rect -23677 13410 -23643 13444
rect -23609 13410 -23575 13444
rect -23541 13411 -23507 13445
rect -23677 13341 -23643 13375
rect -23609 13341 -23575 13375
rect -23541 13342 -23507 13376
rect -23677 13272 -23643 13306
rect -23609 13272 -23575 13306
rect -23541 13273 -23507 13307
rect -23677 13203 -23643 13237
rect -23609 13203 -23575 13237
rect -23541 13204 -23507 13238
rect -23677 13134 -23643 13168
rect -23609 13134 -23575 13168
rect -23541 13135 -23507 13169
rect -23677 13065 -23643 13099
rect -23609 13065 -23575 13099
rect -23541 13066 -23507 13100
rect -23677 12996 -23643 13030
rect -23609 12996 -23575 13030
rect -23541 12997 -23507 13031
rect -23677 12927 -23643 12961
rect -23609 12927 -23575 12961
rect -23541 12928 -23507 12962
rect -23677 12858 -23643 12892
rect -23609 12858 -23575 12892
rect -23541 12859 -23507 12893
rect -23677 12789 -23643 12823
rect -23609 12789 -23575 12823
rect -23541 12790 -23507 12824
rect -23677 12720 -23643 12754
rect -23609 12720 -23575 12754
rect -23541 12721 -23507 12755
rect -23677 12651 -23643 12685
rect -23609 12651 -23575 12685
rect -23541 12652 -23507 12686
rect -23677 12582 -23643 12616
rect -23609 12582 -23575 12616
rect -23541 12583 -23507 12617
rect -23677 12513 -23643 12547
rect -23609 12513 -23575 12547
rect -23541 12514 -23507 12548
rect -23677 12444 -23643 12478
rect -23609 12444 -23575 12478
rect -23541 12445 -23507 12479
rect -23677 12375 -23643 12409
rect -23609 12375 -23575 12409
rect -23541 12376 -23507 12410
rect -23677 12306 -23643 12340
rect -23609 12306 -23575 12340
rect -23541 12307 -23507 12341
rect -23677 12237 -23643 12271
rect -23609 12237 -23575 12271
rect -23541 12238 -23507 12272
rect -23677 12168 -23643 12202
rect -23609 12168 -23575 12202
rect -23541 12169 -23507 12203
rect -23677 12099 -23643 12133
rect -23609 12099 -23575 12133
rect -23541 12100 -23507 12134
rect -23677 12030 -23643 12064
rect -23609 12030 -23575 12064
rect -23541 12031 -23507 12065
rect -23677 11961 -23643 11995
rect -23609 11961 -23575 11995
rect -23541 11962 -23507 11996
rect -23677 11892 -23643 11926
rect -23609 11892 -23575 11926
rect -23541 11893 -23507 11927
rect -23677 11823 -23643 11857
rect -23609 11823 -23575 11857
rect -23541 11824 -23507 11858
rect -23677 11754 -23643 11788
rect -23609 11754 -23575 11788
rect -23541 11755 -23507 11789
rect -23677 11685 -23643 11719
rect -23609 11685 -23575 11719
rect -23541 11686 -23507 11720
rect -23677 11616 -23643 11650
rect -23609 11616 -23575 11650
rect -23541 11617 -23507 11651
rect -23677 11547 -23643 11581
rect -23609 11547 -23575 11581
rect -23541 11548 -23507 11582
rect -23677 11478 -23643 11512
rect -23609 11478 -23575 11512
rect -23541 11479 -23507 11513
rect -23677 11409 -23643 11443
rect -23609 11409 -23575 11443
rect -23541 11410 -23507 11444
rect -23677 11340 -23643 11374
rect -23609 11340 -23575 11374
rect -23541 11341 -23507 11375
rect -23677 11271 -23643 11305
rect -23609 11271 -23575 11305
rect -23541 11272 -23507 11306
rect -23677 11202 -23643 11236
rect -23609 11202 -23575 11236
rect -23541 11203 -23507 11237
rect -23677 11133 -23643 11167
rect -23609 11133 -23575 11167
rect -23541 11134 -23507 11168
rect -23677 11064 -23643 11098
rect -23609 11064 -23575 11098
rect -23541 11065 -23507 11099
rect -23677 10995 -23643 11029
rect -23609 10995 -23575 11029
rect -23541 10996 -23507 11030
rect -23677 10926 -23643 10960
rect -23609 10926 -23575 10960
rect -23541 10927 -23507 10961
rect -23677 10857 -23643 10891
rect -23609 10857 -23575 10891
rect -23541 10858 -23507 10892
rect -23677 10788 -23643 10822
rect -23609 10788 -23575 10822
rect -23541 10789 -23507 10823
rect -23677 10719 -23643 10753
rect -23609 10719 -23575 10753
rect -23541 10720 -23507 10754
rect -23677 10650 -23643 10684
rect -23609 10650 -23575 10684
rect -23541 10651 -23507 10685
rect -23677 10581 -23643 10615
rect -23609 10581 -23575 10615
rect -23541 10582 -23507 10616
rect -23677 10512 -23643 10546
rect -23609 10512 -23575 10546
rect -23541 10513 -23507 10547
rect -23677 10443 -23643 10477
rect -23609 10443 -23575 10477
rect -23541 10444 -23507 10478
rect -23677 10374 -23643 10408
rect -23609 10374 -23575 10408
rect -23541 10375 -23507 10409
rect -23677 10305 -23643 10339
rect -23609 10305 -23575 10339
rect -23541 10306 -23507 10340
rect -23677 10236 -23643 10270
rect -23609 10236 -23575 10270
rect -23541 10237 -23507 10271
rect -23677 10167 -23643 10201
rect -23609 10167 -23575 10201
rect -23541 10168 -23507 10202
rect -23677 10098 -23643 10132
rect -23609 10098 -23575 10132
rect -23541 10099 -23507 10133
rect -23677 10029 -23643 10063
rect -23609 10029 -23575 10063
rect -23541 10030 -23507 10064
rect -23677 9960 -23643 9994
rect -23609 9960 -23575 9994
rect -23541 9961 -23507 9995
rect -23677 9891 -23643 9925
rect -23609 9891 -23575 9925
rect -23541 9892 -23507 9926
rect -23677 9788 -23575 9856
rect -23541 9823 -23507 9857
rect -23677 7646 -23507 9788
rect -22236 7944 -22066 14308
rect -22236 7875 -22202 7909
rect -22168 7875 -22134 7909
rect -22100 7875 -22066 7909
rect -22236 7806 -22202 7840
rect -22168 7806 -22134 7840
rect -22100 7806 -22066 7840
rect -22236 7737 -22202 7771
rect -22168 7737 -22134 7771
rect -22100 7737 -22066 7771
rect -23472 7646 -23438 7680
rect -23403 7646 -23369 7680
rect -23334 7646 -23300 7680
rect -23265 7646 -23231 7680
rect -23196 7646 -23162 7680
rect -23127 7646 -23093 7680
rect -23058 7646 -23024 7680
rect -22989 7646 -22955 7680
rect -22920 7646 -22886 7680
rect -22851 7646 -22817 7680
rect -22782 7646 -22748 7680
rect -22713 7646 -22679 7680
rect -23677 7578 -23575 7646
rect -22644 7612 -22270 7680
rect -22236 7668 -22202 7702
rect -22168 7668 -22134 7702
rect -22100 7668 -22066 7702
rect -23540 7578 -23506 7612
rect -23471 7578 -23437 7612
rect -23402 7578 -23368 7612
rect -23333 7578 -23299 7612
rect -23264 7578 -23230 7612
rect -23195 7578 -23161 7612
rect -23126 7578 -23092 7612
rect -23057 7578 -23023 7612
rect -22988 7578 -22954 7612
rect -22919 7578 -22885 7612
rect -22850 7578 -22816 7612
rect -22781 7578 -22747 7612
rect -23609 7510 -23575 7544
rect -23540 7510 -23506 7544
rect -23471 7510 -23437 7544
rect -23402 7510 -23368 7544
rect -23333 7510 -23299 7544
rect -23264 7510 -23230 7544
rect -23195 7510 -23161 7544
rect -23126 7510 -23092 7544
rect -23057 7510 -23023 7544
rect -22988 7510 -22954 7544
rect -22919 7510 -22885 7544
rect -22850 7510 -22816 7544
rect -22781 7510 -22747 7544
rect -22712 7510 -22270 7612
rect -22236 7599 -22202 7633
rect -22168 7599 -22134 7633
rect -22100 7599 -22066 7633
rect -22236 7530 -22202 7564
rect -22168 7530 -22134 7564
rect -22100 7530 -22066 7564
rect -22236 7461 -22202 7495
rect -22168 7461 -22134 7495
rect -22100 7461 -22066 7495
rect -22236 7392 -22202 7426
rect -22168 7392 -22134 7426
rect -22100 7392 -22066 7426
rect -22236 7323 -22202 7357
rect -22168 7323 -22134 7357
rect -22100 7323 -22066 7357
rect -22236 7254 -22202 7288
rect -22168 7254 -22134 7288
rect -22100 7254 -22066 7288
rect -22236 7185 -22202 7219
rect -22168 7185 -22134 7219
rect -22100 7185 -22066 7219
rect -22236 7116 -22202 7150
rect -22168 7116 -22134 7150
rect -22100 7116 -22066 7150
<< poly >>
rect -23120 9503 -23020 9526
rect -23120 9469 -23087 9503
rect -23053 9469 -23020 9503
rect -23120 9420 -23020 9469
rect -22964 9503 -22864 9526
rect -22964 9469 -22931 9503
rect -22897 9469 -22864 9503
rect -22964 9420 -22864 9469
rect -23120 8794 -23020 8820
rect -22964 8794 -22864 8820
rect -23164 3680 -22908 3696
rect -23164 3646 -23148 3680
rect -23114 3646 -23053 3680
rect -23019 3646 -22958 3680
rect -22924 3646 -22908 3680
rect -23164 3630 -22908 3646
rect -23164 3598 -23064 3630
rect -23008 3598 -22908 3630
rect -23164 2966 -23064 2998
rect -23008 2966 -22908 2998
rect -1040 983 -934 999
rect -1040 949 -1017 983
rect -983 949 -934 983
rect -1040 911 -934 949
rect -1040 877 -1017 911
rect -983 899 -934 911
rect 1066 983 1172 999
rect 1066 949 1115 983
rect 1149 949 1172 983
rect 1066 911 1172 949
rect 1066 899 1115 911
rect -983 877 -960 899
rect -1040 843 -960 877
rect 1092 877 1115 899
rect 1149 877 1172 911
rect 1092 843 1172 877
rect -1040 839 -934 843
rect -1040 805 -1017 839
rect -983 805 -934 839
rect -1040 767 -934 805
rect -1040 733 -1017 767
rect -983 743 -934 767
rect 1066 839 1172 843
rect 1066 805 1115 839
rect 1149 805 1172 839
rect 1066 767 1172 805
rect 1066 743 1115 767
rect -983 733 -960 743
rect -1040 695 -960 733
rect -1040 661 -1017 695
rect -983 687 -960 695
rect 1092 733 1115 743
rect 1149 733 1172 767
rect 1092 695 1172 733
rect 1092 687 1115 695
rect -983 661 -934 687
rect -1040 623 -934 661
rect -1040 589 -1017 623
rect -983 589 -934 623
rect -1040 587 -934 589
rect 1066 661 1115 687
rect 1149 661 1172 695
rect 1066 623 1172 661
rect 1066 589 1115 623
rect 1149 589 1172 623
rect 1066 587 1172 589
rect -1040 551 -960 587
rect -1040 517 -1017 551
rect -983 531 -960 551
rect 1092 551 1172 587
rect 1092 531 1115 551
rect -983 517 -934 531
rect -1040 478 -934 517
rect -1040 444 -1017 478
rect -983 444 -934 478
rect -1040 431 -934 444
rect 1066 517 1115 531
rect 1149 517 1172 551
rect 1066 478 1172 517
rect 1066 444 1115 478
rect 1149 444 1172 478
rect 1066 431 1172 444
rect -1040 405 -960 431
rect -1040 371 -1017 405
rect -983 375 -960 405
rect 1092 405 1172 431
rect 1092 375 1115 405
rect -983 371 -934 375
rect -1040 332 -934 371
rect -1040 298 -1017 332
rect -983 298 -934 332
rect -1040 275 -934 298
rect 1066 371 1115 375
rect 1149 371 1172 405
rect 1066 332 1172 371
rect 1066 298 1115 332
rect 1149 298 1172 332
rect 1066 275 1172 298
rect -1040 259 -960 275
rect -1040 225 -1017 259
rect -983 225 -960 259
rect -1040 219 -960 225
rect 1092 259 1172 275
rect 1092 225 1115 259
rect 1149 225 1172 259
rect 1092 219 1172 225
rect -1040 186 -934 219
rect -1040 152 -1017 186
rect -983 152 -934 186
rect -1040 119 -934 152
rect 1066 186 1172 219
rect 1066 152 1115 186
rect 1149 152 1172 186
rect 1066 119 1172 152
<< polycont >>
rect -23087 9469 -23053 9503
rect -22931 9469 -22897 9503
rect -23148 3646 -23114 3680
rect -23053 3646 -23019 3680
rect -22958 3646 -22924 3680
rect -1017 949 -983 983
rect -1017 877 -983 911
rect 1115 949 1149 983
rect 1115 877 1149 911
rect -1017 805 -983 839
rect -1017 733 -983 767
rect 1115 805 1149 839
rect -1017 661 -983 695
rect 1115 733 1149 767
rect -1017 589 -983 623
rect 1115 661 1149 695
rect 1115 589 1149 623
rect -1017 517 -983 551
rect -1017 444 -983 478
rect 1115 517 1149 551
rect 1115 444 1149 478
rect -1017 371 -983 405
rect -1017 298 -983 332
rect 1115 371 1149 405
rect 1115 298 1149 332
rect -1017 225 -983 259
rect 1115 225 1149 259
rect -1017 152 -983 186
rect 1115 152 1149 186
<< locali >>
rect -22236 16886 -22066 16920
rect -23687 14482 -22236 14488
rect -23687 14478 -23608 14482
rect -23574 14478 -23535 14482
rect -23501 14478 -23462 14482
rect -23428 14478 -23389 14482
rect -23355 14478 -23316 14482
rect -23282 14478 -23243 14482
rect -23209 14478 -23169 14482
rect -23135 14478 -23095 14482
rect -23061 14478 -23021 14482
rect -22987 14478 -22947 14482
rect -22913 14478 -22873 14482
rect -22839 14478 -22799 14482
rect -22765 14478 -22725 14482
rect -22691 14478 -22651 14482
rect -22617 14478 -22577 14482
rect -22543 14478 -22503 14482
rect -22469 14478 -22429 14482
rect -22395 14478 -22355 14482
rect -22321 14478 -22281 14482
rect -22247 14478 -22236 14482
rect -23687 14410 -23609 14478
rect -23135 14448 -23132 14478
rect -23167 14444 -23132 14448
rect -23098 14448 -23095 14478
rect -23029 14448 -23021 14478
rect -22960 14448 -22947 14478
rect -22891 14448 -22873 14478
rect -22822 14448 -22799 14478
rect -22753 14448 -22725 14478
rect -22684 14448 -22651 14478
rect -23098 14444 -23063 14448
rect -23029 14444 -22994 14448
rect -22960 14444 -22925 14448
rect -22891 14444 -22856 14448
rect -22822 14444 -22787 14448
rect -22753 14444 -22718 14448
rect -22684 14444 -22649 14448
rect -22615 14444 -22580 14478
rect -22543 14448 -22511 14478
rect -22469 14448 -22442 14478
rect -22395 14448 -22373 14478
rect -22321 14448 -22304 14478
rect -22546 14444 -22511 14448
rect -22477 14444 -22442 14448
rect -22408 14444 -22373 14448
rect -22339 14444 -22304 14448
rect -23167 14410 -22304 14444
rect -23687 14376 -23681 14410
rect -23643 14376 -23609 14410
rect -23135 14376 -23132 14410
rect -23098 14376 -23095 14410
rect -23029 14376 -23021 14410
rect -22960 14376 -22947 14410
rect -22891 14376 -22873 14410
rect -22822 14376 -22799 14410
rect -22753 14376 -22725 14410
rect -22684 14376 -22651 14410
rect -22615 14376 -22580 14410
rect -22543 14376 -22511 14410
rect -22469 14376 -22442 14410
rect -22395 14376 -22373 14410
rect -22321 14376 -22304 14410
rect -23687 14341 -23541 14376
rect -23687 14337 -23677 14341
rect -23687 14303 -23681 14337
rect -23643 14307 -23609 14341
rect -23575 14308 -23541 14341
rect -23167 14342 -22304 14376
rect -23167 14338 -23132 14342
rect -23135 14308 -23132 14338
rect -23098 14338 -23063 14342
rect -23029 14338 -22994 14342
rect -22960 14338 -22925 14342
rect -22891 14338 -22856 14342
rect -22822 14338 -22787 14342
rect -22753 14338 -22718 14342
rect -22684 14338 -22649 14342
rect -23098 14308 -23095 14338
rect -23029 14308 -23021 14338
rect -22960 14308 -22947 14338
rect -22891 14308 -22873 14338
rect -22822 14308 -22799 14338
rect -22753 14308 -22725 14338
rect -22684 14308 -22651 14338
rect -22615 14308 -22580 14342
rect -22546 14338 -22511 14342
rect -22477 14338 -22442 14342
rect -22408 14338 -22373 14342
rect -22339 14338 -22304 14342
rect -22543 14308 -22511 14338
rect -22469 14308 -22442 14338
rect -22395 14308 -22373 14338
rect -22321 14308 -22304 14338
rect -23647 14303 -23609 14307
rect -23575 14304 -23537 14308
rect -23503 14304 -23464 14308
rect -23430 14304 -23391 14308
rect -23357 14304 -23317 14308
rect -23283 14304 -23243 14308
rect -23209 14304 -23169 14308
rect -23135 14304 -23095 14308
rect -23061 14304 -23021 14308
rect -22987 14304 -22947 14308
rect -22913 14304 -22873 14308
rect -22839 14304 -22799 14308
rect -22765 14304 -22725 14308
rect -22691 14304 -22651 14308
rect -22617 14304 -22577 14308
rect -22543 14304 -22503 14308
rect -22469 14304 -22429 14308
rect -22395 14304 -22355 14308
rect -22321 14304 -22281 14308
rect -22247 14304 -22236 14308
rect -23575 14303 -22236 14304
rect -23687 14298 -22236 14303
rect -23687 14273 -23497 14298
rect -23687 14272 -23541 14273
rect -23687 14264 -23677 14272
rect -23687 14230 -23681 14264
rect -23643 14238 -23609 14272
rect -23575 14239 -23541 14272
rect -23507 14265 -23497 14273
rect -23647 14230 -23609 14238
rect -23575 14231 -23537 14239
rect -23503 14231 -23497 14265
rect -23575 14230 -23497 14231
rect -23687 14204 -23497 14230
rect -23687 14203 -23541 14204
rect -23687 14191 -23677 14203
rect -23687 14157 -23681 14191
rect -23643 14169 -23609 14203
rect -23575 14170 -23541 14203
rect -23507 14192 -23497 14204
rect -23647 14157 -23609 14169
rect -23575 14158 -23537 14170
rect -23503 14158 -23497 14192
rect -23575 14157 -23497 14158
rect -23687 14135 -23497 14157
rect -23687 14134 -23541 14135
rect -23687 14118 -23677 14134
rect -23687 14084 -23681 14118
rect -23643 14100 -23609 14134
rect -23575 14101 -23541 14134
rect -23507 14119 -23497 14135
rect -23647 14084 -23609 14100
rect -23575 14085 -23537 14101
rect -23503 14085 -23497 14119
rect -23575 14084 -23497 14085
rect -23687 14066 -23497 14084
rect -23687 14065 -23541 14066
rect -23687 14045 -23677 14065
rect -23687 14011 -23681 14045
rect -23643 14031 -23609 14065
rect -23575 14032 -23541 14065
rect -23507 14046 -23497 14066
rect -23647 14011 -23609 14031
rect -23575 14012 -23537 14032
rect -23503 14012 -23497 14046
rect -23575 14011 -23497 14012
rect -23687 13997 -23497 14011
rect -23687 13996 -23541 13997
rect -23687 13972 -23677 13996
rect -23687 13938 -23681 13972
rect -23643 13962 -23609 13996
rect -23575 13963 -23541 13996
rect -23507 13973 -23497 13997
rect -23647 13938 -23609 13962
rect -23575 13939 -23537 13963
rect -23503 13939 -23497 13973
rect -23575 13938 -23497 13939
rect -23687 13928 -23497 13938
rect -23687 13927 -23541 13928
rect -23687 13899 -23677 13927
rect -23687 13865 -23681 13899
rect -23643 13893 -23609 13927
rect -23575 13894 -23541 13927
rect -23507 13900 -23497 13928
rect -23647 13865 -23609 13893
rect -23575 13866 -23537 13894
rect -23503 13866 -23497 13900
rect -23575 13865 -23497 13866
rect -23687 13859 -23497 13865
rect -23687 13858 -23541 13859
rect -23687 13826 -23677 13858
rect -23687 13792 -23681 13826
rect -23643 13824 -23609 13858
rect -23575 13825 -23541 13858
rect -23507 13827 -23497 13859
rect -23647 13792 -23609 13824
rect -23575 13793 -23537 13825
rect -23503 13793 -23497 13827
rect -23575 13792 -23497 13793
rect -23687 13790 -23497 13792
rect -23687 13789 -23541 13790
rect -23687 13755 -23677 13789
rect -23643 13755 -23609 13789
rect -23575 13756 -23541 13789
rect -23507 13756 -23497 13790
rect -23575 13755 -23497 13756
rect -23687 13754 -23497 13755
rect -23687 13753 -23537 13754
rect -23687 13719 -23681 13753
rect -23647 13720 -23609 13753
rect -23575 13721 -23537 13753
rect -23687 13686 -23677 13719
rect -23643 13686 -23609 13720
rect -23575 13687 -23541 13721
rect -23503 13720 -23497 13754
rect -23507 13687 -23497 13720
rect -23575 13686 -23497 13687
rect -23687 13681 -23497 13686
rect -23687 13680 -23537 13681
rect -23687 13646 -23681 13680
rect -23647 13651 -23609 13680
rect -23575 13652 -23537 13680
rect -23687 13617 -23677 13646
rect -23643 13617 -23609 13651
rect -23575 13618 -23541 13652
rect -23503 13647 -23497 13681
rect -23507 13618 -23497 13647
rect -23575 13617 -23497 13618
rect -23687 13608 -23497 13617
rect -23687 13607 -23537 13608
rect -23687 13573 -23681 13607
rect -23647 13582 -23609 13607
rect -23575 13583 -23537 13607
rect -23687 13548 -23677 13573
rect -23643 13548 -23609 13582
rect -23575 13549 -23541 13583
rect -23503 13574 -23497 13608
rect -23507 13549 -23497 13574
rect -23575 13548 -23497 13549
rect -23687 13535 -23497 13548
rect -23687 13534 -23537 13535
rect -23687 13500 -23681 13534
rect -23647 13513 -23609 13534
rect -23575 13514 -23537 13534
rect -23687 13479 -23677 13500
rect -23643 13479 -23609 13513
rect -23575 13480 -23541 13514
rect -23503 13501 -23497 13535
rect -23507 13480 -23497 13501
rect -23575 13479 -23497 13480
rect -23687 13462 -23497 13479
rect -23687 13461 -23537 13462
rect -23687 13427 -23681 13461
rect -23647 13444 -23609 13461
rect -23575 13445 -23537 13461
rect -23687 13410 -23677 13427
rect -23643 13410 -23609 13444
rect -23575 13411 -23541 13445
rect -23503 13428 -23497 13462
rect -23507 13411 -23497 13428
rect -23575 13410 -23497 13411
rect -23687 13389 -23497 13410
rect -23687 13388 -23537 13389
rect -23687 13354 -23681 13388
rect -23647 13375 -23609 13388
rect -23575 13376 -23537 13388
rect -23687 13341 -23677 13354
rect -23643 13341 -23609 13375
rect -23575 13342 -23541 13376
rect -23503 13355 -23497 13389
rect -23507 13342 -23497 13355
rect -23575 13341 -23497 13342
rect -23687 13316 -23497 13341
rect -23687 13315 -23537 13316
rect -23687 13281 -23681 13315
rect -23647 13306 -23609 13315
rect -23575 13307 -23537 13315
rect -23687 13272 -23677 13281
rect -23643 13272 -23609 13306
rect -23575 13273 -23541 13307
rect -23503 13282 -23497 13316
rect -23507 13273 -23497 13282
rect -23575 13272 -23497 13273
rect -23687 13243 -23497 13272
rect -23687 13242 -23537 13243
rect -23687 13208 -23681 13242
rect -23647 13237 -23609 13242
rect -23575 13238 -23537 13242
rect -23687 13203 -23677 13208
rect -23643 13203 -23609 13237
rect -23575 13204 -23541 13238
rect -23503 13209 -23497 13243
rect -23507 13204 -23497 13209
rect -23575 13203 -23497 13204
rect -23687 13170 -23497 13203
rect -23687 13169 -23537 13170
rect -23687 13135 -23681 13169
rect -23647 13168 -23609 13169
rect -23687 13134 -23677 13135
rect -23643 13134 -23609 13168
rect -23575 13135 -23541 13169
rect -23503 13136 -23497 13170
rect -23507 13135 -23497 13136
rect -23575 13134 -23497 13135
rect -23687 13100 -23497 13134
rect -23687 13099 -23541 13100
rect -23687 13096 -23677 13099
rect -23687 13062 -23681 13096
rect -23643 13065 -23609 13099
rect -23575 13066 -23541 13099
rect -23507 13097 -23497 13100
rect -23647 13062 -23609 13065
rect -23575 13063 -23537 13066
rect -23503 13063 -23497 13097
rect -23575 13062 -23497 13063
rect -23687 13031 -23497 13062
rect -23687 13030 -23541 13031
rect -23687 13023 -23677 13030
rect -23687 12989 -23681 13023
rect -23643 12996 -23609 13030
rect -23575 12997 -23541 13030
rect -23507 13024 -23497 13031
rect -23647 12989 -23609 12996
rect -23575 12990 -23537 12997
rect -23503 12990 -23497 13024
rect -23575 12989 -23497 12990
rect -23687 12962 -23497 12989
rect -23687 12961 -23541 12962
rect -23687 12950 -23677 12961
rect -23687 12916 -23681 12950
rect -23643 12927 -23609 12961
rect -23575 12928 -23541 12961
rect -23507 12951 -23497 12962
rect -23647 12916 -23609 12927
rect -23575 12917 -23537 12928
rect -23503 12917 -23497 12951
rect -23575 12916 -23497 12917
rect -23687 12893 -23497 12916
rect -23687 12892 -23541 12893
rect -23687 12877 -23677 12892
rect -23687 12843 -23681 12877
rect -23643 12858 -23609 12892
rect -23575 12859 -23541 12892
rect -23507 12878 -23497 12893
rect -23647 12843 -23609 12858
rect -23575 12844 -23537 12859
rect -23503 12844 -23497 12878
rect -23575 12843 -23497 12844
rect -23687 12824 -23497 12843
rect -23687 12823 -23541 12824
rect -23687 12804 -23677 12823
rect -23687 12770 -23681 12804
rect -23643 12789 -23609 12823
rect -23575 12790 -23541 12823
rect -23507 12805 -23497 12824
rect -23647 12770 -23609 12789
rect -23575 12771 -23537 12790
rect -23503 12771 -23497 12805
rect -23575 12770 -23497 12771
rect -23687 12755 -23497 12770
rect -23687 12754 -23541 12755
rect -23687 12731 -23677 12754
rect -23687 12697 -23681 12731
rect -23643 12720 -23609 12754
rect -23575 12721 -23541 12754
rect -23507 12732 -23497 12755
rect -23647 12697 -23609 12720
rect -23575 12698 -23537 12721
rect -23503 12698 -23497 12732
rect -23575 12697 -23497 12698
rect -23687 12686 -23497 12697
rect -23687 12685 -23541 12686
rect -23687 12658 -23677 12685
rect -23687 12624 -23681 12658
rect -23643 12651 -23609 12685
rect -23575 12652 -23541 12685
rect -23507 12659 -23497 12686
rect -23647 12624 -23609 12651
rect -23575 12625 -23537 12652
rect -23503 12625 -23497 12659
rect -23575 12624 -23497 12625
rect -23687 12617 -23497 12624
rect -23687 12616 -23541 12617
rect -23687 12585 -23677 12616
rect -23687 12551 -23681 12585
rect -23643 12582 -23609 12616
rect -23575 12583 -23541 12616
rect -23507 12586 -23497 12617
rect -23647 12551 -23609 12582
rect -23575 12552 -23537 12583
rect -23503 12552 -23497 12586
rect -23575 12551 -23497 12552
rect -23687 12548 -23497 12551
rect -23687 12547 -23541 12548
rect -23687 12513 -23677 12547
rect -23643 12513 -23609 12547
rect -23575 12514 -23541 12547
rect -23507 12514 -23497 12548
rect -23575 12513 -23497 12514
rect -23687 12512 -23537 12513
rect -23687 12478 -23681 12512
rect -23647 12478 -23609 12512
rect -23575 12479 -23537 12512
rect -23503 12479 -23497 12513
rect -23687 12444 -23677 12478
rect -23643 12444 -23609 12478
rect -23575 12445 -23541 12479
rect -23507 12445 -23497 12479
rect -23575 12444 -23497 12445
rect -23687 12440 -23497 12444
rect -23687 12439 -23537 12440
rect -23687 12405 -23681 12439
rect -23647 12409 -23609 12439
rect -23575 12410 -23537 12439
rect -23687 12375 -23677 12405
rect -23643 12375 -23609 12409
rect -23575 12376 -23541 12410
rect -23503 12406 -23497 12440
rect -23507 12376 -23497 12406
rect -23575 12375 -23497 12376
rect -23687 12367 -23497 12375
rect -23687 12366 -23537 12367
rect -23687 12332 -23681 12366
rect -23647 12340 -23609 12366
rect -23575 12341 -23537 12366
rect -23687 12306 -23677 12332
rect -23643 12306 -23609 12340
rect -23575 12307 -23541 12341
rect -23503 12333 -23497 12367
rect -23507 12307 -23497 12333
rect -23575 12306 -23497 12307
rect -23687 12294 -23497 12306
rect -23687 12293 -23537 12294
rect -23687 12259 -23681 12293
rect -23647 12271 -23609 12293
rect -23575 12272 -23537 12293
rect -23687 12237 -23677 12259
rect -23643 12237 -23609 12271
rect -23575 12238 -23541 12272
rect -23503 12260 -23497 12294
rect -23507 12238 -23497 12260
rect -23575 12237 -23497 12238
rect -23687 12221 -23497 12237
rect -23687 12220 -23537 12221
rect -23687 12186 -23681 12220
rect -23647 12202 -23609 12220
rect -23575 12203 -23537 12220
rect -23687 12168 -23677 12186
rect -23643 12168 -23609 12202
rect -23575 12169 -23541 12203
rect -23503 12187 -23497 12221
rect -23507 12169 -23497 12187
rect -23575 12168 -23497 12169
rect -23687 12148 -23497 12168
rect -23687 12147 -23537 12148
rect -23687 7577 -23681 12147
rect -23575 12134 -23537 12147
rect -23575 12100 -23541 12134
rect -23503 12114 -23497 12148
rect -23507 12100 -23497 12114
rect -23575 12075 -23497 12100
rect -23503 7689 -23497 12075
rect -23363 14158 -22621 14164
rect -23363 14122 -23279 14158
rect -23245 14124 -23201 14158
rect -23167 14156 -23123 14158
rect -23089 14156 -23045 14158
rect -23011 14156 -22967 14158
rect -22933 14156 -22889 14158
rect -22855 14156 -22811 14158
rect -22777 14156 -22733 14158
rect -22699 14156 -22621 14158
rect -23167 14124 -23139 14156
rect -23245 14122 -23139 14124
rect -23363 14088 -23139 14122
rect -23363 14086 -23355 14088
rect -23253 14086 -23139 14088
rect -22697 14086 -22621 14156
rect -23363 14052 -23357 14086
rect -23251 14052 -23201 14086
rect -23167 14054 -23139 14086
rect -23167 14052 -23123 14054
rect -23089 14052 -23045 14054
rect -23011 14052 -22967 14054
rect -22933 14052 -22889 14054
rect -22855 14052 -22811 14054
rect -22777 14052 -22733 14054
rect -23363 14013 -23355 14052
rect -23253 14046 -22733 14052
rect -23253 14013 -23245 14046
rect -23363 13979 -23357 14013
rect -23251 13979 -23245 14013
rect -23363 13940 -23355 13979
rect -23253 13940 -23245 13979
rect -23363 13906 -23357 13940
rect -23251 13906 -23245 13940
rect -23363 13867 -23355 13906
rect -23253 13867 -23245 13906
rect -23363 13833 -23357 13867
rect -23251 13833 -23245 13867
rect -23363 13794 -23355 13833
rect -23253 13794 -23245 13833
rect -23363 13760 -23357 13794
rect -23251 13760 -23245 13794
rect -23363 13721 -23355 13760
rect -23253 13721 -23245 13760
rect -23363 13687 -23357 13721
rect -23251 13687 -23245 13721
rect -23363 13648 -23355 13687
rect -23253 13648 -23245 13687
rect -23363 13614 -23357 13648
rect -23251 13614 -23245 13648
rect -23363 13575 -23355 13614
rect -23253 13575 -23245 13614
rect -23363 13541 -23357 13575
rect -23251 13541 -23245 13575
rect -23363 13502 -23355 13541
rect -23253 13502 -23245 13541
rect -23363 13468 -23357 13502
rect -23251 13468 -23245 13502
rect -23363 13429 -23355 13468
rect -23253 13429 -23245 13468
rect -23363 7923 -23357 13429
rect -23251 7963 -23245 13429
rect -22739 13980 -22733 14046
rect -22627 13980 -22621 14086
rect -22739 13941 -22731 13980
rect -22629 13941 -22621 13980
rect -22739 13907 -22733 13941
rect -22627 13907 -22621 13941
rect -22739 13868 -22731 13907
rect -22629 13868 -22621 13907
rect -22739 13834 -22733 13868
rect -22627 13834 -22621 13868
rect -22739 13795 -22731 13834
rect -22629 13795 -22621 13834
rect -22739 13761 -22733 13795
rect -22627 13761 -22621 13795
rect -22739 13722 -22731 13761
rect -22629 13722 -22621 13761
rect -22739 13688 -22733 13722
rect -22627 13688 -22621 13722
rect -22739 13649 -22731 13688
rect -22629 13649 -22621 13688
rect -22739 13615 -22733 13649
rect -22627 13615 -22621 13649
rect -22739 13576 -22731 13615
rect -22629 13576 -22621 13615
rect -22739 13542 -22733 13576
rect -22627 13542 -22621 13576
rect -22739 13503 -22731 13542
rect -22629 13503 -22621 13542
rect -22739 13469 -22733 13503
rect -22627 13469 -22621 13503
rect -22739 13430 -22731 13469
rect -22629 13430 -22621 13469
rect -22739 13396 -22733 13430
rect -22627 13396 -22621 13430
rect -22739 13357 -22731 13396
rect -22629 13357 -22621 13396
rect -22739 13323 -22733 13357
rect -22627 13323 -22621 13357
rect -22739 13284 -22731 13323
rect -22629 13284 -22621 13323
rect -22739 13250 -22733 13284
rect -22627 13250 -22621 13284
rect -22739 13211 -22731 13250
rect -22629 13211 -22621 13250
rect -22739 13177 -22733 13211
rect -22627 13177 -22621 13211
rect -22739 13138 -22731 13177
rect -22629 13138 -22621 13177
rect -22739 13104 -22733 13138
rect -22627 13104 -22621 13138
rect -22739 13065 -22731 13104
rect -22629 13065 -22621 13104
rect -22739 13031 -22733 13065
rect -22627 13031 -22621 13065
rect -22739 12992 -22731 13031
rect -22629 12992 -22621 13031
rect -22739 12958 -22733 12992
rect -22627 12958 -22621 12992
rect -22739 12919 -22731 12958
rect -22629 12919 -22621 12958
rect -22739 12885 -22733 12919
rect -22627 12885 -22621 12919
rect -22739 12846 -22731 12885
rect -22629 12846 -22621 12885
rect -22739 12812 -22733 12846
rect -22627 12812 -22621 12846
rect -22739 12773 -22731 12812
rect -22629 12773 -22621 12812
rect -22739 12739 -22733 12773
rect -22627 12739 -22621 12773
rect -22739 12700 -22731 12739
rect -22629 12700 -22621 12739
rect -22739 12666 -22733 12700
rect -22627 12666 -22621 12700
rect -22739 12627 -22731 12666
rect -22629 12627 -22621 12666
rect -22739 12593 -22733 12627
rect -22627 12593 -22621 12627
rect -22739 12529 -22731 12593
rect -22629 12529 -22621 12593
rect -22739 12495 -22733 12529
rect -22627 12495 -22621 12529
rect -22739 12456 -22731 12495
rect -22629 12456 -22621 12495
rect -22739 12422 -22733 12456
rect -22627 12422 -22621 12456
rect -22739 12383 -22731 12422
rect -22629 12383 -22621 12422
rect -22739 12349 -22733 12383
rect -22627 12349 -22621 12383
rect -22739 12310 -22731 12349
rect -22629 12310 -22621 12349
rect -22739 12276 -22733 12310
rect -22627 12276 -22621 12310
rect -22739 12237 -22731 12276
rect -22629 12237 -22621 12276
rect -22739 12203 -22733 12237
rect -22627 12203 -22621 12237
rect -22739 12164 -22731 12203
rect -22629 12164 -22621 12203
rect -22739 12130 -22733 12164
rect -22627 12130 -22621 12164
rect -22739 12091 -22731 12130
rect -22629 12091 -22621 12130
rect -22739 12057 -22733 12091
rect -22627 12057 -22621 12091
rect -22739 12018 -22731 12057
rect -22629 12018 -22621 12057
rect -22739 11984 -22733 12018
rect -22627 11984 -22621 12018
rect -22739 11945 -22731 11984
rect -22629 11945 -22621 11984
rect -22739 11911 -22733 11945
rect -22627 11911 -22621 11945
rect -22739 11872 -22731 11911
rect -22629 11872 -22621 11911
rect -22739 11838 -22733 11872
rect -22627 11838 -22621 11872
rect -22739 11799 -22731 11838
rect -22629 11799 -22621 11838
rect -22739 11765 -22733 11799
rect -22627 11765 -22621 11799
rect -22739 11726 -22731 11765
rect -22629 11726 -22621 11765
rect -22739 11692 -22733 11726
rect -22627 11692 -22621 11726
rect -22739 11653 -22731 11692
rect -22629 11653 -22621 11692
rect -22739 11619 -22733 11653
rect -22627 11619 -22621 11653
rect -22739 11580 -22731 11619
rect -22629 11580 -22621 11619
rect -22739 11546 -22733 11580
rect -22627 11546 -22621 11580
rect -22739 11507 -22731 11546
rect -22629 11507 -22621 11546
rect -22739 11473 -22733 11507
rect -22627 11473 -22621 11507
rect -22739 11434 -22731 11473
rect -22629 11434 -22621 11473
rect -22739 11400 -22733 11434
rect -22627 11400 -22621 11434
rect -22739 11361 -22731 11400
rect -22629 11361 -22621 11400
rect -22739 11327 -22733 11361
rect -22627 11327 -22621 11361
rect -22739 11288 -22731 11327
rect -22629 11288 -22621 11327
rect -22739 11254 -22733 11288
rect -22627 11254 -22621 11288
rect -22739 11215 -22731 11254
rect -22629 11215 -22621 11254
rect -22739 11181 -22733 11215
rect -22627 11181 -22621 11215
rect -22739 11142 -22731 11181
rect -22629 11142 -22621 11181
rect -22739 11108 -22733 11142
rect -22627 11108 -22621 11142
rect -22739 11069 -22731 11108
rect -22629 11069 -22621 11108
rect -22739 11035 -22733 11069
rect -22627 11035 -22621 11069
rect -22739 10996 -22731 11035
rect -22629 10996 -22621 11035
rect -22739 10962 -22733 10996
rect -22627 10962 -22621 10996
rect -22739 10923 -22731 10962
rect -22629 10923 -22621 10962
rect -22739 10889 -22733 10923
rect -22627 10889 -22621 10923
rect -22739 10850 -22731 10889
rect -22629 10850 -22621 10889
rect -22739 10816 -22733 10850
rect -22627 10816 -22621 10850
rect -22739 10777 -22731 10816
rect -22629 10777 -22621 10816
rect -22739 10743 -22733 10777
rect -22627 10743 -22621 10777
rect -22739 10704 -22731 10743
rect -22629 10704 -22621 10743
rect -22739 10670 -22733 10704
rect -22627 10670 -22621 10704
rect -22739 10631 -22731 10670
rect -22629 10631 -22621 10670
rect -22739 10597 -22733 10631
rect -22627 10597 -22621 10631
rect -22739 10558 -22731 10597
rect -22629 10558 -22621 10597
rect -22739 10524 -22733 10558
rect -22627 10524 -22621 10558
rect -22739 10485 -22731 10524
rect -22629 10485 -22621 10524
rect -22739 10451 -22733 10485
rect -22627 10451 -22621 10485
rect -22739 10412 -22731 10451
rect -22629 10412 -22621 10451
rect -22739 10378 -22733 10412
rect -22627 10378 -22621 10412
rect -22739 10339 -22731 10378
rect -22629 10339 -22621 10378
rect -22739 10305 -22733 10339
rect -22627 10305 -22621 10339
rect -22739 10266 -22731 10305
rect -22629 10266 -22621 10305
rect -22739 10232 -22733 10266
rect -22627 10232 -22621 10266
rect -22739 10193 -22731 10232
rect -22629 10193 -22621 10232
rect -22739 10159 -22733 10193
rect -22627 10159 -22621 10193
rect -22739 10120 -22731 10159
rect -22629 10120 -22621 10159
rect -22739 10086 -22733 10120
rect -22627 10086 -22621 10120
rect -22739 10047 -22731 10086
rect -22629 10047 -22621 10086
rect -22739 10013 -22733 10047
rect -22627 10013 -22621 10047
rect -22739 9974 -22731 10013
rect -22629 9974 -22621 10013
rect -23103 9505 -23087 9510
rect -23053 9505 -22931 9510
rect -22897 9505 -22880 9510
rect -23103 9503 -22880 9505
rect -23103 9469 -23087 9503
rect -23053 9469 -22931 9503
rect -22897 9469 -22880 9503
rect -23103 9467 -22880 9469
rect -23103 9462 -23087 9467
rect -23053 9462 -22931 9467
rect -22897 9462 -22880 9467
rect -23165 9354 -23131 9358
rect -23165 9282 -23131 9308
rect -23165 9210 -23131 9240
rect -23165 9138 -23131 9172
rect -23165 9070 -23131 9104
rect -23165 9002 -23131 9032
rect -23165 8934 -23131 8960
rect -23165 8866 -23131 8888
rect -23009 9354 -22975 9358
rect -23009 9282 -22975 9308
rect -23009 9210 -22975 9240
rect -23009 9138 -22975 9172
rect -23009 9070 -22975 9104
rect -23009 9002 -22975 9032
rect -23009 8934 -22975 8960
rect -23009 8866 -22975 8888
rect -22853 9354 -22819 9358
rect -22853 9282 -22819 9308
rect -22853 9210 -22819 9240
rect -22853 9138 -22819 9172
rect -22853 9070 -22819 9104
rect -22853 9002 -22819 9032
rect -22853 8934 -22819 8960
rect -22853 8866 -22819 8888
rect -22739 7996 -22733 9974
rect -22627 7996 -22621 9974
rect -22739 7963 -22731 7996
rect -23251 7957 -22731 7963
rect -23251 7955 -23209 7957
rect -23175 7955 -23133 7957
rect -23099 7955 -23058 7957
rect -23024 7955 -22983 7957
rect -22949 7955 -22908 7957
rect -22874 7955 -22833 7957
rect -22799 7955 -22758 7957
rect -22777 7923 -22758 7955
rect -23363 7853 -23287 7923
rect -22777 7921 -22731 7923
rect -22629 7921 -22621 7996
rect -22777 7908 -22621 7921
rect -22777 7887 -22661 7908
rect -22777 7853 -22743 7887
rect -22709 7885 -22661 7887
rect -22705 7874 -22661 7885
rect -22627 7874 -22621 7908
rect -23363 7851 -23285 7853
rect -23251 7851 -23207 7853
rect -23173 7851 -23129 7853
rect -23095 7851 -23051 7853
rect -23017 7851 -22973 7853
rect -22939 7851 -22895 7853
rect -22861 7851 -22817 7853
rect -22783 7851 -22739 7853
rect -22705 7851 -22621 7874
rect -23363 7845 -22621 7851
rect -22236 7909 -22066 7944
rect -22202 7875 -22168 7909
rect -22134 7875 -22100 7909
rect -22236 7840 -22066 7875
rect -22202 7806 -22168 7840
rect -22134 7806 -22100 7840
rect -22236 7771 -22066 7806
rect -22202 7737 -22168 7771
rect -22134 7737 -22100 7771
rect -22236 7702 -22066 7737
rect -23503 7683 -22236 7689
rect -23503 7680 -23463 7683
rect -23429 7680 -23389 7683
rect -23355 7680 -23315 7683
rect -23281 7680 -23241 7683
rect -23207 7680 -23167 7683
rect -23133 7680 -23093 7683
rect -23503 7649 -23472 7680
rect -23429 7649 -23403 7680
rect -23355 7649 -23334 7680
rect -23281 7649 -23265 7680
rect -23207 7649 -23196 7680
rect -23133 7649 -23127 7680
rect -23507 7646 -23472 7649
rect -23438 7646 -23403 7649
rect -23369 7646 -23334 7649
rect -23300 7646 -23265 7649
rect -23231 7646 -23196 7649
rect -23162 7646 -23127 7649
rect -23059 7680 -23019 7683
rect -22985 7680 -22945 7683
rect -22911 7680 -22871 7683
rect -22837 7680 -22797 7683
rect -22763 7680 -22723 7683
rect -22689 7680 -22649 7683
rect -22615 7680 -22575 7683
rect -22541 7680 -22501 7683
rect -22467 7680 -22427 7683
rect -22393 7680 -22354 7683
rect -22320 7680 -22281 7683
rect -23059 7649 -23058 7680
rect -23093 7646 -23058 7649
rect -23024 7649 -23019 7680
rect -22955 7649 -22945 7680
rect -22886 7649 -22871 7680
rect -22817 7649 -22797 7680
rect -22748 7649 -22723 7680
rect -22679 7649 -22649 7680
rect -22247 7668 -22236 7683
rect -22202 7668 -22168 7702
rect -22134 7668 -22100 7702
rect -22247 7649 -22066 7668
rect -23024 7646 -22989 7649
rect -22955 7646 -22920 7649
rect -22886 7646 -22851 7649
rect -22817 7646 -22782 7649
rect -22748 7646 -22713 7649
rect -22679 7646 -22644 7649
rect -23575 7612 -22644 7646
rect -22270 7633 -22066 7649
rect -23575 7578 -23540 7612
rect -23506 7611 -23471 7612
rect -23437 7611 -23402 7612
rect -23368 7611 -23333 7612
rect -23299 7611 -23264 7612
rect -23230 7611 -23195 7612
rect -23161 7611 -23126 7612
rect -23501 7578 -23471 7611
rect -23427 7578 -23402 7611
rect -23353 7578 -23333 7611
rect -23279 7578 -23264 7611
rect -23205 7578 -23195 7611
rect -23131 7578 -23126 7611
rect -23092 7611 -23057 7612
rect -23092 7578 -23091 7611
rect -23575 7577 -23535 7578
rect -23501 7577 -23461 7578
rect -23427 7577 -23387 7578
rect -23353 7577 -23313 7578
rect -23279 7577 -23239 7578
rect -23205 7577 -23165 7578
rect -23131 7577 -23091 7578
rect -23023 7611 -22988 7612
rect -22954 7611 -22919 7612
rect -22885 7611 -22850 7612
rect -22816 7611 -22781 7612
rect -22747 7611 -22712 7612
rect -22270 7611 -22236 7633
rect -23023 7578 -23017 7611
rect -22954 7578 -22943 7611
rect -22885 7578 -22869 7611
rect -22816 7578 -22795 7611
rect -22747 7578 -22721 7611
rect -23057 7577 -23017 7578
rect -22983 7577 -22943 7578
rect -22909 7577 -22869 7578
rect -22835 7577 -22795 7578
rect -22761 7577 -22721 7578
rect -22247 7599 -22236 7611
rect -22202 7599 -22168 7633
rect -22134 7599 -22100 7633
rect -22247 7577 -22066 7599
rect -23687 7544 -22712 7577
rect -23687 7505 -23609 7544
rect -23575 7510 -23540 7544
rect -23506 7539 -23471 7544
rect -23437 7539 -23402 7544
rect -23368 7539 -23333 7544
rect -23299 7539 -23264 7544
rect -23230 7539 -23195 7544
rect -23161 7539 -23126 7544
rect -23501 7510 -23471 7539
rect -23427 7510 -23402 7539
rect -23353 7510 -23333 7539
rect -23279 7510 -23264 7539
rect -23205 7510 -23195 7539
rect -23131 7510 -23126 7539
rect -23092 7539 -23057 7544
rect -23092 7510 -23091 7539
rect -23575 7505 -23535 7510
rect -23501 7505 -23461 7510
rect -23427 7505 -23387 7510
rect -23353 7505 -23313 7510
rect -23279 7505 -23239 7510
rect -23205 7505 -23165 7510
rect -23131 7505 -23091 7510
rect -23023 7539 -22988 7544
rect -22954 7539 -22919 7544
rect -22885 7539 -22850 7544
rect -22816 7539 -22781 7544
rect -22747 7539 -22712 7544
rect -22270 7564 -22066 7577
rect -22270 7539 -22236 7564
rect -23023 7510 -23017 7539
rect -22954 7510 -22943 7539
rect -22885 7510 -22869 7539
rect -22816 7510 -22795 7539
rect -22747 7510 -22721 7539
rect -22247 7530 -22236 7539
rect -22202 7530 -22168 7564
rect -22134 7530 -22100 7564
rect -23057 7505 -23017 7510
rect -22983 7505 -22943 7510
rect -22909 7505 -22869 7510
rect -22835 7505 -22795 7510
rect -22761 7505 -22721 7510
rect -22687 7505 -22647 7510
rect -22613 7505 -22573 7510
rect -22539 7505 -22500 7510
rect -22466 7505 -22427 7510
rect -22393 7505 -22354 7510
rect -22320 7505 -22281 7510
rect -22247 7505 -22066 7530
rect -23687 7499 -22066 7505
rect -22236 7495 -22066 7499
rect -22202 7461 -22168 7495
rect -22134 7461 -22100 7495
rect -22236 7426 -22066 7461
rect -22202 7392 -22168 7426
rect -22134 7392 -22100 7426
rect -22236 7357 -22066 7392
rect -22202 7323 -22168 7357
rect -22134 7323 -22100 7357
rect -22236 7288 -22066 7323
rect -22202 7254 -22168 7288
rect -22134 7254 -22100 7288
rect -22236 7219 -22066 7254
rect -22202 7185 -22168 7219
rect -22134 7185 -22100 7219
rect -22236 7150 -22066 7185
rect -22202 7116 -22168 7150
rect -22134 7116 -22100 7150
rect -22236 7082 -22066 7116
rect -23164 3646 -23148 3680
rect -23114 3646 -23053 3680
rect -23019 3646 -22958 3680
rect -22924 3646 -22908 3680
rect -23209 3586 -23175 3602
rect -23209 3545 -23175 3552
rect -23209 3472 -23175 3484
rect -23209 3398 -23175 3416
rect -23209 3314 -23175 3348
rect -23209 3246 -23175 3280
rect -23209 3178 -23175 3212
rect -23209 3110 -23175 3144
rect -23209 3060 -23175 3076
rect -23053 3586 -23019 3602
rect -23053 3518 -23019 3552
rect -22897 3586 -22863 3602
rect -22897 3545 -22863 3552
rect -23053 3450 -23019 3484
rect -23053 3382 -23019 3416
rect -22884 3518 -22863 3545
rect -22918 3484 -22897 3511
rect -22918 3472 -22863 3484
rect -22884 3450 -22863 3472
rect -22918 3416 -22897 3438
rect -22918 3398 -22863 3416
rect -22884 3382 -22863 3398
rect -23053 3314 -23019 3348
rect -23053 3246 -23019 3270
rect -23053 3178 -23019 3198
rect -23053 3110 -23019 3144
rect -23053 3060 -23019 3076
rect -22897 3314 -22863 3348
rect -22897 3246 -22863 3280
rect -22897 3178 -22863 3212
rect -22897 3110 -22863 3144
rect -22897 3060 -22863 3076
rect -850 1010 -836 1044
rect -782 1010 -764 1044
rect -714 1010 -692 1044
rect -646 1010 -620 1044
rect -578 1010 -548 1044
rect -510 1010 -476 1044
rect -442 1010 -408 1044
rect -370 1010 -340 1044
rect -298 1010 -272 1044
rect -226 1010 -204 1044
rect -154 1010 -136 1044
rect -82 1010 -68 1044
rect -10 1010 0 1044
rect 62 1010 68 1044
rect 134 1010 136 1044
rect 170 1010 172 1044
rect 238 1010 244 1044
rect 306 1010 316 1044
rect 374 1010 388 1044
rect 442 1010 460 1044
rect 510 1010 532 1044
rect 578 1010 604 1044
rect 646 1010 676 1044
rect 714 1010 748 1044
rect 782 1010 816 1044
rect 854 1010 884 1044
rect 926 1010 952 1044
rect 998 1010 1020 1044
rect -1024 986 -976 999
rect -1024 949 -1017 986
rect -983 975 -976 986
rect 1108 983 1156 999
rect 1108 975 1115 983
rect -983 949 1115 975
rect 1149 975 1156 983
rect 1149 949 1158 975
rect -1024 923 1158 949
rect -1024 912 -976 923
rect -1024 877 -1017 912
rect -983 877 -976 912
rect 1108 911 1156 923
rect -1024 839 -976 877
rect -850 854 -836 888
rect -782 854 -764 888
rect -714 854 -692 888
rect -646 854 -620 888
rect -578 854 -548 888
rect -510 854 -476 888
rect -442 854 -408 888
rect -370 854 -340 888
rect -298 854 -272 888
rect -226 854 -204 888
rect -154 854 -136 888
rect -82 854 -68 888
rect -10 854 0 888
rect 62 854 68 888
rect 134 854 136 888
rect 170 854 172 888
rect 238 854 244 888
rect 306 854 316 888
rect 374 854 388 888
rect 442 854 460 888
rect 510 854 532 888
rect 578 854 604 888
rect 646 854 676 888
rect 714 854 748 888
rect 782 854 816 888
rect 854 854 884 888
rect 926 854 952 888
rect 998 854 1020 888
rect 1108 877 1115 911
rect 1149 877 1156 911
rect -1024 805 -1017 839
rect -983 819 -976 839
rect 1108 839 1156 877
rect 1108 819 1115 839
rect -983 805 1115 819
rect 1149 819 1156 839
rect 1149 805 1158 819
rect -1024 767 1158 805
rect -1024 732 -1017 767
rect -983 732 -976 767
rect 1108 733 1115 767
rect 1149 733 1156 767
rect -1024 695 -976 732
rect -850 698 -836 732
rect -782 698 -764 732
rect -714 698 -692 732
rect -646 698 -620 732
rect -578 698 -548 732
rect -510 698 -476 732
rect -442 698 -408 732
rect -370 698 -340 732
rect -298 698 -272 732
rect -226 698 -204 732
rect -154 698 -136 732
rect -82 698 -68 732
rect -10 698 0 732
rect 62 698 68 732
rect 134 698 136 732
rect 170 698 172 732
rect 238 698 244 732
rect 306 698 316 732
rect 374 698 388 732
rect 442 698 460 732
rect 510 698 532 732
rect 578 698 604 732
rect 646 698 676 732
rect 714 698 748 732
rect 782 698 816 732
rect 854 698 884 732
rect 926 698 952 732
rect 998 698 1020 732
rect -1024 659 -1017 695
rect -983 663 -976 695
rect 1108 695 1156 733
rect 1108 663 1115 695
rect -983 661 1115 663
rect 1149 663 1156 695
rect 1149 661 1158 663
rect -983 659 1158 661
rect -1024 623 1158 659
rect -1024 586 -1017 623
rect -983 611 1115 623
rect -983 586 -976 611
rect -1024 551 -976 586
rect 1108 589 1115 611
rect 1149 611 1158 623
rect 1149 589 1156 611
rect -1024 513 -1017 551
rect -983 513 -976 551
rect -850 542 -836 576
rect -782 542 -764 576
rect -714 542 -692 576
rect -646 542 -620 576
rect -578 542 -548 576
rect -510 542 -476 576
rect -442 542 -408 576
rect -370 542 -340 576
rect -298 542 -272 576
rect -226 542 -204 576
rect -154 542 -136 576
rect -82 542 -68 576
rect -10 542 0 576
rect 62 542 68 576
rect 134 542 136 576
rect 170 542 172 576
rect 238 542 244 576
rect 306 542 316 576
rect 374 542 388 576
rect 442 542 460 576
rect 510 542 532 576
rect 578 542 604 576
rect 646 542 676 576
rect 714 542 748 576
rect 782 542 816 576
rect 854 542 884 576
rect 926 542 952 576
rect 998 542 1020 576
rect 1108 551 1156 589
rect -1024 507 -976 513
rect 1108 517 1115 551
rect 1149 517 1156 551
rect 1108 507 1156 517
rect -1024 478 1158 507
rect -1024 440 -1017 478
rect -983 455 1115 478
rect -983 440 -976 455
rect -1024 405 -976 440
rect 1108 444 1115 455
rect 1149 455 1158 478
rect 1149 444 1156 455
rect -1024 367 -1017 405
rect -983 367 -976 405
rect -850 386 -836 420
rect -782 386 -764 420
rect -714 386 -692 420
rect -646 386 -620 420
rect -578 386 -548 420
rect -510 386 -476 420
rect -442 386 -408 420
rect -370 386 -340 420
rect -298 386 -272 420
rect -226 386 -204 420
rect -154 386 -136 420
rect -82 386 -68 420
rect -10 386 0 420
rect 62 386 68 420
rect 134 386 136 420
rect 170 386 172 420
rect 238 386 244 420
rect 306 386 316 420
rect 374 386 388 420
rect 442 386 460 420
rect 510 386 532 420
rect 578 386 604 420
rect 646 386 676 420
rect 714 386 748 420
rect 782 386 816 420
rect 854 386 884 420
rect 926 386 952 420
rect 998 386 1020 420
rect 1108 405 1156 444
rect -1024 351 -976 367
rect 1108 371 1115 405
rect 1149 371 1156 405
rect 1108 359 1156 371
rect 1106 351 1158 359
rect -1024 332 1158 351
rect -1024 294 -1017 332
rect -983 299 1115 332
rect -983 294 -976 299
rect -1024 259 -976 294
rect 1106 298 1115 299
rect 1149 298 1158 332
rect -1024 221 -1017 259
rect -983 221 -976 259
rect -850 230 -836 264
rect -782 230 -764 264
rect -714 230 -692 264
rect -646 230 -620 264
rect -578 230 -548 264
rect -510 230 -476 264
rect -442 230 -408 264
rect -370 230 -340 264
rect -298 230 -272 264
rect -226 230 -204 264
rect -154 230 -136 264
rect -82 230 -68 264
rect -10 230 0 264
rect 62 230 68 264
rect 134 230 136 264
rect 170 230 172 264
rect 238 230 244 264
rect 306 230 316 264
rect 374 230 388 264
rect 442 230 460 264
rect 510 230 532 264
rect 578 230 604 264
rect 646 230 676 264
rect 714 230 748 264
rect 782 230 816 264
rect 854 230 884 264
rect 926 230 952 264
rect 998 230 1020 264
rect 1106 259 1158 298
rect -1024 186 -976 221
rect 1106 225 1115 259
rect 1149 225 1158 259
rect 1106 186 1158 225
rect -1024 148 -1017 186
rect -983 148 -976 186
rect 1113 152 1115 186
rect 1149 152 1151 186
rect -1024 136 -976 148
rect 1106 136 1158 152
rect -850 74 -836 108
rect -782 74 -764 108
rect -714 74 -692 108
rect -646 74 -620 108
rect -578 74 -548 108
rect -510 74 -476 108
rect -442 74 -408 108
rect -370 74 -340 108
rect -298 74 -272 108
rect -226 74 -204 108
rect -154 74 -136 108
rect -82 74 -68 108
rect -10 74 0 108
rect 62 74 68 108
rect 134 74 136 108
rect 170 74 172 108
rect 238 74 244 108
rect 306 74 316 108
rect 374 74 388 108
rect 442 74 460 108
rect 510 74 532 108
rect 578 74 604 108
rect 646 74 676 108
rect 714 74 748 108
rect 782 74 816 108
rect 854 74 884 108
rect 926 74 952 108
rect 998 74 1020 108
<< viali >>
rect -23608 14478 -23574 14482
rect -23535 14478 -23501 14482
rect -23462 14478 -23428 14482
rect -23389 14478 -23355 14482
rect -23316 14478 -23282 14482
rect -23243 14478 -23209 14482
rect -23169 14478 -23135 14482
rect -23095 14478 -23061 14482
rect -23021 14478 -22987 14482
rect -22947 14478 -22913 14482
rect -22873 14478 -22839 14482
rect -22799 14478 -22765 14482
rect -22725 14478 -22691 14482
rect -22651 14478 -22617 14482
rect -22577 14478 -22543 14482
rect -22503 14478 -22469 14482
rect -22429 14478 -22395 14482
rect -22355 14478 -22321 14482
rect -22281 14478 -22247 14482
rect -23608 14448 -23574 14478
rect -23535 14448 -23501 14478
rect -23462 14448 -23428 14478
rect -23389 14448 -23355 14478
rect -23316 14448 -23282 14478
rect -23243 14448 -23209 14478
rect -23169 14448 -23167 14478
rect -23167 14448 -23135 14478
rect -23095 14448 -23063 14478
rect -23063 14448 -23061 14478
rect -23021 14448 -22994 14478
rect -22994 14448 -22987 14478
rect -22947 14448 -22925 14478
rect -22925 14448 -22913 14478
rect -22873 14448 -22856 14478
rect -22856 14448 -22839 14478
rect -22799 14448 -22787 14478
rect -22787 14448 -22765 14478
rect -22725 14448 -22718 14478
rect -22718 14448 -22691 14478
rect -22651 14448 -22649 14478
rect -22649 14448 -22617 14478
rect -22577 14448 -22546 14478
rect -22546 14448 -22543 14478
rect -22503 14448 -22477 14478
rect -22477 14448 -22469 14478
rect -22429 14448 -22408 14478
rect -22408 14448 -22395 14478
rect -22355 14448 -22339 14478
rect -22339 14448 -22321 14478
rect -22281 14448 -22247 14478
rect -23681 14376 -23677 14410
rect -23677 14376 -23647 14410
rect -23609 14376 -23575 14410
rect -23535 14376 -23501 14410
rect -23462 14376 -23428 14410
rect -23389 14376 -23355 14410
rect -23316 14376 -23282 14410
rect -23243 14376 -23209 14410
rect -23169 14376 -23167 14410
rect -23167 14376 -23135 14410
rect -23095 14376 -23063 14410
rect -23063 14376 -23061 14410
rect -23021 14376 -22994 14410
rect -22994 14376 -22987 14410
rect -22947 14376 -22925 14410
rect -22925 14376 -22913 14410
rect -22873 14376 -22856 14410
rect -22856 14376 -22839 14410
rect -22799 14376 -22787 14410
rect -22787 14376 -22765 14410
rect -22725 14376 -22718 14410
rect -22718 14376 -22691 14410
rect -22651 14376 -22649 14410
rect -22649 14376 -22617 14410
rect -22577 14376 -22546 14410
rect -22546 14376 -22543 14410
rect -22503 14376 -22477 14410
rect -22477 14376 -22469 14410
rect -22429 14376 -22408 14410
rect -22408 14376 -22395 14410
rect -22355 14376 -22339 14410
rect -22339 14376 -22321 14410
rect -22281 14376 -22247 14410
rect -23681 14307 -23677 14337
rect -23677 14307 -23647 14337
rect -23609 14307 -23575 14337
rect -23537 14308 -23503 14338
rect -23464 14308 -23430 14338
rect -23391 14308 -23357 14338
rect -23317 14308 -23283 14338
rect -23243 14308 -23209 14338
rect -23169 14308 -23167 14338
rect -23167 14308 -23135 14338
rect -23095 14308 -23063 14338
rect -23063 14308 -23061 14338
rect -23021 14308 -22994 14338
rect -22994 14308 -22987 14338
rect -22947 14308 -22925 14338
rect -22925 14308 -22913 14338
rect -22873 14308 -22856 14338
rect -22856 14308 -22839 14338
rect -22799 14308 -22787 14338
rect -22787 14308 -22765 14338
rect -22725 14308 -22718 14338
rect -22718 14308 -22691 14338
rect -22651 14308 -22649 14338
rect -22649 14308 -22617 14338
rect -22577 14308 -22546 14338
rect -22546 14308 -22543 14338
rect -22503 14308 -22477 14338
rect -22477 14308 -22469 14338
rect -22429 14308 -22408 14338
rect -22408 14308 -22395 14338
rect -22355 14308 -22339 14338
rect -22339 14308 -22321 14338
rect -22281 14308 -22247 14338
rect -23681 14303 -23647 14307
rect -23609 14303 -23575 14307
rect -23537 14304 -23503 14308
rect -23464 14304 -23430 14308
rect -23391 14304 -23357 14308
rect -23317 14304 -23283 14308
rect -23243 14304 -23209 14308
rect -23169 14304 -23135 14308
rect -23095 14304 -23061 14308
rect -23021 14304 -22987 14308
rect -22947 14304 -22913 14308
rect -22873 14304 -22839 14308
rect -22799 14304 -22765 14308
rect -22725 14304 -22691 14308
rect -22651 14304 -22617 14308
rect -22577 14304 -22543 14308
rect -22503 14304 -22469 14308
rect -22429 14304 -22395 14308
rect -22355 14304 -22321 14308
rect -22281 14304 -22247 14308
rect -23681 14238 -23677 14264
rect -23677 14238 -23647 14264
rect -23609 14238 -23575 14264
rect -23537 14239 -23507 14265
rect -23507 14239 -23503 14265
rect -23681 14230 -23647 14238
rect -23609 14230 -23575 14238
rect -23537 14231 -23503 14239
rect -23681 14169 -23677 14191
rect -23677 14169 -23647 14191
rect -23609 14169 -23575 14191
rect -23537 14170 -23507 14192
rect -23507 14170 -23503 14192
rect -23681 14157 -23647 14169
rect -23609 14157 -23575 14169
rect -23537 14158 -23503 14170
rect -23681 14100 -23677 14118
rect -23677 14100 -23647 14118
rect -23609 14100 -23575 14118
rect -23537 14101 -23507 14119
rect -23507 14101 -23503 14119
rect -23681 14084 -23647 14100
rect -23609 14084 -23575 14100
rect -23537 14085 -23503 14101
rect -23681 14031 -23677 14045
rect -23677 14031 -23647 14045
rect -23609 14031 -23575 14045
rect -23537 14032 -23507 14046
rect -23507 14032 -23503 14046
rect -23681 14011 -23647 14031
rect -23609 14011 -23575 14031
rect -23537 14012 -23503 14032
rect -23681 13962 -23677 13972
rect -23677 13962 -23647 13972
rect -23609 13962 -23575 13972
rect -23537 13963 -23507 13973
rect -23507 13963 -23503 13973
rect -23681 13938 -23647 13962
rect -23609 13938 -23575 13962
rect -23537 13939 -23503 13963
rect -23681 13893 -23677 13899
rect -23677 13893 -23647 13899
rect -23609 13893 -23575 13899
rect -23537 13894 -23507 13900
rect -23507 13894 -23503 13900
rect -23681 13865 -23647 13893
rect -23609 13865 -23575 13893
rect -23537 13866 -23503 13894
rect -23681 13824 -23677 13826
rect -23677 13824 -23647 13826
rect -23609 13824 -23575 13826
rect -23537 13825 -23507 13827
rect -23507 13825 -23503 13827
rect -23681 13792 -23647 13824
rect -23609 13792 -23575 13824
rect -23537 13793 -23503 13825
rect -23681 13720 -23647 13753
rect -23609 13720 -23575 13753
rect -23537 13721 -23503 13754
rect -23681 13719 -23677 13720
rect -23677 13719 -23647 13720
rect -23609 13719 -23575 13720
rect -23537 13720 -23507 13721
rect -23507 13720 -23503 13721
rect -23681 13651 -23647 13680
rect -23609 13651 -23575 13680
rect -23537 13652 -23503 13681
rect -23681 13646 -23677 13651
rect -23677 13646 -23647 13651
rect -23609 13646 -23575 13651
rect -23537 13647 -23507 13652
rect -23507 13647 -23503 13652
rect -23681 13582 -23647 13607
rect -23609 13582 -23575 13607
rect -23537 13583 -23503 13608
rect -23681 13573 -23677 13582
rect -23677 13573 -23647 13582
rect -23609 13573 -23575 13582
rect -23537 13574 -23507 13583
rect -23507 13574 -23503 13583
rect -23681 13513 -23647 13534
rect -23609 13513 -23575 13534
rect -23537 13514 -23503 13535
rect -23681 13500 -23677 13513
rect -23677 13500 -23647 13513
rect -23609 13500 -23575 13513
rect -23537 13501 -23507 13514
rect -23507 13501 -23503 13514
rect -23681 13444 -23647 13461
rect -23609 13444 -23575 13461
rect -23537 13445 -23503 13462
rect -23681 13427 -23677 13444
rect -23677 13427 -23647 13444
rect -23609 13427 -23575 13444
rect -23537 13428 -23507 13445
rect -23507 13428 -23503 13445
rect -23681 13375 -23647 13388
rect -23609 13375 -23575 13388
rect -23537 13376 -23503 13389
rect -23681 13354 -23677 13375
rect -23677 13354 -23647 13375
rect -23609 13354 -23575 13375
rect -23537 13355 -23507 13376
rect -23507 13355 -23503 13376
rect -23681 13306 -23647 13315
rect -23609 13306 -23575 13315
rect -23537 13307 -23503 13316
rect -23681 13281 -23677 13306
rect -23677 13281 -23647 13306
rect -23609 13281 -23575 13306
rect -23537 13282 -23507 13307
rect -23507 13282 -23503 13307
rect -23681 13237 -23647 13242
rect -23609 13237 -23575 13242
rect -23537 13238 -23503 13243
rect -23681 13208 -23677 13237
rect -23677 13208 -23647 13237
rect -23609 13208 -23575 13237
rect -23537 13209 -23507 13238
rect -23507 13209 -23503 13238
rect -23537 13169 -23503 13170
rect -23681 13168 -23647 13169
rect -23609 13168 -23575 13169
rect -23681 13135 -23677 13168
rect -23677 13135 -23647 13168
rect -23609 13135 -23575 13168
rect -23537 13136 -23507 13169
rect -23507 13136 -23503 13169
rect -23681 13065 -23677 13096
rect -23677 13065 -23647 13096
rect -23609 13065 -23575 13096
rect -23537 13066 -23507 13097
rect -23507 13066 -23503 13097
rect -23681 13062 -23647 13065
rect -23609 13062 -23575 13065
rect -23537 13063 -23503 13066
rect -23681 12996 -23677 13023
rect -23677 12996 -23647 13023
rect -23609 12996 -23575 13023
rect -23537 12997 -23507 13024
rect -23507 12997 -23503 13024
rect -23681 12989 -23647 12996
rect -23609 12989 -23575 12996
rect -23537 12990 -23503 12997
rect -23681 12927 -23677 12950
rect -23677 12927 -23647 12950
rect -23609 12927 -23575 12950
rect -23537 12928 -23507 12951
rect -23507 12928 -23503 12951
rect -23681 12916 -23647 12927
rect -23609 12916 -23575 12927
rect -23537 12917 -23503 12928
rect -23681 12858 -23677 12877
rect -23677 12858 -23647 12877
rect -23609 12858 -23575 12877
rect -23537 12859 -23507 12878
rect -23507 12859 -23503 12878
rect -23681 12843 -23647 12858
rect -23609 12843 -23575 12858
rect -23537 12844 -23503 12859
rect -23681 12789 -23677 12804
rect -23677 12789 -23647 12804
rect -23609 12789 -23575 12804
rect -23537 12790 -23507 12805
rect -23507 12790 -23503 12805
rect -23681 12770 -23647 12789
rect -23609 12770 -23575 12789
rect -23537 12771 -23503 12790
rect -23681 12720 -23677 12731
rect -23677 12720 -23647 12731
rect -23609 12720 -23575 12731
rect -23537 12721 -23507 12732
rect -23507 12721 -23503 12732
rect -23681 12697 -23647 12720
rect -23609 12697 -23575 12720
rect -23537 12698 -23503 12721
rect -23681 12651 -23677 12658
rect -23677 12651 -23647 12658
rect -23609 12651 -23575 12658
rect -23537 12652 -23507 12659
rect -23507 12652 -23503 12659
rect -23681 12624 -23647 12651
rect -23609 12624 -23575 12651
rect -23537 12625 -23503 12652
rect -23681 12582 -23677 12585
rect -23677 12582 -23647 12585
rect -23609 12582 -23575 12585
rect -23537 12583 -23507 12586
rect -23507 12583 -23503 12586
rect -23681 12551 -23647 12582
rect -23609 12551 -23575 12582
rect -23537 12552 -23503 12583
rect -23681 12478 -23647 12512
rect -23609 12478 -23575 12512
rect -23537 12479 -23503 12513
rect -23681 12409 -23647 12439
rect -23609 12409 -23575 12439
rect -23537 12410 -23503 12440
rect -23681 12405 -23677 12409
rect -23677 12405 -23647 12409
rect -23609 12405 -23575 12409
rect -23537 12406 -23507 12410
rect -23507 12406 -23503 12410
rect -23681 12340 -23647 12366
rect -23609 12340 -23575 12366
rect -23537 12341 -23503 12367
rect -23681 12332 -23677 12340
rect -23677 12332 -23647 12340
rect -23609 12332 -23575 12340
rect -23537 12333 -23507 12341
rect -23507 12333 -23503 12341
rect -23681 12271 -23647 12293
rect -23609 12271 -23575 12293
rect -23537 12272 -23503 12294
rect -23681 12259 -23677 12271
rect -23677 12259 -23647 12271
rect -23609 12259 -23575 12271
rect -23537 12260 -23507 12272
rect -23507 12260 -23503 12272
rect -23681 12202 -23647 12220
rect -23609 12202 -23575 12220
rect -23537 12203 -23503 12221
rect -23681 12186 -23677 12202
rect -23677 12186 -23647 12202
rect -23609 12186 -23575 12202
rect -23537 12187 -23507 12203
rect -23507 12187 -23503 12203
rect -23681 12133 -23575 12147
rect -23537 12134 -23503 12148
rect -23681 12099 -23677 12133
rect -23677 12099 -23643 12133
rect -23643 12099 -23609 12133
rect -23609 12099 -23575 12133
rect -23537 12114 -23507 12134
rect -23507 12114 -23503 12134
rect -23681 12075 -23575 12099
rect -23681 12065 -23503 12075
rect -23681 12064 -23541 12065
rect -23681 12030 -23677 12064
rect -23677 12030 -23643 12064
rect -23643 12030 -23609 12064
rect -23609 12030 -23575 12064
rect -23575 12031 -23541 12064
rect -23541 12031 -23507 12065
rect -23507 12031 -23503 12065
rect -23575 12030 -23503 12031
rect -23681 11996 -23503 12030
rect -23681 11995 -23541 11996
rect -23681 11961 -23677 11995
rect -23677 11961 -23643 11995
rect -23643 11961 -23609 11995
rect -23609 11961 -23575 11995
rect -23575 11962 -23541 11995
rect -23541 11962 -23507 11996
rect -23507 11962 -23503 11996
rect -23575 11961 -23503 11962
rect -23681 11927 -23503 11961
rect -23681 11926 -23541 11927
rect -23681 11892 -23677 11926
rect -23677 11892 -23643 11926
rect -23643 11892 -23609 11926
rect -23609 11892 -23575 11926
rect -23575 11893 -23541 11926
rect -23541 11893 -23507 11927
rect -23507 11893 -23503 11927
rect -23575 11892 -23503 11893
rect -23681 11858 -23503 11892
rect -23681 11857 -23541 11858
rect -23681 11823 -23677 11857
rect -23677 11823 -23643 11857
rect -23643 11823 -23609 11857
rect -23609 11823 -23575 11857
rect -23575 11824 -23541 11857
rect -23541 11824 -23507 11858
rect -23507 11824 -23503 11858
rect -23575 11823 -23503 11824
rect -23681 11789 -23503 11823
rect -23681 11788 -23541 11789
rect -23681 11754 -23677 11788
rect -23677 11754 -23643 11788
rect -23643 11754 -23609 11788
rect -23609 11754 -23575 11788
rect -23575 11755 -23541 11788
rect -23541 11755 -23507 11789
rect -23507 11755 -23503 11789
rect -23575 11754 -23503 11755
rect -23681 11720 -23503 11754
rect -23681 11719 -23541 11720
rect -23681 11685 -23677 11719
rect -23677 11685 -23643 11719
rect -23643 11685 -23609 11719
rect -23609 11685 -23575 11719
rect -23575 11686 -23541 11719
rect -23541 11686 -23507 11720
rect -23507 11686 -23503 11720
rect -23575 11685 -23503 11686
rect -23681 11651 -23503 11685
rect -23681 11650 -23541 11651
rect -23681 11616 -23677 11650
rect -23677 11616 -23643 11650
rect -23643 11616 -23609 11650
rect -23609 11616 -23575 11650
rect -23575 11617 -23541 11650
rect -23541 11617 -23507 11651
rect -23507 11617 -23503 11651
rect -23575 11616 -23503 11617
rect -23681 11582 -23503 11616
rect -23681 11581 -23541 11582
rect -23681 11547 -23677 11581
rect -23677 11547 -23643 11581
rect -23643 11547 -23609 11581
rect -23609 11547 -23575 11581
rect -23575 11548 -23541 11581
rect -23541 11548 -23507 11582
rect -23507 11548 -23503 11582
rect -23575 11547 -23503 11548
rect -23681 11513 -23503 11547
rect -23681 11512 -23541 11513
rect -23681 11478 -23677 11512
rect -23677 11478 -23643 11512
rect -23643 11478 -23609 11512
rect -23609 11478 -23575 11512
rect -23575 11479 -23541 11512
rect -23541 11479 -23507 11513
rect -23507 11479 -23503 11513
rect -23575 11478 -23503 11479
rect -23681 11444 -23503 11478
rect -23681 11443 -23541 11444
rect -23681 11409 -23677 11443
rect -23677 11409 -23643 11443
rect -23643 11409 -23609 11443
rect -23609 11409 -23575 11443
rect -23575 11410 -23541 11443
rect -23541 11410 -23507 11444
rect -23507 11410 -23503 11444
rect -23575 11409 -23503 11410
rect -23681 11375 -23503 11409
rect -23681 11374 -23541 11375
rect -23681 11340 -23677 11374
rect -23677 11340 -23643 11374
rect -23643 11340 -23609 11374
rect -23609 11340 -23575 11374
rect -23575 11341 -23541 11374
rect -23541 11341 -23507 11375
rect -23507 11341 -23503 11375
rect -23575 11340 -23503 11341
rect -23681 11306 -23503 11340
rect -23681 11305 -23541 11306
rect -23681 11271 -23677 11305
rect -23677 11271 -23643 11305
rect -23643 11271 -23609 11305
rect -23609 11271 -23575 11305
rect -23575 11272 -23541 11305
rect -23541 11272 -23507 11306
rect -23507 11272 -23503 11306
rect -23575 11271 -23503 11272
rect -23681 11237 -23503 11271
rect -23681 11236 -23541 11237
rect -23681 11202 -23677 11236
rect -23677 11202 -23643 11236
rect -23643 11202 -23609 11236
rect -23609 11202 -23575 11236
rect -23575 11203 -23541 11236
rect -23541 11203 -23507 11237
rect -23507 11203 -23503 11237
rect -23575 11202 -23503 11203
rect -23681 11168 -23503 11202
rect -23681 11167 -23541 11168
rect -23681 11133 -23677 11167
rect -23677 11133 -23643 11167
rect -23643 11133 -23609 11167
rect -23609 11133 -23575 11167
rect -23575 11134 -23541 11167
rect -23541 11134 -23507 11168
rect -23507 11134 -23503 11168
rect -23575 11133 -23503 11134
rect -23681 11099 -23503 11133
rect -23681 11098 -23541 11099
rect -23681 11064 -23677 11098
rect -23677 11064 -23643 11098
rect -23643 11064 -23609 11098
rect -23609 11064 -23575 11098
rect -23575 11065 -23541 11098
rect -23541 11065 -23507 11099
rect -23507 11065 -23503 11099
rect -23575 11064 -23503 11065
rect -23681 11030 -23503 11064
rect -23681 11029 -23541 11030
rect -23681 10995 -23677 11029
rect -23677 10995 -23643 11029
rect -23643 10995 -23609 11029
rect -23609 10995 -23575 11029
rect -23575 10996 -23541 11029
rect -23541 10996 -23507 11030
rect -23507 10996 -23503 11030
rect -23575 10995 -23503 10996
rect -23681 10961 -23503 10995
rect -23681 10960 -23541 10961
rect -23681 10926 -23677 10960
rect -23677 10926 -23643 10960
rect -23643 10926 -23609 10960
rect -23609 10926 -23575 10960
rect -23575 10927 -23541 10960
rect -23541 10927 -23507 10961
rect -23507 10927 -23503 10961
rect -23575 10926 -23503 10927
rect -23681 10892 -23503 10926
rect -23681 10891 -23541 10892
rect -23681 10857 -23677 10891
rect -23677 10857 -23643 10891
rect -23643 10857 -23609 10891
rect -23609 10857 -23575 10891
rect -23575 10858 -23541 10891
rect -23541 10858 -23507 10892
rect -23507 10858 -23503 10892
rect -23575 10857 -23503 10858
rect -23681 10823 -23503 10857
rect -23681 10822 -23541 10823
rect -23681 10788 -23677 10822
rect -23677 10788 -23643 10822
rect -23643 10788 -23609 10822
rect -23609 10788 -23575 10822
rect -23575 10789 -23541 10822
rect -23541 10789 -23507 10823
rect -23507 10789 -23503 10823
rect -23575 10788 -23503 10789
rect -23681 10754 -23503 10788
rect -23681 10753 -23541 10754
rect -23681 10719 -23677 10753
rect -23677 10719 -23643 10753
rect -23643 10719 -23609 10753
rect -23609 10719 -23575 10753
rect -23575 10720 -23541 10753
rect -23541 10720 -23507 10754
rect -23507 10720 -23503 10754
rect -23575 10719 -23503 10720
rect -23681 10685 -23503 10719
rect -23681 10684 -23541 10685
rect -23681 10650 -23677 10684
rect -23677 10650 -23643 10684
rect -23643 10650 -23609 10684
rect -23609 10650 -23575 10684
rect -23575 10651 -23541 10684
rect -23541 10651 -23507 10685
rect -23507 10651 -23503 10685
rect -23575 10650 -23503 10651
rect -23681 10616 -23503 10650
rect -23681 10615 -23541 10616
rect -23681 10581 -23677 10615
rect -23677 10581 -23643 10615
rect -23643 10581 -23609 10615
rect -23609 10581 -23575 10615
rect -23575 10582 -23541 10615
rect -23541 10582 -23507 10616
rect -23507 10582 -23503 10616
rect -23575 10581 -23503 10582
rect -23681 10547 -23503 10581
rect -23681 10546 -23541 10547
rect -23681 10512 -23677 10546
rect -23677 10512 -23643 10546
rect -23643 10512 -23609 10546
rect -23609 10512 -23575 10546
rect -23575 10513 -23541 10546
rect -23541 10513 -23507 10547
rect -23507 10513 -23503 10547
rect -23575 10512 -23503 10513
rect -23681 10478 -23503 10512
rect -23681 10477 -23541 10478
rect -23681 10443 -23677 10477
rect -23677 10443 -23643 10477
rect -23643 10443 -23609 10477
rect -23609 10443 -23575 10477
rect -23575 10444 -23541 10477
rect -23541 10444 -23507 10478
rect -23507 10444 -23503 10478
rect -23575 10443 -23503 10444
rect -23681 10409 -23503 10443
rect -23681 10408 -23541 10409
rect -23681 10374 -23677 10408
rect -23677 10374 -23643 10408
rect -23643 10374 -23609 10408
rect -23609 10374 -23575 10408
rect -23575 10375 -23541 10408
rect -23541 10375 -23507 10409
rect -23507 10375 -23503 10409
rect -23575 10374 -23503 10375
rect -23681 10340 -23503 10374
rect -23681 10339 -23541 10340
rect -23681 10305 -23677 10339
rect -23677 10305 -23643 10339
rect -23643 10305 -23609 10339
rect -23609 10305 -23575 10339
rect -23575 10306 -23541 10339
rect -23541 10306 -23507 10340
rect -23507 10306 -23503 10340
rect -23575 10305 -23503 10306
rect -23681 10271 -23503 10305
rect -23681 10270 -23541 10271
rect -23681 10236 -23677 10270
rect -23677 10236 -23643 10270
rect -23643 10236 -23609 10270
rect -23609 10236 -23575 10270
rect -23575 10237 -23541 10270
rect -23541 10237 -23507 10271
rect -23507 10237 -23503 10271
rect -23575 10236 -23503 10237
rect -23681 10202 -23503 10236
rect -23681 10201 -23541 10202
rect -23681 10167 -23677 10201
rect -23677 10167 -23643 10201
rect -23643 10167 -23609 10201
rect -23609 10167 -23575 10201
rect -23575 10168 -23541 10201
rect -23541 10168 -23507 10202
rect -23507 10168 -23503 10202
rect -23575 10167 -23503 10168
rect -23681 10133 -23503 10167
rect -23681 10132 -23541 10133
rect -23681 10098 -23677 10132
rect -23677 10098 -23643 10132
rect -23643 10098 -23609 10132
rect -23609 10098 -23575 10132
rect -23575 10099 -23541 10132
rect -23541 10099 -23507 10133
rect -23507 10099 -23503 10133
rect -23575 10098 -23503 10099
rect -23681 10064 -23503 10098
rect -23681 10063 -23541 10064
rect -23681 10029 -23677 10063
rect -23677 10029 -23643 10063
rect -23643 10029 -23609 10063
rect -23609 10029 -23575 10063
rect -23575 10030 -23541 10063
rect -23541 10030 -23507 10064
rect -23507 10030 -23503 10064
rect -23575 10029 -23503 10030
rect -23681 9995 -23503 10029
rect -23681 9994 -23541 9995
rect -23681 9960 -23677 9994
rect -23677 9960 -23643 9994
rect -23643 9960 -23609 9994
rect -23609 9960 -23575 9994
rect -23575 9961 -23541 9994
rect -23541 9961 -23507 9995
rect -23507 9961 -23503 9995
rect -23575 9960 -23503 9961
rect -23681 9926 -23503 9960
rect -23681 9925 -23541 9926
rect -23681 9891 -23677 9925
rect -23677 9891 -23643 9925
rect -23643 9891 -23609 9925
rect -23609 9891 -23575 9925
rect -23575 9892 -23541 9925
rect -23541 9892 -23507 9926
rect -23507 9892 -23503 9926
rect -23575 9891 -23503 9892
rect -23681 9857 -23503 9891
rect -23681 9856 -23541 9857
rect -23681 7578 -23677 9856
rect -23677 9788 -23575 9856
rect -23575 9823 -23541 9856
rect -23541 9823 -23507 9857
rect -23507 9823 -23503 9857
rect -23575 9788 -23503 9823
rect -23677 7649 -23507 9788
rect -23507 7649 -23503 9788
rect -23279 14156 -23245 14158
rect -23279 14124 -23245 14156
rect -23201 14124 -23167 14158
rect -23123 14156 -23089 14158
rect -23045 14156 -23011 14158
rect -22967 14156 -22933 14158
rect -22889 14156 -22855 14158
rect -22811 14156 -22777 14158
rect -22733 14156 -22699 14158
rect -23123 14124 -23089 14156
rect -23045 14124 -23011 14156
rect -22967 14124 -22933 14156
rect -22889 14124 -22855 14156
rect -22811 14124 -22777 14156
rect -22733 14124 -22699 14156
rect -23357 14052 -23355 14086
rect -23355 14052 -23323 14086
rect -23285 14052 -23253 14086
rect -23253 14052 -23251 14086
rect -23201 14052 -23167 14086
rect -23123 14054 -23089 14086
rect -23045 14054 -23011 14086
rect -22967 14054 -22933 14086
rect -22889 14054 -22855 14086
rect -22811 14054 -22777 14086
rect -22733 14054 -22697 14086
rect -22697 14075 -22627 14086
rect -22697 14054 -22663 14075
rect -23123 14052 -23089 14054
rect -23045 14052 -23011 14054
rect -22967 14052 -22933 14054
rect -22889 14052 -22855 14054
rect -22811 14052 -22777 14054
rect -23357 13979 -23355 14013
rect -23355 13979 -23323 14013
rect -23285 13979 -23253 14013
rect -23253 13979 -23251 14013
rect -23357 13906 -23355 13940
rect -23355 13906 -23323 13940
rect -23285 13906 -23253 13940
rect -23253 13906 -23251 13940
rect -23357 13833 -23355 13867
rect -23355 13833 -23323 13867
rect -23285 13833 -23253 13867
rect -23253 13833 -23251 13867
rect -23357 13760 -23355 13794
rect -23355 13760 -23323 13794
rect -23285 13760 -23253 13794
rect -23253 13760 -23251 13794
rect -23357 13687 -23355 13721
rect -23355 13687 -23323 13721
rect -23285 13687 -23253 13721
rect -23253 13687 -23251 13721
rect -23357 13614 -23355 13648
rect -23355 13614 -23323 13648
rect -23285 13614 -23253 13648
rect -23253 13614 -23251 13648
rect -23357 13541 -23355 13575
rect -23355 13541 -23323 13575
rect -23285 13541 -23253 13575
rect -23253 13541 -23251 13575
rect -23357 13468 -23355 13502
rect -23355 13468 -23323 13502
rect -23285 13468 -23253 13502
rect -23253 13468 -23251 13502
rect -23357 8002 -23355 13429
rect -23355 8002 -23253 13429
rect -23253 8002 -23251 13429
rect -23357 7968 -23251 8002
rect -23357 7934 -23355 7968
rect -23355 7934 -23321 7968
rect -23321 7955 -23251 7968
rect -22733 14041 -22663 14054
rect -22663 14041 -22629 14075
rect -22629 14041 -22627 14075
rect -22733 14007 -22627 14041
rect -22733 13980 -22731 14007
rect -22731 13980 -22629 14007
rect -22629 13980 -22627 14007
rect -22733 13907 -22731 13941
rect -22731 13907 -22699 13941
rect -22661 13907 -22629 13941
rect -22629 13907 -22627 13941
rect -22733 13834 -22731 13868
rect -22731 13834 -22699 13868
rect -22661 13834 -22629 13868
rect -22629 13834 -22627 13868
rect -22733 13761 -22731 13795
rect -22731 13761 -22699 13795
rect -22661 13761 -22629 13795
rect -22629 13761 -22627 13795
rect -22733 13688 -22731 13722
rect -22731 13688 -22699 13722
rect -22661 13688 -22629 13722
rect -22629 13688 -22627 13722
rect -22733 13615 -22731 13649
rect -22731 13615 -22699 13649
rect -22661 13615 -22629 13649
rect -22629 13615 -22627 13649
rect -22733 13542 -22731 13576
rect -22731 13542 -22699 13576
rect -22661 13542 -22629 13576
rect -22629 13542 -22627 13576
rect -22733 13469 -22731 13503
rect -22731 13469 -22699 13503
rect -22661 13469 -22629 13503
rect -22629 13469 -22627 13503
rect -22733 13396 -22731 13430
rect -22731 13396 -22699 13430
rect -22661 13396 -22629 13430
rect -22629 13396 -22627 13430
rect -22733 13323 -22731 13357
rect -22731 13323 -22699 13357
rect -22661 13323 -22629 13357
rect -22629 13323 -22627 13357
rect -22733 13250 -22731 13284
rect -22731 13250 -22699 13284
rect -22661 13250 -22629 13284
rect -22629 13250 -22627 13284
rect -22733 13177 -22731 13211
rect -22731 13177 -22699 13211
rect -22661 13177 -22629 13211
rect -22629 13177 -22627 13211
rect -22733 13104 -22731 13138
rect -22731 13104 -22699 13138
rect -22661 13104 -22629 13138
rect -22629 13104 -22627 13138
rect -22733 13031 -22731 13065
rect -22731 13031 -22699 13065
rect -22661 13031 -22629 13065
rect -22629 13031 -22627 13065
rect -22733 12958 -22731 12992
rect -22731 12958 -22699 12992
rect -22661 12958 -22629 12992
rect -22629 12958 -22627 12992
rect -22733 12885 -22731 12919
rect -22731 12885 -22699 12919
rect -22661 12885 -22629 12919
rect -22629 12885 -22627 12919
rect -22733 12812 -22731 12846
rect -22731 12812 -22699 12846
rect -22661 12812 -22629 12846
rect -22629 12812 -22627 12846
rect -22733 12739 -22731 12773
rect -22731 12739 -22699 12773
rect -22661 12739 -22629 12773
rect -22629 12739 -22627 12773
rect -22733 12666 -22731 12700
rect -22731 12666 -22699 12700
rect -22661 12666 -22629 12700
rect -22629 12666 -22627 12700
rect -22733 12593 -22731 12627
rect -22731 12593 -22699 12627
rect -22661 12593 -22629 12627
rect -22629 12593 -22627 12627
rect -22733 12495 -22731 12529
rect -22731 12495 -22699 12529
rect -22661 12495 -22629 12529
rect -22629 12495 -22627 12529
rect -22733 12422 -22731 12456
rect -22731 12422 -22699 12456
rect -22661 12422 -22629 12456
rect -22629 12422 -22627 12456
rect -22733 12349 -22731 12383
rect -22731 12349 -22699 12383
rect -22661 12349 -22629 12383
rect -22629 12349 -22627 12383
rect -22733 12276 -22731 12310
rect -22731 12276 -22699 12310
rect -22661 12276 -22629 12310
rect -22629 12276 -22627 12310
rect -22733 12203 -22731 12237
rect -22731 12203 -22699 12237
rect -22661 12203 -22629 12237
rect -22629 12203 -22627 12237
rect -22733 12130 -22731 12164
rect -22731 12130 -22699 12164
rect -22661 12130 -22629 12164
rect -22629 12130 -22627 12164
rect -22733 12057 -22731 12091
rect -22731 12057 -22699 12091
rect -22661 12057 -22629 12091
rect -22629 12057 -22627 12091
rect -22733 11984 -22731 12018
rect -22731 11984 -22699 12018
rect -22661 11984 -22629 12018
rect -22629 11984 -22627 12018
rect -22733 11911 -22731 11945
rect -22731 11911 -22699 11945
rect -22661 11911 -22629 11945
rect -22629 11911 -22627 11945
rect -22733 11838 -22731 11872
rect -22731 11838 -22699 11872
rect -22661 11838 -22629 11872
rect -22629 11838 -22627 11872
rect -22733 11765 -22731 11799
rect -22731 11765 -22699 11799
rect -22661 11765 -22629 11799
rect -22629 11765 -22627 11799
rect -22733 11692 -22731 11726
rect -22731 11692 -22699 11726
rect -22661 11692 -22629 11726
rect -22629 11692 -22627 11726
rect -22733 11619 -22731 11653
rect -22731 11619 -22699 11653
rect -22661 11619 -22629 11653
rect -22629 11619 -22627 11653
rect -22733 11546 -22731 11580
rect -22731 11546 -22699 11580
rect -22661 11546 -22629 11580
rect -22629 11546 -22627 11580
rect -22733 11473 -22731 11507
rect -22731 11473 -22699 11507
rect -22661 11473 -22629 11507
rect -22629 11473 -22627 11507
rect -22733 11400 -22731 11434
rect -22731 11400 -22699 11434
rect -22661 11400 -22629 11434
rect -22629 11400 -22627 11434
rect -22733 11327 -22731 11361
rect -22731 11327 -22699 11361
rect -22661 11327 -22629 11361
rect -22629 11327 -22627 11361
rect -22733 11254 -22731 11288
rect -22731 11254 -22699 11288
rect -22661 11254 -22629 11288
rect -22629 11254 -22627 11288
rect -22733 11181 -22731 11215
rect -22731 11181 -22699 11215
rect -22661 11181 -22629 11215
rect -22629 11181 -22627 11215
rect -22733 11108 -22731 11142
rect -22731 11108 -22699 11142
rect -22661 11108 -22629 11142
rect -22629 11108 -22627 11142
rect -22733 11035 -22731 11069
rect -22731 11035 -22699 11069
rect -22661 11035 -22629 11069
rect -22629 11035 -22627 11069
rect -22733 10962 -22731 10996
rect -22731 10962 -22699 10996
rect -22661 10962 -22629 10996
rect -22629 10962 -22627 10996
rect -22733 10889 -22731 10923
rect -22731 10889 -22699 10923
rect -22661 10889 -22629 10923
rect -22629 10889 -22627 10923
rect -22733 10816 -22731 10850
rect -22731 10816 -22699 10850
rect -22661 10816 -22629 10850
rect -22629 10816 -22627 10850
rect -22733 10743 -22731 10777
rect -22731 10743 -22699 10777
rect -22661 10743 -22629 10777
rect -22629 10743 -22627 10777
rect -22733 10670 -22731 10704
rect -22731 10670 -22699 10704
rect -22661 10670 -22629 10704
rect -22629 10670 -22627 10704
rect -22733 10597 -22731 10631
rect -22731 10597 -22699 10631
rect -22661 10597 -22629 10631
rect -22629 10597 -22627 10631
rect -22733 10524 -22731 10558
rect -22731 10524 -22699 10558
rect -22661 10524 -22629 10558
rect -22629 10524 -22627 10558
rect -22733 10451 -22731 10485
rect -22731 10451 -22699 10485
rect -22661 10451 -22629 10485
rect -22629 10451 -22627 10485
rect -22733 10378 -22731 10412
rect -22731 10378 -22699 10412
rect -22661 10378 -22629 10412
rect -22629 10378 -22627 10412
rect -22733 10305 -22731 10339
rect -22731 10305 -22699 10339
rect -22661 10305 -22629 10339
rect -22629 10305 -22627 10339
rect -22733 10232 -22731 10266
rect -22731 10232 -22699 10266
rect -22661 10232 -22629 10266
rect -22629 10232 -22627 10266
rect -22733 10159 -22731 10193
rect -22731 10159 -22699 10193
rect -22661 10159 -22629 10193
rect -22629 10159 -22627 10193
rect -22733 10086 -22731 10120
rect -22731 10086 -22699 10120
rect -22661 10086 -22629 10120
rect -22629 10086 -22627 10120
rect -22733 10013 -22731 10047
rect -22731 10013 -22699 10047
rect -22661 10013 -22629 10047
rect -22629 10013 -22627 10047
rect -23087 9505 -23053 9539
rect -22931 9505 -22897 9539
rect -23087 9433 -23053 9467
rect -22931 9433 -22897 9467
rect -23165 9342 -23131 9354
rect -23165 9320 -23131 9342
rect -23165 9274 -23131 9282
rect -23165 9248 -23131 9274
rect -23165 9206 -23131 9210
rect -23165 9176 -23131 9206
rect -23165 9104 -23131 9138
rect -23165 9036 -23131 9066
rect -23165 9032 -23131 9036
rect -23165 8968 -23131 8994
rect -23165 8960 -23131 8968
rect -23165 8900 -23131 8922
rect -23165 8888 -23131 8900
rect -23165 8832 -23131 8850
rect -23165 8816 -23131 8832
rect -23009 9342 -22975 9354
rect -23009 9320 -22975 9342
rect -23009 9274 -22975 9282
rect -23009 9248 -22975 9274
rect -23009 9206 -22975 9210
rect -23009 9176 -22975 9206
rect -23009 9104 -22975 9138
rect -23009 9036 -22975 9066
rect -23009 9032 -22975 9036
rect -23009 8968 -22975 8994
rect -23009 8960 -22975 8968
rect -23009 8900 -22975 8922
rect -23009 8888 -22975 8900
rect -23009 8832 -22975 8850
rect -23009 8816 -22975 8832
rect -22853 9342 -22819 9354
rect -22853 9320 -22819 9342
rect -22853 9274 -22819 9282
rect -22853 9248 -22819 9274
rect -22853 9206 -22819 9210
rect -22853 9176 -22819 9206
rect -22853 9104 -22819 9138
rect -22853 9036 -22819 9066
rect -22853 9032 -22819 9036
rect -22853 8968 -22819 8994
rect -22853 8960 -22819 8968
rect -22853 8900 -22819 8922
rect -22853 8888 -22819 8900
rect -22853 8832 -22819 8850
rect -22853 8816 -22819 8832
rect -22733 7996 -22731 9974
rect -22731 7996 -22629 9974
rect -22629 7996 -22627 9974
rect -23209 7955 -23175 7957
rect -23133 7955 -23099 7957
rect -23058 7955 -23024 7957
rect -22983 7955 -22949 7957
rect -22908 7955 -22874 7957
rect -22833 7955 -22799 7957
rect -23321 7934 -23287 7955
rect -23357 7923 -23287 7934
rect -23287 7923 -23251 7955
rect -23209 7923 -23175 7955
rect -23133 7923 -23099 7955
rect -23058 7923 -23024 7955
rect -22983 7923 -22949 7955
rect -22908 7923 -22874 7955
rect -22833 7923 -22799 7955
rect -22758 7923 -22731 7957
rect -22731 7923 -22724 7957
rect -23285 7853 -23251 7885
rect -23207 7853 -23173 7885
rect -23129 7853 -23095 7885
rect -23051 7853 -23017 7885
rect -22973 7853 -22939 7885
rect -22895 7853 -22861 7885
rect -22817 7853 -22783 7885
rect -22739 7853 -22709 7885
rect -22709 7853 -22705 7885
rect -22661 7874 -22627 7908
rect -23285 7851 -23251 7853
rect -23207 7851 -23173 7853
rect -23129 7851 -23095 7853
rect -23051 7851 -23017 7853
rect -22973 7851 -22939 7853
rect -22895 7851 -22861 7853
rect -22817 7851 -22783 7853
rect -22739 7851 -22705 7853
rect -23463 7680 -23429 7683
rect -23389 7680 -23355 7683
rect -23315 7680 -23281 7683
rect -23241 7680 -23207 7683
rect -23167 7680 -23133 7683
rect -23463 7649 -23438 7680
rect -23438 7649 -23429 7680
rect -23389 7649 -23369 7680
rect -23369 7649 -23355 7680
rect -23315 7649 -23300 7680
rect -23300 7649 -23281 7680
rect -23241 7649 -23231 7680
rect -23231 7649 -23207 7680
rect -23167 7649 -23162 7680
rect -23162 7649 -23133 7680
rect -23677 7578 -23575 7649
rect -23093 7649 -23059 7683
rect -23019 7680 -22985 7683
rect -22945 7680 -22911 7683
rect -22871 7680 -22837 7683
rect -22797 7680 -22763 7683
rect -22723 7680 -22689 7683
rect -22649 7680 -22615 7683
rect -22575 7680 -22541 7683
rect -22501 7680 -22467 7683
rect -22427 7680 -22393 7683
rect -22354 7680 -22320 7683
rect -22281 7680 -22247 7683
rect -23019 7649 -22989 7680
rect -22989 7649 -22985 7680
rect -22945 7649 -22920 7680
rect -22920 7649 -22911 7680
rect -22871 7649 -22851 7680
rect -22851 7649 -22837 7680
rect -22797 7649 -22782 7680
rect -22782 7649 -22763 7680
rect -22723 7649 -22713 7680
rect -22713 7649 -22689 7680
rect -22649 7649 -22644 7680
rect -22644 7649 -22615 7680
rect -22575 7649 -22541 7680
rect -22501 7649 -22467 7680
rect -22427 7649 -22393 7680
rect -22354 7649 -22320 7680
rect -22281 7649 -22270 7680
rect -22270 7649 -22247 7680
rect -23535 7578 -23506 7611
rect -23506 7578 -23501 7611
rect -23461 7578 -23437 7611
rect -23437 7578 -23427 7611
rect -23387 7578 -23368 7611
rect -23368 7578 -23353 7611
rect -23313 7578 -23299 7611
rect -23299 7578 -23279 7611
rect -23239 7578 -23230 7611
rect -23230 7578 -23205 7611
rect -23165 7578 -23161 7611
rect -23161 7578 -23131 7611
rect -23681 7577 -23575 7578
rect -23535 7577 -23501 7578
rect -23461 7577 -23427 7578
rect -23387 7577 -23353 7578
rect -23313 7577 -23279 7578
rect -23239 7577 -23205 7578
rect -23165 7577 -23131 7578
rect -23091 7577 -23057 7611
rect -23017 7578 -22988 7611
rect -22988 7578 -22983 7611
rect -22943 7578 -22919 7611
rect -22919 7578 -22909 7611
rect -22869 7578 -22850 7611
rect -22850 7578 -22835 7611
rect -22795 7578 -22781 7611
rect -22781 7578 -22761 7611
rect -23017 7577 -22983 7578
rect -22943 7577 -22909 7578
rect -22869 7577 -22835 7578
rect -22795 7577 -22761 7578
rect -22721 7577 -22712 7611
rect -22712 7577 -22687 7611
rect -22647 7577 -22613 7611
rect -22573 7577 -22539 7611
rect -22500 7577 -22466 7611
rect -22427 7577 -22393 7611
rect -22354 7577 -22320 7611
rect -22281 7577 -22270 7611
rect -22270 7577 -22247 7611
rect -23609 7510 -23575 7539
rect -23535 7510 -23506 7539
rect -23506 7510 -23501 7539
rect -23461 7510 -23437 7539
rect -23437 7510 -23427 7539
rect -23387 7510 -23368 7539
rect -23368 7510 -23353 7539
rect -23313 7510 -23299 7539
rect -23299 7510 -23279 7539
rect -23239 7510 -23230 7539
rect -23230 7510 -23205 7539
rect -23165 7510 -23161 7539
rect -23161 7510 -23131 7539
rect -23609 7505 -23575 7510
rect -23535 7505 -23501 7510
rect -23461 7505 -23427 7510
rect -23387 7505 -23353 7510
rect -23313 7505 -23279 7510
rect -23239 7505 -23205 7510
rect -23165 7505 -23131 7510
rect -23091 7505 -23057 7539
rect -23017 7510 -22988 7539
rect -22988 7510 -22983 7539
rect -22943 7510 -22919 7539
rect -22919 7510 -22909 7539
rect -22869 7510 -22850 7539
rect -22850 7510 -22835 7539
rect -22795 7510 -22781 7539
rect -22781 7510 -22761 7539
rect -22721 7510 -22712 7539
rect -22712 7510 -22687 7539
rect -22647 7510 -22613 7539
rect -22573 7510 -22539 7539
rect -22500 7510 -22466 7539
rect -22427 7510 -22393 7539
rect -22354 7510 -22320 7539
rect -22281 7510 -22270 7539
rect -22270 7510 -22247 7539
rect -23017 7505 -22983 7510
rect -22943 7505 -22909 7510
rect -22869 7505 -22835 7510
rect -22795 7505 -22761 7510
rect -22721 7505 -22687 7510
rect -22647 7505 -22613 7510
rect -22573 7505 -22539 7510
rect -22500 7505 -22466 7510
rect -22427 7505 -22393 7510
rect -22354 7505 -22320 7510
rect -22281 7505 -22247 7510
rect -23209 3518 -23175 3545
rect -23209 3511 -23175 3518
rect -23209 3450 -23175 3472
rect -23209 3438 -23175 3450
rect -23209 3382 -23175 3398
rect -23209 3364 -23175 3382
rect -22918 3518 -22884 3545
rect -22918 3511 -22897 3518
rect -22897 3511 -22884 3518
rect -22918 3450 -22884 3472
rect -22918 3438 -22897 3450
rect -22897 3438 -22884 3450
rect -22918 3382 -22884 3398
rect -22918 3364 -22897 3382
rect -22897 3364 -22884 3382
rect -23053 3280 -23019 3304
rect -23053 3270 -23019 3280
rect -23053 3212 -23019 3232
rect -23053 3198 -23019 3212
rect -908 1010 -884 1044
rect -884 1010 -874 1044
rect -836 1010 -816 1044
rect -816 1010 -802 1044
rect -764 1010 -748 1044
rect -748 1010 -730 1044
rect -692 1010 -680 1044
rect -680 1010 -658 1044
rect -620 1010 -612 1044
rect -612 1010 -586 1044
rect -548 1010 -544 1044
rect -544 1010 -514 1044
rect -476 1010 -442 1044
rect -404 1010 -374 1044
rect -374 1010 -370 1044
rect -332 1010 -306 1044
rect -306 1010 -298 1044
rect -260 1010 -238 1044
rect -238 1010 -226 1044
rect -188 1010 -170 1044
rect -170 1010 -154 1044
rect -116 1010 -102 1044
rect -102 1010 -82 1044
rect -44 1010 -34 1044
rect -34 1010 -10 1044
rect 28 1010 34 1044
rect 34 1010 62 1044
rect 100 1010 102 1044
rect 102 1010 134 1044
rect 172 1010 204 1044
rect 204 1010 206 1044
rect 244 1010 272 1044
rect 272 1010 278 1044
rect 316 1010 340 1044
rect 340 1010 350 1044
rect 388 1010 408 1044
rect 408 1010 422 1044
rect 460 1010 476 1044
rect 476 1010 494 1044
rect 532 1010 544 1044
rect 544 1010 566 1044
rect 604 1010 612 1044
rect 612 1010 638 1044
rect 676 1010 680 1044
rect 680 1010 710 1044
rect 748 1010 782 1044
rect 820 1010 850 1044
rect 850 1010 854 1044
rect 892 1010 918 1044
rect 918 1010 926 1044
rect 964 1010 986 1044
rect 986 1010 998 1044
rect 1036 1010 1054 1044
rect 1054 1010 1070 1044
rect -1017 983 -983 986
rect -1017 952 -983 983
rect -1017 911 -983 912
rect -1017 878 -983 911
rect -908 854 -884 888
rect -884 854 -874 888
rect -836 854 -816 888
rect -816 854 -802 888
rect -764 854 -748 888
rect -748 854 -730 888
rect -692 854 -680 888
rect -680 854 -658 888
rect -620 854 -612 888
rect -612 854 -586 888
rect -548 854 -544 888
rect -544 854 -514 888
rect -476 854 -442 888
rect -404 854 -374 888
rect -374 854 -370 888
rect -332 854 -306 888
rect -306 854 -298 888
rect -260 854 -238 888
rect -238 854 -226 888
rect -188 854 -170 888
rect -170 854 -154 888
rect -116 854 -102 888
rect -102 854 -82 888
rect -44 854 -34 888
rect -34 854 -10 888
rect 28 854 34 888
rect 34 854 62 888
rect 100 854 102 888
rect 102 854 134 888
rect 172 854 204 888
rect 204 854 206 888
rect 244 854 272 888
rect 272 854 278 888
rect 316 854 340 888
rect 340 854 350 888
rect 388 854 408 888
rect 408 854 422 888
rect 460 854 476 888
rect 476 854 494 888
rect 532 854 544 888
rect 544 854 566 888
rect 604 854 612 888
rect 612 854 638 888
rect 676 854 680 888
rect 680 854 710 888
rect 748 854 782 888
rect 820 854 850 888
rect 850 854 854 888
rect 892 854 918 888
rect 918 854 926 888
rect 964 854 986 888
rect 986 854 998 888
rect 1036 854 1054 888
rect 1054 854 1070 888
rect -1017 805 -983 839
rect -1017 733 -983 766
rect -1017 732 -983 733
rect -908 698 -884 732
rect -884 698 -874 732
rect -836 698 -816 732
rect -816 698 -802 732
rect -764 698 -748 732
rect -748 698 -730 732
rect -692 698 -680 732
rect -680 698 -658 732
rect -620 698 -612 732
rect -612 698 -586 732
rect -548 698 -544 732
rect -544 698 -514 732
rect -476 698 -442 732
rect -404 698 -374 732
rect -374 698 -370 732
rect -332 698 -306 732
rect -306 698 -298 732
rect -260 698 -238 732
rect -238 698 -226 732
rect -188 698 -170 732
rect -170 698 -154 732
rect -116 698 -102 732
rect -102 698 -82 732
rect -44 698 -34 732
rect -34 698 -10 732
rect 28 698 34 732
rect 34 698 62 732
rect 100 698 102 732
rect 102 698 134 732
rect 172 698 204 732
rect 204 698 206 732
rect 244 698 272 732
rect 272 698 278 732
rect 316 698 340 732
rect 340 698 350 732
rect 388 698 408 732
rect 408 698 422 732
rect 460 698 476 732
rect 476 698 494 732
rect 532 698 544 732
rect 544 698 566 732
rect 604 698 612 732
rect 612 698 638 732
rect 676 698 680 732
rect 680 698 710 732
rect 748 698 782 732
rect 820 698 850 732
rect 850 698 854 732
rect 892 698 918 732
rect 918 698 926 732
rect 964 698 986 732
rect 986 698 998 732
rect 1036 698 1054 732
rect 1054 698 1070 732
rect -1017 661 -983 693
rect -1017 659 -983 661
rect -1017 589 -983 620
rect -1017 586 -983 589
rect -1017 517 -983 547
rect -1017 513 -983 517
rect -908 542 -884 576
rect -884 542 -874 576
rect -836 542 -816 576
rect -816 542 -802 576
rect -764 542 -748 576
rect -748 542 -730 576
rect -692 542 -680 576
rect -680 542 -658 576
rect -620 542 -612 576
rect -612 542 -586 576
rect -548 542 -544 576
rect -544 542 -514 576
rect -476 542 -442 576
rect -404 542 -374 576
rect -374 542 -370 576
rect -332 542 -306 576
rect -306 542 -298 576
rect -260 542 -238 576
rect -238 542 -226 576
rect -188 542 -170 576
rect -170 542 -154 576
rect -116 542 -102 576
rect -102 542 -82 576
rect -44 542 -34 576
rect -34 542 -10 576
rect 28 542 34 576
rect 34 542 62 576
rect 100 542 102 576
rect 102 542 134 576
rect 172 542 204 576
rect 204 542 206 576
rect 244 542 272 576
rect 272 542 278 576
rect 316 542 340 576
rect 340 542 350 576
rect 388 542 408 576
rect 408 542 422 576
rect 460 542 476 576
rect 476 542 494 576
rect 532 542 544 576
rect 544 542 566 576
rect 604 542 612 576
rect 612 542 638 576
rect 676 542 680 576
rect 680 542 710 576
rect 748 542 782 576
rect 820 542 850 576
rect 850 542 854 576
rect 892 542 918 576
rect 918 542 926 576
rect 964 542 986 576
rect 986 542 998 576
rect 1036 542 1054 576
rect 1054 542 1070 576
rect -1017 444 -983 474
rect -1017 440 -983 444
rect -1017 371 -983 401
rect -1017 367 -983 371
rect -908 386 -884 420
rect -884 386 -874 420
rect -836 386 -816 420
rect -816 386 -802 420
rect -764 386 -748 420
rect -748 386 -730 420
rect -692 386 -680 420
rect -680 386 -658 420
rect -620 386 -612 420
rect -612 386 -586 420
rect -548 386 -544 420
rect -544 386 -514 420
rect -476 386 -442 420
rect -404 386 -374 420
rect -374 386 -370 420
rect -332 386 -306 420
rect -306 386 -298 420
rect -260 386 -238 420
rect -238 386 -226 420
rect -188 386 -170 420
rect -170 386 -154 420
rect -116 386 -102 420
rect -102 386 -82 420
rect -44 386 -34 420
rect -34 386 -10 420
rect 28 386 34 420
rect 34 386 62 420
rect 100 386 102 420
rect 102 386 134 420
rect 172 386 204 420
rect 204 386 206 420
rect 244 386 272 420
rect 272 386 278 420
rect 316 386 340 420
rect 340 386 350 420
rect 388 386 408 420
rect 408 386 422 420
rect 460 386 476 420
rect 476 386 494 420
rect 532 386 544 420
rect 544 386 566 420
rect 604 386 612 420
rect 612 386 638 420
rect 676 386 680 420
rect 680 386 710 420
rect 748 386 782 420
rect 820 386 850 420
rect 850 386 854 420
rect 892 386 918 420
rect 918 386 926 420
rect 964 386 986 420
rect 986 386 998 420
rect 1036 386 1054 420
rect 1054 386 1070 420
rect -1017 298 -983 328
rect -1017 294 -983 298
rect -1017 225 -983 255
rect -1017 221 -983 225
rect -908 230 -884 264
rect -884 230 -874 264
rect -836 230 -816 264
rect -816 230 -802 264
rect -764 230 -748 264
rect -748 230 -730 264
rect -692 230 -680 264
rect -680 230 -658 264
rect -620 230 -612 264
rect -612 230 -586 264
rect -548 230 -544 264
rect -544 230 -514 264
rect -476 230 -442 264
rect -404 230 -374 264
rect -374 230 -370 264
rect -332 230 -306 264
rect -306 230 -298 264
rect -260 230 -238 264
rect -238 230 -226 264
rect -188 230 -170 264
rect -170 230 -154 264
rect -116 230 -102 264
rect -102 230 -82 264
rect -44 230 -34 264
rect -34 230 -10 264
rect 28 230 34 264
rect 34 230 62 264
rect 100 230 102 264
rect 102 230 134 264
rect 172 230 204 264
rect 204 230 206 264
rect 244 230 272 264
rect 272 230 278 264
rect 316 230 340 264
rect 340 230 350 264
rect 388 230 408 264
rect 408 230 422 264
rect 460 230 476 264
rect 476 230 494 264
rect 532 230 544 264
rect 544 230 566 264
rect 604 230 612 264
rect 612 230 638 264
rect 676 230 680 264
rect 680 230 710 264
rect 748 230 782 264
rect 820 230 850 264
rect 850 230 854 264
rect 892 230 918 264
rect 918 230 926 264
rect 964 230 986 264
rect 986 230 998 264
rect 1036 230 1054 264
rect 1054 230 1070 264
rect -1017 152 -983 182
rect -1017 148 -983 152
rect 1079 152 1113 186
rect 1151 152 1185 186
rect -908 74 -884 108
rect -884 74 -874 108
rect -836 74 -816 108
rect -816 74 -802 108
rect -764 74 -748 108
rect -748 74 -730 108
rect -692 74 -680 108
rect -680 74 -658 108
rect -620 74 -612 108
rect -612 74 -586 108
rect -548 74 -544 108
rect -544 74 -514 108
rect -476 74 -442 108
rect -404 74 -374 108
rect -374 74 -370 108
rect -332 74 -306 108
rect -306 74 -298 108
rect -260 74 -238 108
rect -238 74 -226 108
rect -188 74 -170 108
rect -170 74 -154 108
rect -116 74 -102 108
rect -102 74 -82 108
rect -44 74 -34 108
rect -34 74 -10 108
rect 28 74 34 108
rect 34 74 62 108
rect 100 74 102 108
rect 102 74 134 108
rect 172 74 204 108
rect 204 74 206 108
rect 244 74 272 108
rect 272 74 278 108
rect 316 74 340 108
rect 340 74 350 108
rect 388 74 408 108
rect 408 74 422 108
rect 460 74 476 108
rect 476 74 494 108
rect 532 74 544 108
rect 544 74 566 108
rect 604 74 612 108
rect 612 74 638 108
rect 676 74 680 108
rect 680 74 710 108
rect 748 74 782 108
rect 820 74 850 108
rect 850 74 854 108
rect 892 74 918 108
rect 918 74 926 108
rect 964 74 986 108
rect 986 74 998 108
rect 1036 74 1054 108
rect 1054 74 1070 108
<< metal1 >>
rect -23687 14482 -22215 14488
rect -23687 14448 -23608 14482
rect -23574 14448 -23535 14482
rect -23501 14448 -23462 14482
rect -23428 14448 -23389 14482
rect -23355 14448 -23316 14482
rect -23282 14448 -23243 14482
rect -23209 14448 -23169 14482
rect -23135 14448 -23095 14482
rect -23061 14448 -23021 14482
rect -22987 14448 -22947 14482
rect -22913 14448 -22873 14482
rect -22839 14448 -22799 14482
rect -22765 14448 -22725 14482
rect -22691 14448 -22651 14482
rect -22617 14448 -22577 14482
rect -22543 14448 -22503 14482
rect -22469 14448 -22429 14482
rect -22395 14448 -22355 14482
rect -22321 14448 -22281 14482
rect -22247 14448 -22215 14482
rect -23687 14410 -22215 14448
rect -23687 14376 -23681 14410
rect -23647 14376 -23609 14410
rect -23575 14376 -23535 14410
rect -23501 14376 -23462 14410
rect -23428 14376 -23389 14410
rect -23355 14376 -23316 14410
rect -23282 14376 -23243 14410
rect -23209 14376 -23169 14410
rect -23135 14376 -23095 14410
rect -23061 14376 -23021 14410
rect -22987 14376 -22947 14410
rect -22913 14376 -22873 14410
rect -22839 14376 -22799 14410
rect -22765 14376 -22725 14410
rect -22691 14376 -22651 14410
rect -22617 14376 -22577 14410
rect -22543 14376 -22503 14410
rect -22469 14376 -22429 14410
rect -22395 14376 -22355 14410
rect -22321 14376 -22281 14410
rect -22247 14376 -22215 14410
rect -23687 14338 -22215 14376
rect -23687 14337 -23537 14338
rect -23687 14303 -23681 14337
rect -23647 14303 -23609 14337
rect -23575 14304 -23537 14337
rect -23503 14304 -23464 14338
rect -23430 14304 -23391 14338
rect -23357 14304 -23317 14338
rect -23283 14304 -23243 14338
rect -23209 14304 -23169 14338
rect -23135 14304 -23095 14338
rect -23061 14304 -23021 14338
rect -22987 14304 -22947 14338
rect -22913 14304 -22873 14338
rect -22839 14304 -22799 14338
rect -22765 14304 -22725 14338
rect -22691 14304 -22651 14338
rect -22617 14304 -22577 14338
rect -22543 14304 -22503 14338
rect -22469 14304 -22429 14338
rect -22395 14304 -22355 14338
rect -22321 14304 -22281 14338
rect -22247 14304 -22215 14338
rect -23575 14303 -22215 14304
rect -23687 14298 -22215 14303
rect -23687 14265 -23497 14298
rect -23687 14264 -23537 14265
rect -23687 14230 -23681 14264
rect -23647 14230 -23609 14264
rect -23575 14231 -23537 14264
rect -23503 14231 -23497 14265
rect -23575 14230 -23497 14231
rect -23687 14192 -23497 14230
rect -23687 14191 -23537 14192
rect -23687 14157 -23681 14191
rect -23647 14157 -23609 14191
rect -23575 14158 -23537 14191
rect -23503 14158 -23497 14192
rect -23575 14157 -23497 14158
rect -23687 14119 -23497 14157
rect -23687 14118 -23537 14119
rect -23687 14084 -23681 14118
rect -23647 14084 -23609 14118
rect -23575 14085 -23537 14118
rect -23503 14085 -23497 14119
rect -23575 14084 -23497 14085
rect -23687 14046 -23497 14084
rect -23687 14045 -23537 14046
rect -23687 14011 -23681 14045
rect -23647 14011 -23609 14045
rect -23575 14012 -23537 14045
rect -23503 14012 -23497 14046
rect -23575 14011 -23497 14012
rect -23687 13973 -23497 14011
rect -23687 13972 -23537 13973
rect -23687 13938 -23681 13972
rect -23647 13938 -23609 13972
rect -23575 13939 -23537 13972
rect -23503 13939 -23497 13973
rect -23575 13938 -23497 13939
rect -23687 13900 -23497 13938
rect -23687 13899 -23537 13900
rect -23687 13865 -23681 13899
rect -23647 13865 -23609 13899
rect -23575 13866 -23537 13899
rect -23503 13866 -23497 13900
rect -23575 13865 -23497 13866
rect -23687 13827 -23497 13865
rect -23687 13826 -23537 13827
rect -23687 13792 -23681 13826
rect -23647 13792 -23609 13826
rect -23575 13793 -23537 13826
rect -23503 13793 -23497 13827
rect -23575 13792 -23497 13793
rect -23687 13754 -23497 13792
rect -23687 13753 -23537 13754
rect -23687 13719 -23681 13753
rect -23647 13719 -23609 13753
rect -23575 13720 -23537 13753
rect -23503 13720 -23497 13754
rect -23575 13719 -23497 13720
rect -23687 13681 -23497 13719
rect -23687 13680 -23537 13681
rect -23687 13646 -23681 13680
rect -23647 13646 -23609 13680
rect -23575 13647 -23537 13680
rect -23503 13647 -23497 13681
rect -23575 13646 -23497 13647
rect -23687 13608 -23497 13646
rect -23687 13607 -23537 13608
rect -23687 13573 -23681 13607
rect -23647 13573 -23609 13607
rect -23575 13574 -23537 13607
rect -23503 13574 -23497 13608
rect -23575 13573 -23497 13574
rect -23687 13535 -23497 13573
rect -23687 13534 -23537 13535
rect -23687 13500 -23681 13534
rect -23647 13500 -23609 13534
rect -23575 13501 -23537 13534
rect -23503 13501 -23497 13535
rect -23575 13500 -23497 13501
rect -23687 13462 -23497 13500
rect -23687 13461 -23537 13462
rect -23687 13427 -23681 13461
rect -23647 13427 -23609 13461
rect -23575 13428 -23537 13461
rect -23503 13428 -23497 13462
rect -23575 13427 -23497 13428
rect -23687 13389 -23497 13427
rect -23687 13388 -23537 13389
rect -23687 13354 -23681 13388
rect -23647 13354 -23609 13388
rect -23575 13355 -23537 13388
rect -23503 13355 -23497 13389
rect -23575 13354 -23497 13355
rect -23687 13316 -23497 13354
rect -23687 13315 -23537 13316
rect -23687 13281 -23681 13315
rect -23647 13281 -23609 13315
rect -23575 13282 -23537 13315
rect -23503 13282 -23497 13316
rect -23575 13281 -23497 13282
rect -23687 13243 -23497 13281
rect -23687 13242 -23537 13243
rect -23687 13208 -23681 13242
rect -23647 13208 -23609 13242
rect -23575 13209 -23537 13242
rect -23503 13209 -23497 13243
rect -23575 13208 -23497 13209
rect -23687 13170 -23497 13208
rect -23687 13169 -23537 13170
rect -23687 13135 -23681 13169
rect -23647 13135 -23609 13169
rect -23575 13136 -23537 13169
rect -23503 13136 -23497 13170
rect -23575 13135 -23497 13136
rect -23687 13097 -23497 13135
rect -23687 13096 -23537 13097
rect -23687 13062 -23681 13096
rect -23647 13062 -23609 13096
rect -23575 13063 -23537 13096
rect -23503 13063 -23497 13097
rect -23575 13062 -23497 13063
rect -23687 13024 -23497 13062
rect -23687 13023 -23537 13024
rect -23687 12989 -23681 13023
rect -23647 12989 -23609 13023
rect -23575 12990 -23537 13023
rect -23503 12990 -23497 13024
rect -23575 12989 -23497 12990
rect -23687 12951 -23497 12989
rect -23687 12950 -23537 12951
rect -23687 12916 -23681 12950
rect -23647 12916 -23609 12950
rect -23575 12917 -23537 12950
rect -23503 12917 -23497 12951
rect -23575 12916 -23497 12917
rect -23687 12878 -23497 12916
rect -23687 12877 -23537 12878
rect -23687 12843 -23681 12877
rect -23647 12843 -23609 12877
rect -23575 12844 -23537 12877
rect -23503 12844 -23497 12878
rect -23575 12843 -23497 12844
rect -23687 12805 -23497 12843
rect -23687 12804 -23537 12805
rect -23687 12770 -23681 12804
rect -23647 12770 -23609 12804
rect -23575 12771 -23537 12804
rect -23503 12771 -23497 12805
rect -23575 12770 -23497 12771
rect -23687 12732 -23497 12770
rect -23687 12731 -23537 12732
rect -23687 12697 -23681 12731
rect -23647 12697 -23609 12731
rect -23575 12698 -23537 12731
rect -23503 12698 -23497 12732
rect -23575 12697 -23497 12698
rect -23687 12659 -23497 12697
rect -23687 12658 -23537 12659
rect -23687 12624 -23681 12658
rect -23647 12624 -23609 12658
rect -23575 12625 -23537 12658
rect -23503 12625 -23497 12659
rect -23575 12624 -23497 12625
rect -23687 12586 -23497 12624
rect -23687 12585 -23537 12586
rect -23687 12551 -23681 12585
rect -23647 12551 -23609 12585
rect -23575 12552 -23537 12585
rect -23503 12552 -23497 12586
rect -23575 12551 -23497 12552
rect -23687 12513 -23497 12551
rect -23687 12512 -23537 12513
rect -23687 12478 -23681 12512
rect -23647 12478 -23609 12512
rect -23575 12479 -23537 12512
rect -23503 12479 -23497 12513
rect -23575 12478 -23497 12479
rect -23687 12440 -23497 12478
rect -23687 12439 -23537 12440
rect -23687 12405 -23681 12439
rect -23647 12405 -23609 12439
rect -23575 12406 -23537 12439
rect -23503 12406 -23497 12440
rect -23575 12405 -23497 12406
rect -23687 12367 -23497 12405
rect -23687 12366 -23537 12367
rect -23687 12332 -23681 12366
rect -23647 12332 -23609 12366
rect -23575 12333 -23537 12366
rect -23503 12333 -23497 12367
rect -23575 12332 -23497 12333
rect -23687 12294 -23497 12332
rect -23687 12293 -23537 12294
rect -23687 12259 -23681 12293
rect -23647 12259 -23609 12293
rect -23575 12260 -23537 12293
rect -23503 12260 -23497 12294
rect -23575 12259 -23497 12260
rect -23687 12221 -23497 12259
rect -23687 12220 -23537 12221
rect -23687 12186 -23681 12220
rect -23647 12186 -23609 12220
rect -23575 12187 -23537 12220
rect -23503 12187 -23497 12221
rect -23575 12186 -23497 12187
rect -23687 12148 -23497 12186
rect -23687 12147 -23537 12148
rect -23687 7577 -23681 12147
rect -23575 12114 -23537 12147
rect -23503 12114 -23497 12148
rect -23575 12075 -23497 12114
rect -23503 7689 -23497 12075
rect -23363 14158 -22621 14164
rect -23363 14124 -23279 14158
rect -23245 14124 -23201 14158
rect -23167 14124 -23123 14158
rect -23089 14124 -23045 14158
rect -23011 14124 -22967 14158
rect -22933 14124 -22889 14158
rect -22855 14124 -22811 14158
rect -22777 14124 -22733 14158
rect -22699 14124 -22621 14158
rect -23363 14086 -22621 14124
rect -23363 14052 -23357 14086
rect -23323 14052 -23285 14086
rect -23251 14052 -23201 14086
rect -23167 14052 -23123 14086
rect -23089 14052 -23045 14086
rect -23011 14052 -22967 14086
rect -22933 14052 -22889 14086
rect -22855 14052 -22811 14086
rect -22777 14052 -22733 14086
rect -23363 14046 -22733 14052
rect -23363 14013 -23245 14046
rect -23363 13979 -23357 14013
rect -23323 13979 -23285 14013
rect -23251 13979 -23245 14013
rect -23363 13940 -23245 13979
rect -23363 13906 -23357 13940
rect -23323 13906 -23285 13940
rect -23251 13906 -23245 13940
rect -23363 13867 -23245 13906
rect -23363 13833 -23357 13867
rect -23323 13833 -23285 13867
rect -23251 13833 -23245 13867
rect -23363 13794 -23245 13833
rect -23363 13760 -23357 13794
rect -23323 13760 -23285 13794
rect -23251 13760 -23245 13794
rect -23363 13721 -23245 13760
rect -23363 13687 -23357 13721
rect -23323 13687 -23285 13721
rect -23251 13687 -23245 13721
rect -23363 13648 -23245 13687
rect -23363 13614 -23357 13648
rect -23323 13614 -23285 13648
rect -23251 13614 -23245 13648
rect -23363 13575 -23245 13614
rect -23363 13541 -23357 13575
rect -23323 13541 -23285 13575
rect -23251 13541 -23245 13575
rect -23363 13502 -23245 13541
rect -23363 13468 -23357 13502
rect -23323 13468 -23285 13502
rect -23251 13468 -23245 13502
rect -23363 13429 -23245 13468
rect -23363 7923 -23357 13429
rect -23251 7996 -23245 13429
rect -22739 13980 -22733 14046
rect -22627 13980 -22621 14086
rect -22739 13941 -22621 13980
rect -22739 13907 -22733 13941
rect -22699 13907 -22661 13941
rect -22627 13907 -22621 13941
rect -22739 13868 -22621 13907
rect -22739 13834 -22733 13868
rect -22699 13834 -22661 13868
rect -22627 13834 -22621 13868
rect -22739 13795 -22621 13834
rect -22739 13761 -22733 13795
rect -22699 13761 -22661 13795
rect -22627 13761 -22621 13795
rect -22739 13722 -22621 13761
rect -22739 13688 -22733 13722
rect -22699 13688 -22661 13722
rect -22627 13688 -22621 13722
rect -22739 13649 -22621 13688
rect -22739 13615 -22733 13649
rect -22699 13615 -22661 13649
rect -22627 13615 -22621 13649
rect -22739 13576 -22621 13615
rect -22739 13542 -22733 13576
rect -22699 13542 -22661 13576
rect -22627 13542 -22621 13576
rect -22739 13503 -22621 13542
rect -22739 13469 -22733 13503
rect -22699 13469 -22661 13503
rect -22627 13469 -22621 13503
rect -22739 13430 -22621 13469
rect -22739 13396 -22733 13430
rect -22699 13396 -22661 13430
rect -22627 13396 -22621 13430
rect -22739 13357 -22621 13396
rect -22739 13323 -22733 13357
rect -22699 13323 -22661 13357
rect -22627 13323 -22621 13357
rect -22739 13284 -22621 13323
rect -22739 13250 -22733 13284
rect -22699 13250 -22661 13284
rect -22627 13250 -22621 13284
rect -22739 13211 -22621 13250
rect -22739 13177 -22733 13211
rect -22699 13177 -22661 13211
rect -22627 13177 -22621 13211
rect -22739 13138 -22621 13177
rect -22739 13104 -22733 13138
rect -22699 13104 -22661 13138
rect -22627 13104 -22621 13138
rect -22739 13065 -22621 13104
rect -22739 13031 -22733 13065
rect -22699 13031 -22661 13065
rect -22627 13031 -22621 13065
rect -22739 12992 -22621 13031
rect -22739 12958 -22733 12992
rect -22699 12958 -22661 12992
rect -22627 12958 -22621 12992
rect -22739 12919 -22621 12958
rect -22739 12885 -22733 12919
rect -22699 12885 -22661 12919
rect -22627 12885 -22621 12919
rect -22739 12846 -22621 12885
rect -22739 12812 -22733 12846
rect -22699 12812 -22661 12846
rect -22627 12812 -22621 12846
rect -22739 12773 -22621 12812
rect -22739 12739 -22733 12773
rect -22699 12739 -22661 12773
rect -22627 12739 -22621 12773
rect -22739 12700 -22621 12739
rect -22739 12666 -22733 12700
rect -22699 12666 -22661 12700
rect -22627 12666 -22621 12700
rect -22739 12627 -22621 12666
rect -22739 12593 -22733 12627
rect -22699 12593 -22661 12627
rect -22627 12593 -22621 12627
rect -22739 12529 -22621 12593
rect -22739 12495 -22733 12529
rect -22699 12495 -22661 12529
rect -22627 12495 -22621 12529
rect -22739 12456 -22621 12495
rect -22739 12422 -22733 12456
rect -22699 12422 -22661 12456
rect -22627 12422 -22621 12456
rect -22739 12383 -22621 12422
rect -22739 12349 -22733 12383
rect -22699 12349 -22661 12383
rect -22627 12349 -22621 12383
rect -22739 12310 -22621 12349
rect -22739 12276 -22733 12310
rect -22699 12276 -22661 12310
rect -22627 12276 -22621 12310
rect -22739 12237 -22621 12276
rect -22739 12203 -22733 12237
rect -22699 12203 -22661 12237
rect -22627 12203 -22621 12237
rect -22739 12164 -22621 12203
rect -22739 12130 -22733 12164
rect -22699 12130 -22661 12164
rect -22627 12130 -22621 12164
rect -22739 12091 -22621 12130
rect -22739 12057 -22733 12091
rect -22699 12057 -22661 12091
rect -22627 12057 -22621 12091
rect -22739 12018 -22621 12057
rect -22739 11984 -22733 12018
rect -22699 11984 -22661 12018
rect -22627 11984 -22621 12018
rect -22739 11945 -22621 11984
rect -22739 11911 -22733 11945
rect -22699 11911 -22661 11945
rect -22627 11911 -22621 11945
rect -22739 11872 -22621 11911
rect -22739 11838 -22733 11872
rect -22699 11838 -22661 11872
rect -22627 11838 -22621 11872
rect -22739 11799 -22621 11838
rect -22739 11765 -22733 11799
rect -22699 11765 -22661 11799
rect -22627 11765 -22621 11799
rect -22739 11726 -22621 11765
rect -22739 11692 -22733 11726
rect -22699 11692 -22661 11726
rect -22627 11692 -22621 11726
rect -22739 11653 -22621 11692
rect -22739 11619 -22733 11653
rect -22699 11619 -22661 11653
rect -22627 11619 -22621 11653
rect -22739 11580 -22621 11619
rect -22739 11546 -22733 11580
rect -22699 11546 -22661 11580
rect -22627 11546 -22621 11580
rect -22739 11507 -22621 11546
rect -22739 11473 -22733 11507
rect -22699 11473 -22661 11507
rect -22627 11473 -22621 11507
rect -22739 11434 -22621 11473
rect -22739 11400 -22733 11434
rect -22699 11400 -22661 11434
rect -22627 11400 -22621 11434
rect -22739 11361 -22621 11400
rect -22739 11327 -22733 11361
rect -22699 11327 -22661 11361
rect -22627 11327 -22621 11361
rect -22739 11288 -22621 11327
rect -22739 11254 -22733 11288
rect -22699 11254 -22661 11288
rect -22627 11254 -22621 11288
rect -22739 11215 -22621 11254
rect -22739 11181 -22733 11215
rect -22699 11181 -22661 11215
rect -22627 11181 -22621 11215
rect -22739 11142 -22621 11181
rect -22739 11108 -22733 11142
rect -22699 11108 -22661 11142
rect -22627 11108 -22621 11142
rect -22739 11069 -22621 11108
rect -22739 11035 -22733 11069
rect -22699 11035 -22661 11069
rect -22627 11035 -22621 11069
rect -22739 10996 -22621 11035
rect -22739 10962 -22733 10996
rect -22699 10962 -22661 10996
rect -22627 10962 -22621 10996
rect -22739 10923 -22621 10962
rect -22739 10889 -22733 10923
rect -22699 10889 -22661 10923
rect -22627 10889 -22621 10923
rect -22739 10850 -22621 10889
rect -22739 10816 -22733 10850
rect -22699 10816 -22661 10850
rect -22627 10816 -22621 10850
rect -22739 10777 -22621 10816
rect -22739 10743 -22733 10777
rect -22699 10743 -22661 10777
rect -22627 10743 -22621 10777
rect -22739 10704 -22621 10743
rect -22739 10670 -22733 10704
rect -22699 10670 -22661 10704
rect -22627 10670 -22621 10704
rect -22739 10631 -22621 10670
rect -22739 10597 -22733 10631
rect -22699 10597 -22661 10631
rect -22627 10597 -22621 10631
rect -22739 10558 -22621 10597
rect -22739 10524 -22733 10558
rect -22699 10524 -22661 10558
rect -22627 10524 -22621 10558
rect -22739 10485 -22621 10524
rect -22739 10451 -22733 10485
rect -22699 10451 -22661 10485
rect -22627 10451 -22621 10485
rect -22739 10412 -22621 10451
rect -22739 10378 -22733 10412
rect -22699 10378 -22661 10412
rect -22627 10378 -22621 10412
rect -22739 10339 -22621 10378
rect -22739 10305 -22733 10339
rect -22699 10305 -22661 10339
rect -22627 10305 -22621 10339
rect -22739 10266 -22621 10305
rect -22739 10232 -22733 10266
rect -22699 10232 -22661 10266
rect -22627 10232 -22621 10266
rect -22739 10193 -22621 10232
rect -22739 10159 -22733 10193
rect -22699 10159 -22661 10193
rect -22627 10159 -22621 10193
rect -22739 10120 -22621 10159
rect -22739 10086 -22733 10120
rect -22699 10086 -22661 10120
rect -22627 10086 -22621 10120
rect -22739 10047 -22621 10086
rect -22739 10013 -22733 10047
rect -22699 10013 -22661 10047
rect -22627 10013 -22621 10047
rect -22739 9974 -22621 10013
rect -23093 9539 -23047 9551
rect -23093 9505 -23087 9539
rect -23053 9505 -23047 9539
rect -23093 9467 -23047 9505
rect -23093 9433 -23087 9467
rect -23053 9433 -23047 9467
rect -23093 9421 -23047 9433
rect -22937 9539 -22891 9551
rect -22937 9505 -22931 9539
rect -22897 9505 -22891 9539
rect -22937 9467 -22891 9505
rect -22937 9433 -22931 9467
rect -22897 9433 -22891 9467
rect -22937 9421 -22891 9433
rect -23171 9354 -23125 9366
rect -23171 9320 -23165 9354
rect -23131 9320 -23125 9354
rect -23171 9282 -23125 9320
rect -23171 9248 -23165 9282
rect -23131 9248 -23125 9282
rect -23171 9210 -23125 9248
rect -23171 9176 -23165 9210
rect -23131 9176 -23125 9210
rect -23171 9138 -23125 9176
rect -23018 9354 -22966 9366
rect -23018 9344 -23009 9354
rect -22975 9344 -22966 9354
rect -23018 9282 -22966 9292
rect -23018 9280 -23009 9282
rect -22975 9280 -22966 9282
rect -23018 9216 -22966 9228
rect -23018 9158 -22966 9164
tri -23018 9155 -23015 9158 ne
rect -23171 9104 -23165 9138
rect -23131 9104 -23125 9138
rect -23171 9066 -23125 9104
rect -23171 9032 -23165 9066
rect -23131 9032 -23125 9066
tri -23174 9012 -23171 9015 se
rect -23171 9012 -23125 9032
rect -23015 9138 -22969 9158
tri -22969 9155 -22966 9158 nw
rect -22859 9354 -22813 9366
rect -22859 9320 -22853 9354
rect -22819 9320 -22813 9354
rect -22859 9282 -22813 9320
rect -22859 9248 -22853 9282
rect -22819 9248 -22813 9282
rect -22859 9210 -22813 9248
rect -22859 9176 -22853 9210
rect -22819 9176 -22813 9210
rect -23015 9104 -23009 9138
rect -22975 9104 -22969 9138
rect -23015 9066 -22969 9104
rect -23015 9032 -23009 9066
rect -22975 9032 -22969 9066
rect -22859 9138 -22813 9176
rect -22859 9104 -22853 9138
rect -22819 9104 -22813 9138
rect -22859 9066 -22813 9104
tri -22864 9032 -22859 9037 se
rect -22859 9032 -22853 9066
rect -22819 9032 -22813 9066
tri -23125 9012 -23122 9015 sw
rect -23174 9006 -23122 9012
rect -23174 8942 -23122 8954
rect -23174 8888 -23165 8890
rect -23131 8888 -23122 8890
rect -23174 8878 -23122 8888
rect -23174 8816 -23165 8826
rect -23131 8816 -23122 8826
rect -23174 8804 -23122 8816
rect -23015 8994 -22969 9032
tri -22884 9012 -22864 9032 se
rect -22864 9012 -22813 9032
tri -22813 9012 -22810 9015 sw
rect -23015 8960 -23009 8994
rect -22975 8960 -22969 8994
rect -23015 8922 -22969 8960
rect -23015 8888 -23009 8922
rect -22975 8888 -22969 8922
rect -23015 8850 -22969 8888
rect -23015 8816 -23009 8850
rect -22975 8816 -22969 8850
rect -22928 9006 -22810 9012
rect -22876 8994 -22810 9006
rect -22876 8960 -22853 8994
rect -22819 8960 -22810 8994
rect -22876 8954 -22810 8960
rect -22928 8942 -22810 8954
rect -22876 8922 -22810 8942
rect -22876 8890 -22853 8922
rect -22928 8888 -22853 8890
rect -22819 8888 -22810 8922
rect -22928 8878 -22810 8888
rect -22876 8850 -22810 8878
rect -22876 8826 -22853 8850
rect -22928 8820 -22853 8826
tri -22878 8816 -22874 8820 ne
rect -22874 8816 -22853 8820
rect -22819 8816 -22810 8850
rect -23015 8804 -22969 8816
tri -22874 8804 -22862 8816 ne
rect -22862 8804 -22810 8816
tri -23245 7996 -23208 8033 sw
tri -22776 7996 -22739 8033 se
rect -22739 7996 -22733 9974
rect -22627 7996 -22621 9974
rect -23251 7963 -23208 7996
tri -23208 7963 -23175 7996 sw
tri -22809 7963 -22776 7996 se
rect -22776 7963 -22621 7996
rect -23251 7957 -22621 7963
rect -23251 7923 -23209 7957
rect -23175 7923 -23133 7957
rect -23099 7923 -23058 7957
rect -23024 7923 -22983 7957
rect -22949 7923 -22908 7957
rect -22874 7923 -22833 7957
rect -22799 7923 -22758 7957
rect -22724 7923 -22621 7957
rect -23363 7908 -22621 7923
rect -23363 7885 -22661 7908
rect -23363 7851 -23285 7885
rect -23251 7851 -23207 7885
rect -23173 7851 -23129 7885
rect -23095 7851 -23051 7885
rect -23017 7851 -22973 7885
rect -22939 7851 -22895 7885
rect -22861 7851 -22817 7885
rect -22783 7851 -22739 7885
rect -22705 7874 -22661 7885
rect -22627 7874 -22621 7908
rect -22705 7851 -22621 7874
rect -23363 7845 -22621 7851
rect -23503 7683 -22215 7689
rect -23503 7649 -23463 7683
rect -23429 7649 -23389 7683
rect -23355 7649 -23315 7683
rect -23281 7649 -23241 7683
rect -23207 7649 -23167 7683
rect -23133 7649 -23093 7683
rect -23059 7649 -23019 7683
rect -22985 7649 -22945 7683
rect -22911 7649 -22871 7683
rect -22837 7649 -22797 7683
rect -22763 7649 -22723 7683
rect -22689 7649 -22649 7683
rect -22615 7649 -22575 7683
rect -22541 7649 -22501 7683
rect -22467 7649 -22427 7683
rect -22393 7649 -22354 7683
rect -22320 7649 -22281 7683
rect -22247 7649 -22215 7683
rect -23575 7611 -22215 7649
rect -23575 7577 -23535 7611
rect -23501 7577 -23461 7611
rect -23427 7577 -23387 7611
rect -23353 7577 -23313 7611
rect -23279 7577 -23239 7611
rect -23205 7577 -23165 7611
rect -23131 7577 -23091 7611
rect -23057 7577 -23017 7611
rect -22983 7577 -22943 7611
rect -22909 7577 -22869 7611
rect -22835 7577 -22795 7611
rect -22761 7577 -22721 7611
rect -22687 7577 -22647 7611
rect -22613 7577 -22573 7611
rect -22539 7577 -22500 7611
rect -22466 7577 -22427 7611
rect -22393 7577 -22354 7611
rect -22320 7577 -22281 7611
rect -22247 7577 -22215 7611
rect -23687 7539 -22215 7577
rect -23687 7505 -23609 7539
rect -23575 7505 -23535 7539
rect -23501 7505 -23461 7539
rect -23427 7505 -23387 7539
rect -23353 7505 -23313 7539
rect -23279 7505 -23239 7539
rect -23205 7505 -23165 7539
rect -23131 7505 -23091 7539
rect -23057 7505 -23017 7539
rect -22983 7505 -22943 7539
rect -22909 7505 -22869 7539
rect -22835 7505 -22795 7539
rect -22761 7505 -22721 7539
rect -22687 7505 -22647 7539
rect -22613 7505 -22573 7539
rect -22539 7505 -22500 7539
rect -22466 7505 -22427 7539
rect -22393 7505 -22354 7539
rect -22320 7505 -22281 7539
rect -22247 7505 -22215 7539
rect -23687 7499 -22215 7505
rect -23215 3551 -22876 3557
rect -23215 3545 -22928 3551
rect -23215 3511 -23209 3545
rect -23175 3511 -22928 3545
rect -23215 3499 -22928 3511
rect -23215 3481 -22876 3499
rect -23215 3472 -22928 3481
rect -23215 3438 -23209 3472
rect -23175 3438 -22928 3472
rect -23215 3429 -22928 3438
rect -23215 3410 -22876 3429
rect -23215 3398 -22928 3410
rect -23215 3364 -23209 3398
rect -23175 3364 -22928 3398
rect -23215 3358 -22928 3364
rect -23215 3352 -22876 3358
rect -23304 3336 -23252 3342
rect -23304 3272 -23252 3284
rect -23059 3304 -23013 3316
rect -23059 3270 -23053 3304
rect -23019 3270 -23013 3304
rect -23059 3246 -23013 3270
rect -23252 3241 -22103 3246
tri -22103 3241 -22098 3246 sw
rect -23252 3232 -22098 3241
rect -23252 3220 -23053 3232
rect -23304 3214 -23053 3220
rect -23059 3198 -23053 3214
rect -23019 3214 -22098 3232
rect -23019 3198 -23013 3214
rect -23059 3186 -23013 3198
tri -22126 3186 -22098 3214 ne
tri -22098 3186 -22043 3241 sw
tri -22098 3154 -22066 3186 ne
rect -22066 3154 -1318 3186
rect -1370 1221 -1318 3154
rect -1370 1152 -1318 1169
rect -1370 1082 -1318 1100
rect -1370 1024 -1318 1030
rect -1074 1221 -1022 1227
rect -1074 1152 -1022 1169
rect -1074 1082 -1022 1100
tri 124 1050 127 1053 se
rect 127 1050 133 1053
rect -1074 1024 -1022 1030
rect -920 1044 133 1050
rect 185 1044 200 1053
rect 252 1044 267 1053
rect 319 1044 335 1053
rect 387 1044 403 1053
rect 455 1044 471 1053
rect 523 1044 539 1053
rect 591 1044 607 1053
rect -920 1010 -908 1044
rect -874 1010 -836 1044
rect -802 1010 -764 1044
rect -730 1010 -692 1044
rect -658 1010 -620 1044
rect -586 1010 -548 1044
rect -514 1010 -476 1044
rect -442 1010 -404 1044
rect -370 1010 -332 1044
rect -298 1010 -260 1044
rect -226 1010 -188 1044
rect -154 1010 -116 1044
rect -82 1010 -44 1044
rect -10 1010 28 1044
rect 62 1010 100 1044
rect 387 1010 388 1044
rect 455 1010 460 1044
rect 523 1010 532 1044
rect 591 1010 604 1044
rect -920 1004 133 1010
tri 124 1001 127 1004 ne
rect 127 1001 133 1004
rect 185 1001 200 1010
rect 252 1001 267 1010
rect 319 1001 335 1010
rect 387 1001 403 1010
rect 455 1001 471 1010
rect 523 1001 539 1010
rect 591 1001 607 1010
rect 659 1001 675 1053
rect 727 1001 743 1053
rect 795 1001 811 1053
rect 863 1001 879 1053
rect 931 1001 947 1053
rect 999 1050 1005 1053
tri 1005 1050 1008 1053 sw
rect 999 1044 1082 1050
rect 999 1010 1036 1044
rect 1070 1010 1082 1044
rect 999 1004 1082 1010
rect 999 1001 1005 1004
tri 1005 1001 1008 1004 nw
rect -1023 986 -977 998
rect -1023 952 -1017 986
rect -983 952 -977 986
rect -1023 912 -977 952
rect -1023 878 -1017 912
rect -983 878 -977 912
tri -847 894 -844 897 se
rect -844 894 -838 897
rect -1023 839 -977 878
rect -920 888 -838 894
rect -920 854 -908 888
rect -874 854 -838 888
rect -920 848 -838 854
tri -847 845 -844 848 ne
rect -844 845 -838 848
rect -786 845 -771 897
rect -719 845 -704 897
rect -652 845 -636 897
rect -584 845 -568 897
rect -516 888 -500 897
rect -448 888 -432 897
rect -380 888 -364 897
rect -312 888 -296 897
rect -244 888 -228 897
rect -176 888 -160 897
rect -108 888 -92 897
rect -40 888 -24 897
rect 28 894 34 897
tri 34 894 37 897 sw
rect 28 888 1082 894
rect -514 854 -500 888
rect -442 854 -432 888
rect -370 854 -364 888
rect -298 854 -296 888
rect 62 854 100 888
rect 134 854 172 888
rect 206 854 244 888
rect 278 854 316 888
rect 350 854 388 888
rect 422 854 460 888
rect 494 854 532 888
rect 566 854 604 888
rect 638 854 676 888
rect 710 854 748 888
rect 782 854 820 888
rect 854 854 892 888
rect 926 854 964 888
rect 998 854 1036 888
rect 1070 854 1082 888
rect -516 845 -500 854
rect -448 845 -432 854
rect -380 845 -364 854
rect -312 845 -296 854
rect -244 845 -228 854
rect -176 845 -160 854
rect -108 845 -92 854
rect -40 845 -24 854
rect 28 848 1082 854
rect 28 845 34 848
tri 34 845 37 848 nw
rect -1023 805 -1017 839
rect -983 805 -977 839
rect -1023 766 -977 805
rect -1023 732 -1017 766
rect -983 732 -977 766
tri 124 738 127 741 se
rect 127 738 133 741
rect -1023 693 -977 732
rect -1023 659 -1017 693
rect -983 659 -977 693
rect -920 732 133 738
rect 185 732 200 741
rect 252 732 267 741
rect 319 732 335 741
rect 387 732 403 741
rect 455 732 471 741
rect 523 732 539 741
rect 591 732 607 741
rect -920 698 -908 732
rect -874 698 -836 732
rect -802 698 -764 732
rect -730 698 -692 732
rect -658 698 -620 732
rect -586 698 -548 732
rect -514 698 -476 732
rect -442 698 -404 732
rect -370 698 -332 732
rect -298 698 -260 732
rect -226 698 -188 732
rect -154 698 -116 732
rect -82 698 -44 732
rect -10 698 28 732
rect 62 698 100 732
rect 387 698 388 732
rect 455 698 460 732
rect 523 698 532 732
rect 591 698 604 732
rect -920 692 133 698
tri 124 689 127 692 ne
rect 127 689 133 692
rect 185 689 200 698
rect 252 689 267 698
rect 319 689 335 698
rect 387 689 403 698
rect 455 689 471 698
rect 523 689 539 698
rect 591 689 607 698
rect 659 689 675 741
rect 727 689 743 741
rect 795 689 811 741
rect 863 689 879 741
rect 931 689 947 741
rect 999 738 1005 741
tri 1005 738 1008 741 sw
rect 999 732 1082 738
rect 999 698 1036 732
rect 1070 698 1082 732
rect 999 692 1082 698
rect 999 689 1005 692
tri 1005 689 1008 692 nw
rect -1023 620 -977 659
rect -1023 586 -1017 620
rect -983 586 -977 620
rect -1023 547 -977 586
tri -847 582 -844 585 se
rect -844 582 -838 585
rect -1023 513 -1017 547
rect -983 513 -977 547
rect -920 576 -838 582
rect -920 542 -908 576
rect -874 542 -838 576
rect -920 536 -838 542
tri -847 533 -844 536 ne
rect -844 533 -838 536
rect -786 533 -771 585
rect -719 533 -704 585
rect -652 533 -636 585
rect -584 533 -568 585
rect -516 576 -500 585
rect -448 576 -432 585
rect -380 576 -364 585
rect -312 576 -296 585
rect -244 576 -228 585
rect -176 576 -160 585
rect -108 576 -92 585
rect -40 576 -24 585
rect 28 582 34 585
tri 34 582 37 585 sw
rect 28 576 1082 582
rect -514 542 -500 576
rect -442 542 -432 576
rect -370 542 -364 576
rect -298 542 -296 576
rect 62 542 100 576
rect 134 542 172 576
rect 206 542 244 576
rect 278 542 316 576
rect 350 542 388 576
rect 422 542 460 576
rect 494 542 532 576
rect 566 542 604 576
rect 638 542 676 576
rect 710 542 748 576
rect 782 542 820 576
rect 854 542 892 576
rect 926 542 964 576
rect 998 542 1036 576
rect 1070 542 1082 576
rect -516 533 -500 542
rect -448 533 -432 542
rect -380 533 -364 542
rect -312 533 -296 542
rect -244 533 -228 542
rect -176 533 -160 542
rect -108 533 -92 542
rect -40 533 -24 542
rect 28 536 1082 542
rect 28 533 34 536
tri 34 533 37 536 nw
rect -1023 474 -977 513
rect -1023 440 -1017 474
rect -983 440 -977 474
rect -1023 401 -977 440
rect 88 429 1186 432
rect 88 426 133 429
rect -1023 367 -1017 401
rect -983 367 -977 401
rect -920 420 133 426
rect 185 420 200 429
rect 252 420 267 429
rect 319 420 335 429
rect 387 420 403 429
rect 455 420 471 429
rect 523 420 539 429
rect 591 420 607 429
rect -920 386 -908 420
rect -874 386 -836 420
rect -802 386 -764 420
rect -730 386 -692 420
rect -658 386 -620 420
rect -586 386 -548 420
rect -514 386 -476 420
rect -442 386 -404 420
rect -370 386 -332 420
rect -298 386 -260 420
rect -226 386 -188 420
rect -154 386 -116 420
rect -82 386 -44 420
rect -10 386 28 420
rect 62 386 100 420
rect 387 386 388 420
rect 455 386 460 420
rect 523 386 532 420
rect 591 386 604 420
rect -920 380 133 386
tri 124 377 127 380 ne
rect 127 377 133 380
rect 185 377 200 386
rect 252 377 267 386
rect 319 377 335 386
rect 387 377 403 386
rect 455 377 471 386
rect 523 377 539 386
rect 591 377 607 386
rect 659 377 675 429
rect 727 377 743 429
rect 795 377 811 429
rect 863 377 879 429
rect 931 377 947 429
rect 999 420 1186 429
rect 999 386 1036 420
rect 1070 386 1186 420
rect 999 380 1186 386
rect 999 377 1005 380
tri 1005 377 1008 380 nw
rect -1023 328 -977 367
rect -1023 294 -1017 328
rect -983 294 -977 328
rect -1023 255 -977 294
tri -847 270 -844 273 se
rect -844 270 -838 273
rect -1023 221 -1017 255
rect -983 221 -977 255
rect -920 264 -838 270
rect -920 230 -908 264
rect -874 230 -838 264
rect -920 224 -838 230
tri -847 221 -844 224 ne
rect -844 221 -838 224
rect -786 221 -771 273
rect -719 221 -704 273
rect -652 221 -636 273
rect -584 221 -568 273
rect -516 264 -500 273
rect -448 264 -432 273
rect -380 264 -364 273
rect -312 264 -296 273
rect -244 264 -228 273
rect -176 264 -160 273
rect -108 264 -92 273
rect -40 264 -24 273
rect 28 270 34 273
tri 34 270 37 273 sw
rect 28 264 1082 270
rect -514 230 -500 264
rect -442 230 -432 264
rect -370 230 -364 264
rect -298 230 -296 264
rect 62 230 100 264
rect 134 230 172 264
rect 206 230 244 264
rect 278 230 316 264
rect 350 230 388 264
rect 422 230 460 264
rect 494 230 532 264
rect 566 230 604 264
rect 638 230 676 264
rect 710 230 748 264
rect 782 230 820 264
rect 854 230 892 264
rect 926 230 964 264
rect 998 230 1036 264
rect 1070 230 1082 264
rect -516 221 -500 230
rect -448 221 -432 230
rect -380 221 -364 230
rect -312 221 -296 230
rect -244 221 -228 230
rect -176 221 -160 230
rect -108 221 -92 230
rect -40 221 -24 230
rect 28 224 1082 230
rect 28 221 34 224
tri 34 221 37 224 nw
rect -1023 182 -977 221
rect -1023 148 -1017 182
rect -983 148 -977 182
rect -1023 136 -977 148
rect -936 186 1197 192
rect -936 152 1079 186
rect 1113 152 1151 186
rect 1185 152 1197 186
rect -936 146 1197 152
tri 124 114 127 117 se
rect 127 114 133 117
rect -920 108 133 114
rect 185 108 200 117
rect 252 108 267 117
rect 319 108 335 117
rect 387 108 403 117
rect 455 108 471 117
rect 523 108 539 117
rect 591 108 607 117
rect -920 74 -908 108
rect -874 74 -836 108
rect -802 74 -764 108
rect -730 74 -692 108
rect -658 74 -620 108
rect -586 74 -548 108
rect -514 74 -476 108
rect -442 74 -404 108
rect -370 74 -332 108
rect -298 74 -260 108
rect -226 74 -188 108
rect -154 74 -116 108
rect -82 74 -44 108
rect -10 74 28 108
rect 62 74 100 108
rect 387 74 388 108
rect 455 74 460 108
rect 523 74 532 108
rect 591 74 604 108
rect -920 68 133 74
tri 124 65 127 68 ne
rect 127 65 133 68
rect 185 65 200 74
rect 252 65 267 74
rect 319 65 335 74
rect 387 65 403 74
rect 455 65 471 74
rect 523 65 539 74
rect 591 65 607 74
rect 659 65 675 117
rect 727 65 743 117
rect 795 65 811 117
rect 863 65 879 117
rect 931 65 947 117
rect 999 114 1005 117
tri 1005 114 1008 117 sw
rect 999 108 1186 114
rect 999 74 1036 108
rect 1070 74 1186 108
rect 999 68 1186 74
rect 999 65 1005 68
tri 1005 65 1008 68 nw
rect -23358 -1858 -23213 -1692
rect -23751 -2818 -23626 -2686
<< via1 >>
rect -23018 9320 -23009 9344
rect -23009 9320 -22975 9344
rect -22975 9320 -22966 9344
rect -23018 9292 -22966 9320
rect -23018 9248 -23009 9280
rect -23009 9248 -22975 9280
rect -22975 9248 -22966 9280
rect -23018 9228 -22966 9248
rect -23018 9210 -22966 9216
rect -23018 9176 -23009 9210
rect -23009 9176 -22975 9210
rect -22975 9176 -22966 9210
rect -23018 9164 -22966 9176
rect -23174 8994 -23122 9006
rect -23174 8960 -23165 8994
rect -23165 8960 -23131 8994
rect -23131 8960 -23122 8994
rect -23174 8954 -23122 8960
rect -23174 8922 -23122 8942
rect -23174 8890 -23165 8922
rect -23165 8890 -23131 8922
rect -23131 8890 -23122 8922
rect -23174 8850 -23122 8878
rect -23174 8826 -23165 8850
rect -23165 8826 -23131 8850
rect -23131 8826 -23122 8850
rect -22928 8954 -22876 9006
rect -22928 8890 -22876 8942
rect -22928 8826 -22876 8878
rect -22928 3545 -22876 3551
rect -22928 3511 -22918 3545
rect -22918 3511 -22884 3545
rect -22884 3511 -22876 3545
rect -22928 3499 -22876 3511
rect -22928 3472 -22876 3481
rect -22928 3438 -22918 3472
rect -22918 3438 -22884 3472
rect -22884 3438 -22876 3472
rect -22928 3429 -22876 3438
rect -22928 3398 -22876 3410
rect -22928 3364 -22918 3398
rect -22918 3364 -22884 3398
rect -22884 3364 -22876 3398
rect -22928 3358 -22876 3364
rect -23304 3284 -23252 3336
rect -23304 3220 -23252 3272
rect -1370 1169 -1318 1221
rect -1370 1100 -1318 1152
rect -1370 1030 -1318 1082
rect -1074 1169 -1022 1221
rect -1074 1100 -1022 1152
rect -1074 1030 -1022 1082
rect 133 1044 185 1053
rect 200 1044 252 1053
rect 267 1044 319 1053
rect 335 1044 387 1053
rect 403 1044 455 1053
rect 471 1044 523 1053
rect 539 1044 591 1053
rect 607 1044 659 1053
rect 133 1010 134 1044
rect 134 1010 172 1044
rect 172 1010 185 1044
rect 200 1010 206 1044
rect 206 1010 244 1044
rect 244 1010 252 1044
rect 267 1010 278 1044
rect 278 1010 316 1044
rect 316 1010 319 1044
rect 335 1010 350 1044
rect 350 1010 387 1044
rect 403 1010 422 1044
rect 422 1010 455 1044
rect 471 1010 494 1044
rect 494 1010 523 1044
rect 539 1010 566 1044
rect 566 1010 591 1044
rect 607 1010 638 1044
rect 638 1010 659 1044
rect 133 1001 185 1010
rect 200 1001 252 1010
rect 267 1001 319 1010
rect 335 1001 387 1010
rect 403 1001 455 1010
rect 471 1001 523 1010
rect 539 1001 591 1010
rect 607 1001 659 1010
rect 675 1044 727 1053
rect 675 1010 676 1044
rect 676 1010 710 1044
rect 710 1010 727 1044
rect 675 1001 727 1010
rect 743 1044 795 1053
rect 743 1010 748 1044
rect 748 1010 782 1044
rect 782 1010 795 1044
rect 743 1001 795 1010
rect 811 1044 863 1053
rect 811 1010 820 1044
rect 820 1010 854 1044
rect 854 1010 863 1044
rect 811 1001 863 1010
rect 879 1044 931 1053
rect 879 1010 892 1044
rect 892 1010 926 1044
rect 926 1010 931 1044
rect 879 1001 931 1010
rect 947 1044 999 1053
rect 947 1010 964 1044
rect 964 1010 998 1044
rect 998 1010 999 1044
rect 947 1001 999 1010
rect -838 888 -786 897
rect -838 854 -836 888
rect -836 854 -802 888
rect -802 854 -786 888
rect -838 845 -786 854
rect -771 888 -719 897
rect -771 854 -764 888
rect -764 854 -730 888
rect -730 854 -719 888
rect -771 845 -719 854
rect -704 888 -652 897
rect -704 854 -692 888
rect -692 854 -658 888
rect -658 854 -652 888
rect -704 845 -652 854
rect -636 888 -584 897
rect -636 854 -620 888
rect -620 854 -586 888
rect -586 854 -584 888
rect -636 845 -584 854
rect -568 888 -516 897
rect -500 888 -448 897
rect -432 888 -380 897
rect -364 888 -312 897
rect -296 888 -244 897
rect -228 888 -176 897
rect -160 888 -108 897
rect -92 888 -40 897
rect -24 888 28 897
rect -568 854 -548 888
rect -548 854 -516 888
rect -500 854 -476 888
rect -476 854 -448 888
rect -432 854 -404 888
rect -404 854 -380 888
rect -364 854 -332 888
rect -332 854 -312 888
rect -296 854 -260 888
rect -260 854 -244 888
rect -228 854 -226 888
rect -226 854 -188 888
rect -188 854 -176 888
rect -160 854 -154 888
rect -154 854 -116 888
rect -116 854 -108 888
rect -92 854 -82 888
rect -82 854 -44 888
rect -44 854 -40 888
rect -24 854 -10 888
rect -10 854 28 888
rect -568 845 -516 854
rect -500 845 -448 854
rect -432 845 -380 854
rect -364 845 -312 854
rect -296 845 -244 854
rect -228 845 -176 854
rect -160 845 -108 854
rect -92 845 -40 854
rect -24 845 28 854
rect 133 732 185 741
rect 200 732 252 741
rect 267 732 319 741
rect 335 732 387 741
rect 403 732 455 741
rect 471 732 523 741
rect 539 732 591 741
rect 607 732 659 741
rect 133 698 134 732
rect 134 698 172 732
rect 172 698 185 732
rect 200 698 206 732
rect 206 698 244 732
rect 244 698 252 732
rect 267 698 278 732
rect 278 698 316 732
rect 316 698 319 732
rect 335 698 350 732
rect 350 698 387 732
rect 403 698 422 732
rect 422 698 455 732
rect 471 698 494 732
rect 494 698 523 732
rect 539 698 566 732
rect 566 698 591 732
rect 607 698 638 732
rect 638 698 659 732
rect 133 689 185 698
rect 200 689 252 698
rect 267 689 319 698
rect 335 689 387 698
rect 403 689 455 698
rect 471 689 523 698
rect 539 689 591 698
rect 607 689 659 698
rect 675 732 727 741
rect 675 698 676 732
rect 676 698 710 732
rect 710 698 727 732
rect 675 689 727 698
rect 743 732 795 741
rect 743 698 748 732
rect 748 698 782 732
rect 782 698 795 732
rect 743 689 795 698
rect 811 732 863 741
rect 811 698 820 732
rect 820 698 854 732
rect 854 698 863 732
rect 811 689 863 698
rect 879 732 931 741
rect 879 698 892 732
rect 892 698 926 732
rect 926 698 931 732
rect 879 689 931 698
rect 947 732 999 741
rect 947 698 964 732
rect 964 698 998 732
rect 998 698 999 732
rect 947 689 999 698
rect -838 576 -786 585
rect -838 542 -836 576
rect -836 542 -802 576
rect -802 542 -786 576
rect -838 533 -786 542
rect -771 576 -719 585
rect -771 542 -764 576
rect -764 542 -730 576
rect -730 542 -719 576
rect -771 533 -719 542
rect -704 576 -652 585
rect -704 542 -692 576
rect -692 542 -658 576
rect -658 542 -652 576
rect -704 533 -652 542
rect -636 576 -584 585
rect -636 542 -620 576
rect -620 542 -586 576
rect -586 542 -584 576
rect -636 533 -584 542
rect -568 576 -516 585
rect -500 576 -448 585
rect -432 576 -380 585
rect -364 576 -312 585
rect -296 576 -244 585
rect -228 576 -176 585
rect -160 576 -108 585
rect -92 576 -40 585
rect -24 576 28 585
rect -568 542 -548 576
rect -548 542 -516 576
rect -500 542 -476 576
rect -476 542 -448 576
rect -432 542 -404 576
rect -404 542 -380 576
rect -364 542 -332 576
rect -332 542 -312 576
rect -296 542 -260 576
rect -260 542 -244 576
rect -228 542 -226 576
rect -226 542 -188 576
rect -188 542 -176 576
rect -160 542 -154 576
rect -154 542 -116 576
rect -116 542 -108 576
rect -92 542 -82 576
rect -82 542 -44 576
rect -44 542 -40 576
rect -24 542 -10 576
rect -10 542 28 576
rect -568 533 -516 542
rect -500 533 -448 542
rect -432 533 -380 542
rect -364 533 -312 542
rect -296 533 -244 542
rect -228 533 -176 542
rect -160 533 -108 542
rect -92 533 -40 542
rect -24 533 28 542
rect 133 420 185 429
rect 200 420 252 429
rect 267 420 319 429
rect 335 420 387 429
rect 403 420 455 429
rect 471 420 523 429
rect 539 420 591 429
rect 607 420 659 429
rect 133 386 134 420
rect 134 386 172 420
rect 172 386 185 420
rect 200 386 206 420
rect 206 386 244 420
rect 244 386 252 420
rect 267 386 278 420
rect 278 386 316 420
rect 316 386 319 420
rect 335 386 350 420
rect 350 386 387 420
rect 403 386 422 420
rect 422 386 455 420
rect 471 386 494 420
rect 494 386 523 420
rect 539 386 566 420
rect 566 386 591 420
rect 607 386 638 420
rect 638 386 659 420
rect 133 377 185 386
rect 200 377 252 386
rect 267 377 319 386
rect 335 377 387 386
rect 403 377 455 386
rect 471 377 523 386
rect 539 377 591 386
rect 607 377 659 386
rect 675 420 727 429
rect 675 386 676 420
rect 676 386 710 420
rect 710 386 727 420
rect 675 377 727 386
rect 743 420 795 429
rect 743 386 748 420
rect 748 386 782 420
rect 782 386 795 420
rect 743 377 795 386
rect 811 420 863 429
rect 811 386 820 420
rect 820 386 854 420
rect 854 386 863 420
rect 811 377 863 386
rect 879 420 931 429
rect 879 386 892 420
rect 892 386 926 420
rect 926 386 931 420
rect 879 377 931 386
rect 947 420 999 429
rect 947 386 964 420
rect 964 386 998 420
rect 998 386 999 420
rect 947 377 999 386
rect -838 264 -786 273
rect -838 230 -836 264
rect -836 230 -802 264
rect -802 230 -786 264
rect -838 221 -786 230
rect -771 264 -719 273
rect -771 230 -764 264
rect -764 230 -730 264
rect -730 230 -719 264
rect -771 221 -719 230
rect -704 264 -652 273
rect -704 230 -692 264
rect -692 230 -658 264
rect -658 230 -652 264
rect -704 221 -652 230
rect -636 264 -584 273
rect -636 230 -620 264
rect -620 230 -586 264
rect -586 230 -584 264
rect -636 221 -584 230
rect -568 264 -516 273
rect -500 264 -448 273
rect -432 264 -380 273
rect -364 264 -312 273
rect -296 264 -244 273
rect -228 264 -176 273
rect -160 264 -108 273
rect -92 264 -40 273
rect -24 264 28 273
rect -568 230 -548 264
rect -548 230 -516 264
rect -500 230 -476 264
rect -476 230 -448 264
rect -432 230 -404 264
rect -404 230 -380 264
rect -364 230 -332 264
rect -332 230 -312 264
rect -296 230 -260 264
rect -260 230 -244 264
rect -228 230 -226 264
rect -226 230 -188 264
rect -188 230 -176 264
rect -160 230 -154 264
rect -154 230 -116 264
rect -116 230 -108 264
rect -92 230 -82 264
rect -82 230 -44 264
rect -44 230 -40 264
rect -24 230 -10 264
rect -10 230 28 264
rect -568 221 -516 230
rect -500 221 -448 230
rect -432 221 -380 230
rect -364 221 -312 230
rect -296 221 -244 230
rect -228 221 -176 230
rect -160 221 -108 230
rect -92 221 -40 230
rect -24 221 28 230
rect 133 108 185 117
rect 200 108 252 117
rect 267 108 319 117
rect 335 108 387 117
rect 403 108 455 117
rect 471 108 523 117
rect 539 108 591 117
rect 607 108 659 117
rect 133 74 134 108
rect 134 74 172 108
rect 172 74 185 108
rect 200 74 206 108
rect 206 74 244 108
rect 244 74 252 108
rect 267 74 278 108
rect 278 74 316 108
rect 316 74 319 108
rect 335 74 350 108
rect 350 74 387 108
rect 403 74 422 108
rect 422 74 455 108
rect 471 74 494 108
rect 494 74 523 108
rect 539 74 566 108
rect 566 74 591 108
rect 607 74 638 108
rect 638 74 659 108
rect 133 65 185 74
rect 200 65 252 74
rect 267 65 319 74
rect 335 65 387 74
rect 403 65 455 74
rect 471 65 523 74
rect 539 65 591 74
rect 607 65 659 74
rect 675 108 727 117
rect 675 74 676 108
rect 676 74 710 108
rect 710 74 727 108
rect 675 65 727 74
rect 743 108 795 117
rect 743 74 748 108
rect 748 74 782 108
rect 782 74 795 108
rect 743 65 795 74
rect 811 108 863 117
rect 811 74 820 108
rect 820 74 854 108
rect 854 74 863 108
rect 811 65 863 74
rect 879 108 931 117
rect 879 74 892 108
rect 892 74 926 108
rect 926 74 931 108
rect 879 65 931 74
rect 947 108 999 117
rect 947 74 964 108
rect 964 74 998 108
rect 998 74 999 108
rect 947 65 999 74
<< metal2 >>
rect -23018 9344 -22966 9350
tri -23049 9305 -23018 9336 se
rect -23484 9292 -23018 9305
rect -23484 9280 -22966 9292
rect -23484 9253 -23018 9280
rect -23484 9228 -23427 9253
tri -23427 9228 -23402 9253 nw
tri -23048 9228 -23023 9253 ne
rect -23023 9228 -23018 9253
rect -23484 3342 -23432 9228
tri -23432 9223 -23427 9228 nw
tri -23023 9223 -23018 9228 ne
rect -23018 9216 -22966 9228
rect -23018 9158 -22966 9164
rect -23174 9006 -22876 9012
rect -23122 8954 -22928 9006
rect -23174 8942 -22876 8954
rect -23122 8890 -22928 8942
rect -23174 8878 -22876 8890
rect -23122 8826 -22928 8878
rect -23174 8820 -22876 8826
rect -22928 3551 -22876 8820
rect -22928 3481 -22876 3499
rect -22928 3410 -22876 3429
rect -22928 3352 -22876 3358
rect -23484 3336 -23252 3342
rect -23484 3290 -23304 3336
rect -23304 3272 -23252 3284
rect -23304 3214 -23252 3220
rect -1370 1221 -1022 1227
rect -1318 1169 -1074 1221
rect -1370 1152 -1022 1169
rect -1318 1100 -1074 1152
rect -1370 1082 -1022 1100
rect -1318 1030 -1074 1082
rect -1370 1024 -1022 1030
rect -844 897 34 1151
rect 127 1053 1005 1080
rect 127 1001 133 1053
rect 185 1001 200 1053
rect 252 1001 267 1053
rect 319 1001 335 1053
rect 387 1001 403 1053
rect 455 1001 471 1053
rect 523 1001 539 1053
rect 591 1001 607 1053
rect 659 1001 675 1053
rect 727 1001 743 1053
rect 795 1001 811 1053
rect 863 1001 879 1053
rect 931 1001 947 1053
rect 999 1001 1005 1053
rect 127 924 1005 1001
rect 128 922 1004 923
rect -844 845 -838 897
rect -786 845 -771 897
rect -719 845 -704 897
rect -652 845 -636 897
rect -584 845 -568 897
rect -516 845 -500 897
rect -448 845 -432 897
rect -380 845 -364 897
rect -312 845 -296 897
rect -244 845 -228 897
rect -176 845 -160 897
rect -108 845 -92 897
rect -40 845 -24 897
rect 28 845 34 897
rect -844 585 34 845
rect -844 533 -838 585
rect -786 533 -771 585
rect -719 533 -704 585
rect -652 533 -636 585
rect -584 533 -568 585
rect -516 533 -500 585
rect -448 533 -432 585
rect -380 533 -364 585
rect -312 533 -296 585
rect -244 533 -228 585
rect -176 533 -160 585
rect -108 533 -92 585
rect -40 533 -24 585
rect 28 533 34 585
rect -844 273 34 533
rect -844 221 -838 273
rect -786 221 -771 273
rect -719 221 -704 273
rect -652 221 -636 273
rect -584 221 -568 273
rect -516 221 -500 273
rect -448 221 -432 273
rect -380 221 -364 273
rect -312 221 -296 273
rect -244 221 -228 273
rect -176 221 -160 273
rect -108 221 -92 273
rect -40 221 -24 273
rect 28 221 34 273
rect 128 861 1004 862
rect 127 741 1005 860
rect 127 689 133 741
rect 185 689 200 741
rect 252 689 267 741
rect 319 689 335 741
rect 387 689 403 741
rect 455 689 471 741
rect 523 689 539 741
rect 591 689 607 741
rect 659 689 675 741
rect 727 689 743 741
rect 795 689 811 741
rect 863 689 879 741
rect 931 689 947 741
rect 999 689 1005 741
rect 127 429 1005 689
rect 127 377 133 429
rect 185 377 200 429
rect 252 377 267 429
rect 319 377 335 429
rect 387 377 403 429
rect 455 377 471 429
rect 523 377 539 429
rect 591 377 607 429
rect 659 377 675 429
rect 727 377 743 429
rect 795 377 811 429
rect 863 377 879 429
rect 931 377 947 429
rect 999 377 1005 429
rect 127 117 1005 377
rect 127 65 133 117
rect 185 65 200 117
rect 252 65 267 117
rect 319 65 335 117
rect 387 65 403 117
rect 455 65 471 117
rect 523 65 539 117
rect 591 65 607 117
rect 659 65 675 117
rect 727 65 743 117
rect 795 65 811 117
rect 863 65 879 117
rect 931 65 947 117
rect 999 65 1005 117
<< rmetal2 >>
rect 127 923 1005 924
rect 127 922 128 923
rect 1004 922 1005 923
rect 127 861 128 862
rect 1004 861 1005 862
rect 127 860 1005 861
use sky130_fd_pr__pfet_01v8__example_5595914180837  sky130_fd_pr__pfet_01v8__example_5595914180837_0
timestamp 1619862920
transform 1 0 -23164 0 -1 3598
box -28 0 284 267
use sky130_fd_pr__pfet_01v8__example_5595914180845  sky130_fd_pr__pfet_01v8__example_5595914180845_0
timestamp 1619862920
transform 0 -1 1066 1 0 119
box -28 0 908 985
use sky130_fd_io__tk_em2o_cdns_5595914180844  sky130_fd_io__tk_em2o_cdns_5595914180844_0
timestamp 1619862920
transform 0 -1 1005 1 0 808
box 0 24 168 28
use sky130_fd_io__gpio_ovtv2_hotswap_guardrings  sky130_fd_io__gpio_ovtv2_hotswap_guardrings_0
timestamp 1619862920
transform 1 0 -24510 0 1 -3388
box 0 0 26980 8664
use sky130_fd_pr__nfet_01v8__example_5595914180834  sky130_fd_pr__nfet_01v8__example_5595914180834_0
timestamp 1619862920
transform 1 0 -23120 0 1 8820
box -28 0 284 265
<< labels >>
flabel metal1 s -23358 -1858 -23213 -1692 3 FreeSans 520 0 0 0 VPB_DRVR
port 1 nsew
flabel metal1 s -23751 -2818 -23626 -2686 3 FreeSans 520 0 0 0 VSSD
port 2 nsew
flabel metal1 s -22716 8796 -22642 8884 3 FreeSans 520 0 0 0 VSSIO
port 3 nsew
flabel metal1 s -22782 3214 -22739 3246 3 FreeSans 520 0 0 0 PUG_H
port 4 nsew
flabel metal2 s -22928 3712 -22876 3763 3 FreeSans 520 0 0 0 PU_H_N
port 5 nsew
flabel metal2 s -628 561 -396 660 3 FreeSans 520 0 0 0 VDDIO
port 6 nsew
flabel metal2 s 416 590 605 664 3 FreeSans 520 0 0 0 PAD
port 7 nsew
flabel locali s -23015 9462 -22971 9510 3 FreeSans 520 0 0 0 NGHS_H
port 8 nsew
flabel locali s -23089 3646 -23054 3680 3 FreeSans 520 0 0 0 PGHS_H
port 9 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 43690064
string GDS_START 43541348
<< end >>
