magic
tech sky130A
magscale 1 2
timestamp 1619862920
<< checkpaint >>
rect -1260 -1402 16260 40711
use sky130_fd_io__top_gpio_pad  sky130_fd_io__top_gpio_pad_0
timestamp 1619862920
transform 1 0 0 0 1 0
box 960 18991 14040 34071
use sky130_fd_io__com_bus_hookup  sky130_fd_io__com_bus_hookup_0
timestamp 1619862920
transform 1 0 0 0 1 0
box 0 -142 15000 39451
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 7008154
string GDS_START 7008048
<< end >>
